-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Apr 5 2020 01:05:17

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    ioFifoData : inout std_logic_vector(7 downto 0);
    P1A9 : out std_logic;
    P1A1 : in std_logic;
    P1A8 : out std_logic;
    oRx_n : out std_logic;
    P1A7 : out std_logic;
    P1A3 : out std_logic;
    iTxE_n : in std_logic;
    iRxF_n : in std_logic;
    iClk : in std_logic;
    P1A2 : out std_logic;
    BTN_N : in std_logic;
    BTN1 : in std_logic;
    oTx_n : out std_logic;
    P1A4 : out std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__17429\ : std_logic;
signal \N__17415\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17406\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17397\ : std_logic;
signal \N__17396\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17378\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17361\ : std_logic;
signal \N__17360\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17352\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17333\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17325\ : std_logic;
signal \N__17324\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17306\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17298\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17287\ : std_logic;
signal \N__17280\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17271\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17262\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17253\ : std_logic;
signal \N__17252\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17244\ : std_logic;
signal \N__17243\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17225\ : std_logic;
signal \N__17222\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17203\ : std_logic;
signal \N__17200\ : std_logic;
signal \N__17195\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17182\ : std_logic;
signal \N__17179\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17168\ : std_logic;
signal \N__17165\ : std_logic;
signal \N__17162\ : std_logic;
signal \N__17159\ : std_logic;
signal \N__17156\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17144\ : std_logic;
signal \N__17141\ : std_logic;
signal \N__17138\ : std_logic;
signal \N__17135\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17111\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17096\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17078\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17069\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17061\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17028\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17016\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17006\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16991\ : std_logic;
signal \N__16990\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16988\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16985\ : std_logic;
signal \N__16984\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16982\ : std_logic;
signal \N__16981\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16979\ : std_logic;
signal \N__16978\ : std_logic;
signal \N__16977\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16974\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16968\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16965\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16962\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16959\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16956\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16950\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16944\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16941\ : std_logic;
signal \N__16940\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16938\ : std_logic;
signal \N__16937\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16935\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16930\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16926\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16921\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16914\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16912\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16903\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16901\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16898\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16699\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16696\ : std_logic;
signal \N__16695\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16693\ : std_logic;
signal \N__16690\ : std_logic;
signal \N__16689\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16683\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16680\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16677\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16674\ : std_logic;
signal \N__16671\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16662\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16660\ : std_logic;
signal \N__16659\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16657\ : std_logic;
signal \N__16654\ : std_logic;
signal \N__16653\ : std_logic;
signal \N__16650\ : std_logic;
signal \N__16649\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16644\ : std_logic;
signal \N__16641\ : std_logic;
signal \N__16640\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16638\ : std_logic;
signal \N__16637\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16622\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16619\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16610\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16594\ : std_logic;
signal \N__16589\ : std_logic;
signal \N__16580\ : std_logic;
signal \N__16577\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16541\ : std_logic;
signal \N__16538\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16518\ : std_logic;
signal \N__16511\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16466\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16455\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16453\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16438\ : std_logic;
signal \N__16437\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16425\ : std_logic;
signal \N__16422\ : std_logic;
signal \N__16421\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16419\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16416\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16413\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16395\ : std_logic;
signal \N__16392\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16386\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16384\ : std_logic;
signal \N__16381\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16375\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16369\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16357\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16352\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16347\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16340\ : std_logic;
signal \N__16217\ : std_logic;
signal \N__16214\ : std_logic;
signal \N__16211\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16196\ : std_logic;
signal \N__16193\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16172\ : std_logic;
signal \N__16169\ : std_logic;
signal \N__16166\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16159\ : std_logic;
signal \N__16156\ : std_logic;
signal \N__16153\ : std_logic;
signal \N__16148\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16137\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16115\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16111\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16105\ : std_logic;
signal \N__16100\ : std_logic;
signal \N__16097\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16082\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16049\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16032\ : std_logic;
signal \N__16029\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16014\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15974\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15969\ : std_logic;
signal \N__15966\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15933\ : std_logic;
signal \N__15930\ : std_logic;
signal \N__15927\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15922\ : std_logic;
signal \N__15921\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15864\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15832\ : std_logic;
signal \N__15829\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15823\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15794\ : std_logic;
signal \N__15791\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15731\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15692\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15688\ : std_logic;
signal \N__15685\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15677\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15671\ : std_logic;
signal \N__15668\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15662\ : std_logic;
signal \N__15659\ : std_logic;
signal \N__15656\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15654\ : std_logic;
signal \N__15651\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15616\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15605\ : std_logic;
signal \N__15602\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15596\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15557\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15545\ : std_logic;
signal \N__15542\ : std_logic;
signal \N__15539\ : std_logic;
signal \N__15536\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15524\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15505\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15497\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15490\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15445\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15431\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15416\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15367\ : std_logic;
signal \N__15366\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15363\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15358\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15320\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15304\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15277\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15257\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15246\ : std_logic;
signal \N__15243\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15203\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15195\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15168\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15149\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15104\ : std_logic;
signal \N__15101\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15099\ : std_logic;
signal \N__15096\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15066\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15042\ : std_logic;
signal \N__15039\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15004\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14949\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14946\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14943\ : std_logic;
signal \N__14940\ : std_logic;
signal \N__14937\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14931\ : std_logic;
signal \N__14928\ : std_logic;
signal \N__14925\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14890\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14884\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14873\ : std_logic;
signal \N__14870\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14852\ : std_logic;
signal \N__14849\ : std_logic;
signal \N__14846\ : std_logic;
signal \N__14843\ : std_logic;
signal \N__14842\ : std_logic;
signal \N__14841\ : std_logic;
signal \N__14840\ : std_logic;
signal \N__14837\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14831\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14807\ : std_logic;
signal \N__14804\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14796\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14756\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14743\ : std_logic;
signal \N__14740\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14728\ : std_logic;
signal \N__14725\ : std_logic;
signal \N__14722\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14668\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14660\ : std_logic;
signal \N__14657\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14639\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14599\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14555\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14549\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14544\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14537\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14529\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14523\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14517\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14501\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14494\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14448\ : std_logic;
signal \N__14445\ : std_logic;
signal \N__14442\ : std_logic;
signal \N__14439\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14428\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14418\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14409\ : std_logic;
signal \N__14406\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14397\ : std_logic;
signal \N__14394\ : std_logic;
signal \N__14391\ : std_logic;
signal \N__14388\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14366\ : std_logic;
signal \N__14363\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14325\ : std_logic;
signal \N__14322\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14309\ : std_logic;
signal \N__14308\ : std_logic;
signal \N__14307\ : std_logic;
signal \N__14304\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14288\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14274\ : std_logic;
signal \N__14271\ : std_logic;
signal \N__14268\ : std_logic;
signal \N__14265\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14255\ : std_logic;
signal \N__14252\ : std_logic;
signal \N__14249\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14238\ : std_logic;
signal \N__14235\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14208\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14183\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14175\ : std_logic;
signal \N__14172\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14156\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14154\ : std_logic;
signal \N__14151\ : std_logic;
signal \N__14148\ : std_logic;
signal \N__14145\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14131\ : std_logic;
signal \N__14130\ : std_logic;
signal \N__14127\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14121\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14108\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14100\ : std_logic;
signal \N__14097\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14082\ : std_logic;
signal \N__14081\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14075\ : std_logic;
signal \N__14072\ : std_logic;
signal \N__14069\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14052\ : std_logic;
signal \N__14049\ : std_logic;
signal \N__14046\ : std_logic;
signal \N__14039\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14022\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14016\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14004\ : std_logic;
signal \N__14003\ : std_logic;
signal \N__14000\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13986\ : std_logic;
signal \N__13983\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13971\ : std_logic;
signal \N__13968\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13956\ : std_logic;
signal \N__13953\ : std_logic;
signal \N__13950\ : std_logic;
signal \N__13947\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13875\ : std_logic;
signal \N__13872\ : std_logic;
signal \N__13869\ : std_logic;
signal \N__13866\ : std_logic;
signal \N__13857\ : std_logic;
signal \N__13854\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13848\ : std_logic;
signal \N__13845\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13836\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13824\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13819\ : std_logic;
signal \N__13818\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13799\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13781\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13779\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13775\ : std_logic;
signal \N__13772\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13746\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13738\ : std_logic;
signal \N__13735\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13707\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13685\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13679\ : std_logic;
signal \N__13676\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13630\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13625\ : std_logic;
signal \N__13622\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13600\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13597\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13592\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13551\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13548\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13545\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13543\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13483\ : std_logic;
signal \N__13480\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13441\ : std_logic;
signal \N__13438\ : std_logic;
signal \N__13435\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13414\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13382\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13372\ : std_logic;
signal \N__13371\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13345\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13337\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13327\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13318\ : std_logic;
signal \N__13317\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13315\ : std_logic;
signal \N__13312\ : std_logic;
signal \N__13309\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13299\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13291\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13263\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13255\ : std_logic;
signal \N__13254\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13242\ : std_logic;
signal \N__13239\ : std_logic;
signal \N__13236\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13146\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13094\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13058\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13034\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13028\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13003\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12968\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12931\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12878\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12851\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12847\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12841\ : std_logic;
signal \N__12838\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12793\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12787\ : std_logic;
signal \N__12784\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12775\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12769\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12757\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12754\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12652\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12634\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12589\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12577\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12515\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12279\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12261\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12189\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11860\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10765\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9710\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7963\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6449\ : std_logic;
signal \INVfifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net\ : std_logic;
signal \INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net\ : std_logic;
signal \BTN_N_c\ : std_logic;
signal \INVfifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net\ : std_logic;
signal \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_0\ : std_logic;
signal \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_1\ : std_logic;
signal \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_2\ : std_logic;
signal \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_3\ : std_logic;
signal \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_4\ : std_logic;
signal \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_5\ : std_logic;
signal \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_6\ : std_logic;
signal \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_7\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_8\ : std_logic;
signal \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_9\ : std_logic;
signal \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_10\ : std_logic;
signal \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_11\ : std_logic;
signal \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_12\ : std_logic;
signal \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_13\ : std_logic;
signal \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_8\ : std_logic;
signal \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_7\ : std_logic;
signal \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_14\ : std_logic;
signal \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_10\ : std_logic;
signal \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_11\ : std_logic;
signal \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_12\ : std_logic;
signal \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_9\ : std_logic;
signal \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_13\ : std_logic;
signal \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_6\ : std_logic;
signal \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_5\ : std_logic;
signal \uart_inst0.uart_inst0.un1_rx_clk_divider_10\ : std_logic;
signal \uart_inst0.uart_inst0.un1_rx_clk_divider_9\ : std_logic;
signal \uart_inst0.uart_inst0.un1_rx_clk_divider_7_cascade_\ : std_logic;
signal \uart_inst0.uart_inst0.un1_rx_clk_divider_0_cascade_\ : std_logic;
signal \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_3\ : std_logic;
signal \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_1\ : std_logic;
signal \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_4\ : std_logic;
signal \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_2\ : std_logic;
signal \uart_inst0.uart_inst0.un1_rx_clk_divider_8\ : std_logic;
signal \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_0\ : std_logic;
signal \uart_inst0.uart_inst0.rx_clk_divider_1_sqmuxa_i\ : std_logic;
signal \P1A3_c\ : std_logic;
signal \N_86_mux\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_0_cascade_\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_6\ : std_logic;
signal \GB_BUFFER_wPllLocked_i_g_THRU_CO\ : std_logic;
signal \fifo_inst_tx_fifo_inst_wRamWrEn_cascade_\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.m68_eZ0Z_5_cascade_\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.m68_eZ0Z_6\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.N_92\ : std_logic;
signal \fifo_inst_tx_fifo_inst_rRamWrAddr_0\ : std_logic;
signal \rRamWrAddr_RNI10581_0\ : std_logic;
signal \bfn_13_2_0_\ : std_logic;
signal \fifo_inst_tx_fifo_inst_rRamWrAddr_1\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_0\ : std_logic;
signal \fifo_inst_tx_fifo_inst_rRamWrAddr_2\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_1\ : std_logic;
signal \fifo_inst_tx_fifo_inst_rRamWrAddr_3\ : std_logic;
signal \un1_rRamWrAddr_cry_2_c_RNISJKU\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_2\ : std_logic;
signal \fifo_inst_tx_fifo_inst_rRamWrAddr_4\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_3\ : std_logic;
signal \fifo_inst_tx_fifo_inst_rRamWrAddr_5\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_4\ : std_logic;
signal \fifo_inst_tx_fifo_inst_rRamWrAddr_6\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_5\ : std_logic;
signal \fifo_inst_tx_fifo_inst_rRamWrAddr_7\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_6\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_7\ : std_logic;
signal \bfn_13_3_0_\ : std_logic;
signal \fifo_inst_tx_fifo_inst_rRamWrAddr_8\ : std_logic;
signal \fifo_inst_ft2232h_inst_un1_rFifoState_12_0_i_cascade_\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rDataCount_ac0_1_a1_1\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.m78_bmZ0\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.m78_nsZ0Z_1_cascade_\ : std_logic;
signal \fifo_inst.ft2232h_inst.un1_rFifoState_12_0_i_0\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c2_d_cascade_\ : std_logic;
signal \N_84_mux_cascade_\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.m65_bmZ0_cascade_\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rDataCount_c2_1_1_0_cascade_\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.m65_nsZ0Z_1\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rDataCount_c2_1\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rDataCount_0_sqmuxa\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rDataCount_ac0_2\ : std_logic;
signal \rUartTxEnZ0\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c3_0_0\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c2_d\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rDataCount_0_sqmuxa\ : std_logic;
signal \uart_inst0.wTxRdEmpty_cascade_\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_0\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_1\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_2\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_3\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_4\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_5\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_6\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_7\ : std_logic;
signal \INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ1Z_0\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNO_0Z0Z_0\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ1Z_1\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_0\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ0Z_2\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_1\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_3\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNO_0Z0Z_3\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_2\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_3\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_4\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_5\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_6\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_7\ : std_logic;
signal \bfn_13_13_0_\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_8\ : std_logic;
signal \uart_inst0.wTxRdData_0\ : std_logic;
signal \uart_inst0.wTxRdData_1\ : std_logic;
signal \uart_inst0.uart_inst0.rTxDataZ0Z_1\ : std_logic;
signal \uart_inst0.wTxRdData_6\ : std_logic;
signal \uart_inst0.wTxRdData_3\ : std_logic;
signal \uart_inst0.wTxRdData_4\ : std_logic;
signal \uart_inst0.uart_inst0.rTxDataZ0Z_4\ : std_logic;
signal \uart_inst0.uart_inst0.rTxDataZ0Z_3\ : std_logic;
signal \uart_inst0.wTxRdData_2\ : std_logic;
signal \uart_inst0.uart_inst0.rTxDataZ0Z_2\ : std_logic;
signal \uart_inst0.uart_inst0.rTxDataZ0Z_6\ : std_logic;
signal \uart_inst0.wTxRdData_5\ : std_logic;
signal \uart_inst0.uart_inst0.rTxDataZ0Z_5\ : std_logic;
signal \uart_inst0.wTxRdData_7\ : std_logic;
signal \uart_inst0.uart_inst0.rTxDataZ0Z_7\ : std_logic;
signal \N_97_cascade_\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.m8_xZ0Z0_cascade_\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rDataCount_axbxc3_2_tz\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rDataCount_axbxc3_a0_2\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rDataCount_c2_0\ : std_logic;
signal \fifo_inst_tx_fifo_inst_wRamWrEn\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rDataCount_ac0_1_a0_0\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rDataCount_c2_1_cascade_\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rDataCount_ac0_2\ : std_logic;
signal \fifo_inst_tx_fifo_inst_un1_rDataCount15_2_0_0\ : std_logic;
signal \fifo_inst_tx_fifo_inst_rDataCount_2\ : std_logic;
signal \fifo_inst_tx_fifo_inst_rDataCount_1\ : std_logic;
signal \fifo_inst_tx_fifo_inst_rDataCount_fast_3\ : std_logic;
signal \fifo_inst_tx_fifo_inst_rDataCount_0\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rDataCount_axbxc3_1_1_cascade_\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.m15_xZ0Z0_cascade_\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rDataCount_axbxc3_1_1\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rDataCount_fast_3\ : std_logic;
signal \P1A4_c\ : std_logic;
signal \fifo_inst_ft2232h_inst_rFifoState_3\ : std_logic;
signal \fifo_inst_rx_fifo_inst_un1_rDataCount15_2_0_0\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rDataCount_fast_0\ : std_logic;
signal \N_84_mux\ : std_logic;
signal \rUartTxEn_4_cascade_\ : std_logic;
signal \rFtdiRxStateZ0Z_0\ : std_logic;
signal \fifo_inst.ft2232h_inst.rFifoStatesr_0\ : std_logic;
signal \fifo_inst.ft2232h_inst.rFifoStateZ0Z_2\ : std_logic;
signal \iRxF_n_c\ : std_logic;
signal \fifo_inst_ft2232h_inst_rFifoState_0\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c2\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.wRamWrEn_1\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rDataCount_axbxc1_0\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_1\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rDataCountZ0Z_2\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_0\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIJHQM1Z0Z_2_cascade_\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.wUartTxFull\ : std_logic;
signal \bfn_14_11_0_\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_0\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_1\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_2\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_3\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_4\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_5\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_6\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_7\ : std_logic;
signal \bfn_14_12_0_\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_7\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_5\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_6\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_4\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_5\ : std_logic;
signal \P1A7_c\ : std_logic;
signal \uart_inst0.uart_inst0.tx_state_81_d\ : std_logic;
signal \uart_inst0.uart_inst0.rTxDataZ0Z_0\ : std_logic;
signal \uart_inst0.uart_inst0.rTx_6_f1_0\ : std_logic;
signal \uart_inst0.uart_inst0.N_141_0\ : std_logic;
signal \uart_inst0.uart_inst0.N_143_0\ : std_logic;
signal \uart_inst0.uart_inst0.N_143_0_cascade_\ : std_logic;
signal \uart_inst0.uart_inst0.N_143_0_0\ : std_logic;
signal \uart_inst0.uart_inst0.un1_m3_0_a2_2_1\ : std_logic;
signal \uart_inst0.uart_inst0.N_136_0_cascade_\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_bits_remaining_c1\ : std_logic;
signal \uart_inst0.uart_inst0.N_136_0\ : std_logic;
signal \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_0\ : std_logic;
signal \wTxRdData_0\ : std_logic;
signal \INVfifo_inst.tx_fifo_inst.ram512x8_inst.RDATA_0C_net\ : std_logic;
signal \bfn_15_3_0_\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_0\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_1\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_2\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_3\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIMJ1QZ0\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_4\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIOM2QZ0\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_5\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIQP3QZ0\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_6\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_7\ : std_logic;
signal \bfn_15_4_0_\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIE7TPZ0\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNISS4QZ0\ : std_logic;
signal \fifo_inst_wRxWrEn\ : std_logic;
signal \bfn_15_5_0_\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_0\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNICK0CZ0\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_1\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_2\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_3\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_4\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIK05CZ0\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_5\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_6\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_7\ : std_logic;
signal \bfn_15_6_0_\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIIT3CZ0\ : std_logic;
signal \rTxEnZ0\ : std_logic;
signal \fifo_inst_wTxRdEn\ : std_logic;
signal \fifo_inst_tx_fifo_inst_rDataCount_0_sqmuxa\ : std_logic;
signal \fifo_inst_ft2232h_inst_rWrDelay\ : std_logic;
signal \fifo_inst_ft2232h_inst_rFifoState_4\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNIO67CZ0\ : std_logic;
signal \rUartTxDataZ0Z_6\ : std_logic;
signal \rUartTxDataZ0Z_5\ : std_logic;
signal \rUartTxDataZ0Z_1\ : std_logic;
signal \rUartRxDataZ0Z_5\ : std_logic;
signal \rUartRxDataZ0Z_6\ : std_logic;
signal \rUartRxDataZ0Z_1\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_2\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNISGZ0Z74\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_5_cascade_\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7_cascade_\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.wRamRdEn_1\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIBDOK2Z0Z_0\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7\ : std_logic;
signal \uart_inst0.wTxRdEn_0\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_5\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_6\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_7\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_0\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_3\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_4\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_3\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIUJZ0Z84\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_4\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_5\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNI2QAZ0Z4\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_6\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI4TBZ0Z4\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_7\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI60DZ0Z4\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_8\ : std_logic;
signal \uart_inst0.uart_inst0.rx_state_srsts_0_o2_3_3_cascade_\ : std_logic;
signal \uart_inst0.uart_inst0.N_257_0_cascade_\ : std_logic;
signal \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_2\ : std_logic;
signal \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_3\ : std_logic;
signal \uart_inst0.uart_inst0.N_157\ : std_logic;
signal \uart_inst0.uart_inst0.N_157_cascade_\ : std_logic;
signal \uart_inst0.uart_inst0.N_147_0_cascade_\ : std_logic;
signal \uart_inst0.uart_inst0.N_277_cascade_\ : std_logic;
signal \uart_inst0.uart_inst0.rx_state_srsts_0_a5_1_0\ : std_logic;
signal \uart_inst0.uart_inst0.N_280_cascade_\ : std_logic;
signal \uart_inst0.uart_inst0.rx_stateZ0Z_4\ : std_logic;
signal \uart_inst0.uart_inst0.N_261_0\ : std_logic;
signal \uart_inst0.wTxRdEmpty\ : std_logic;
signal \uart_inst0.uart_inst0.tx_state_ns_0_0_0_cascade_\ : std_logic;
signal \uart_inst0.uart_inst0.tx_state_1_sqmuxa_1_0_a3_0\ : std_logic;
signal \uart_inst0.uart_inst0.tx_state_RNI1319Z0Z_0\ : std_logic;
signal \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_1\ : std_logic;
signal \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_0\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_bits_remaining_ac0_1_a0_0_cascade_\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_bits_remaining_ac0_1\ : std_logic;
signal \uart_inst0.uart_inst0.un1_rx_state49_i_cascade_\ : std_logic;
signal \uart_inst0.uart_inst0.tx_countdown_RNO_0Z0Z_3_cascade_\ : std_logic;
signal \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_11_3_cascade_\ : std_logic;
signal \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13\ : std_logic;
signal \wTxFull\ : std_logic;
signal \rTxDataZ0Z_0\ : std_logic;
signal \rTxBusReady\ : std_logic;
signal \un1_rRamRdAddr_cry_2_c_RNIMVKN\ : std_logic;
signal m74 : std_logic;
signal \fifo_inst_tx_fifo_inst_rRamRdAddr_5\ : std_logic;
signal \fifo_inst_tx_fifo_inst_rRamRdAddr_7\ : std_logic;
signal \fifo_inst_tx_fifo_inst_rRamRdAddr_6\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.m72_eZ0Z_5_cascade_\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.N_100_cascade_\ : std_logic;
signal m73 : std_logic;
signal \fifo_inst_tx_fifo_inst_rRamRdAddr_3\ : std_logic;
signal \fifo_inst_tx_fifo_inst_rRamRdAddr_1\ : std_logic;
signal \fifo_inst_tx_fifo_inst_rRamRdAddr_8\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.m72_eZ0Z_6\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIKG0QZ0\ : std_logic;
signal \fifo_inst_tx_fifo_inst_rRamRdAddr_4\ : std_logic;
signal \fifo_inst_tx_fifo_inst_wRamRdEn\ : std_logic;
signal \rRamRdAddr_RNI9KL42_0\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.N_100\ : std_logic;
signal \fifo_inst_tx_fifo_inst_rRamRdAddr_0\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIM36CZ0\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIAHVBZ0\ : std_logic;
signal \un1_rRamRdAddr_cry_2_c_RNII9N9\ : std_logic;
signal m60 : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIGQ2CZ0\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rRamRdAddr_3\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rRamRdAddr_1\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rRamRdAddr_8\ : std_logic;
signal \N_101\ : std_logic;
signal \N_97\ : std_logic;
signal \iTxE_n_c\ : std_logic;
signal \N_8_0\ : std_logic;
signal \fifo_inst_ft2232h_inst_un1_rFifoState_1_sqmuxa_0_i_cascade_\ : std_logic;
signal \fifo_inst.ft2232h_inst.un1_rFifoState_1_sqmuxa_0_i_0\ : std_logic;
signal m59 : std_logic;
signal \fifo_inst_rx_fifo_inst_rRamRdAddr_5\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rRamRdAddr_4\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rRamRdAddr_2\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rRamRdAddr_7\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rRamRdAddr_6\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.m58_eZ0Z_5_cascade_\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.m58_eZ0Z_6\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.N_99\ : std_logic;
signal \rRamRdAddr_RNI0S8U_0\ : std_logic;
signal \fifo_inst_rx_fifo_inst_wRamRdEn\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.N_99_cascade_\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rRamRdAddr_0\ : std_logic;
signal \rUartRxDataZ0Z_3\ : std_logic;
signal \rUartTxDataZ0Z_3\ : std_logic;
signal \rUartRxDataZ0Z_4\ : std_logic;
signal \rRxDataZ0Z_4\ : std_logic;
signal \rUartTxDataZ0Z_4\ : std_logic;
signal \rUartRxDataZ0Z_7\ : std_logic;
signal \rUartTxDataZ0Z_7\ : std_logic;
signal \rUartRxDataZ0Z_2\ : std_logic;
signal \rUartTxDataZ0Z_2\ : std_logic;
signal \rUartRxDataZ0Z_0\ : std_logic;
signal \rUartRxFlagZ0\ : std_logic;
signal \rUartTxDataZ0Z_0\ : std_logic;
signal \rUartTxEn_4_0\ : std_logic;
signal \rUartRxState_0_0\ : std_logic;
signal \uart_inst0.uart_inst0.rx_stateZ0Z_0\ : std_logic;
signal \uart_inst0.wRxWrEn_0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_0_0\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ1Z_1\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ0Z_2\ : std_logic;
signal \uart_inst0.uart_inst0.rx_stateZ0Z_5\ : std_logic;
signal \uart_inst0.uart_inst0.N_283_cascade_\ : std_logic;
signal \uart_inst0.uart_inst0.rx_stateZ0Z_6\ : std_logic;
signal \uart_inst0.uart_inst0.rx_state_srsts_0_o2_3_3\ : std_logic;
signal \uart_inst0.uart_inst0.rx_countdown_2_sqmuxa_i_1\ : std_logic;
signal \uart_inst0.uart_inst0.un1_rx_clk_divider_0\ : std_logic;
signal \uart_inst0.uart_inst0.N_258_0_cascade_\ : std_logic;
signal \uart_inst0.uart_inst0.rx_countdownZ0Z_0\ : std_logic;
signal \bfn_16_15_0_\ : std_logic;
signal \uart_inst0.uart_inst0.rx_countdownZ0Z_1\ : std_logic;
signal \uart_inst0.uart_inst0.rx_countdown_s_1\ : std_logic;
signal \uart_inst0.uart_inst0.rx_countdown_cry_0\ : std_logic;
signal \uart_inst0.uart_inst0.rx_countdownZ0Z_2\ : std_logic;
signal \uart_inst0.uart_inst0.rx_countdown_s_2\ : std_logic;
signal \uart_inst0.uart_inst0.rx_countdown_cry_1\ : std_logic;
signal \uart_inst0.uart_inst0.rx_countdownZ0Z_3\ : std_logic;
signal \uart_inst0.uart_inst0.rx_countdown_s_3\ : std_logic;
signal \uart_inst0.uart_inst0.rx_countdown_cry_2\ : std_logic;
signal \uart_inst0.uart_inst0.rx_countdownZ0Z_4\ : std_logic;
signal \uart_inst0.uart_inst0.rx_countdown_cry_3_THRU_CO\ : std_logic;
signal \uart_inst0.uart_inst0.rx_countdown_cry_3\ : std_logic;
signal \uart_inst0.uart_inst0.N_252_0_i\ : std_logic;
signal \uart_inst0.uart_inst0.rx_countdown_cry_4\ : std_logic;
signal \uart_inst0.uart_inst0.rx_countdownZ0Z_5\ : std_logic;
signal \uart_inst0.uart_inst0.rx_countdowne_0_i\ : std_logic;
signal \uart_inst0.uart_inst0.N_258_0\ : std_logic;
signal \uart_inst0.uart_inst0.N_276_cascade_\ : std_logic;
signal \uart_inst0.uart_inst0.tx_stateZ0Z_0\ : std_logic;
signal \uart_inst0.uart_inst0.tx_stateZ0Z_1\ : std_logic;
signal \uart_inst0.uart_inst0.un1_m3_0_a2_0\ : std_logic;
signal \uart_inst0.uart_inst0.N_275\ : std_logic;
signal \uart_inst0.uart_inst0.N_147_0\ : std_logic;
signal \bfn_16_18_0_\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_0_s1_THRU_CO\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_0_s1\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_1_s1_THRU_CO\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_1_s1\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_2_s1\ : std_logic;
signal \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_4\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_3_s1_THRU_CO\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_3_s1\ : std_logic;
signal \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_5\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_4_s1_THRU_CO\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_4_s1\ : std_logic;
signal \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_6\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_5_s1_THRU_CO\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_5_s1\ : std_logic;
signal \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_7\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_6_s1_THRU_CO\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_6_s1\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_7_s1\ : std_logic;
signal \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_8\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_7_s1_THRU_CO\ : std_logic;
signal \bfn_16_19_0_\ : std_logic;
signal \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_9\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_8_s1_THRU_CO\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_8_s1\ : std_logic;
signal \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_10\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_9_s1_THRU_CO\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_9_s1\ : std_logic;
signal \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_11\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_10_s1_THRU_CO\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_10_s1\ : std_logic;
signal \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_12\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_11_s1_THRU_CO\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_11_s1\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_13\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_12_s1_THRU_CO\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_12_s1\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_13_s1\ : std_logic;
signal \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_14\ : std_logic;
signal \uart_inst0.uart_inst0.N_147_0_i_0\ : std_logic;
signal \bfn_17_2_0_\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_0\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_1\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_2\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_3\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_4\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_5\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_6\ : std_logic;
signal \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_7\ : std_logic;
signal \bfn_17_3_0_\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIGAUPZ0\ : std_logic;
signal \fifo_inst_tx_fifo_inst_rRamRdAddr_2\ : std_logic;
signal \fifo_inst_wRxWrFull\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rDataCount_2\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rDataCount_0\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rDataCount_1\ : std_logic;
signal \rRxDataZ0Z_6\ : std_logic;
signal \rRxDataZ0Z_1\ : std_logic;
signal \rRxDataZ0Z_2\ : std_logic;
signal \rRxDataZ0Z_3\ : std_logic;
signal \rRxDataZ0Z_0\ : std_logic;
signal \rRxDataZ0Z_5\ : std_logic;
signal \rRxDataZ0Z_7\ : std_logic;
signal \N_27_0\ : std_logic;
signal \bfn_17_6_0_\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_1\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_2\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_3\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_4\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_5\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_6\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_7\ : std_logic;
signal \bfn_17_7_0_\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNO_0_0_3\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNO_0_0_0\ : std_logic;
signal \wUartRxEmpty_cascade_\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.wRamWrEn\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rDataCount_RNI3V391Z0Z_2_cascade_\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rDataCount15_2_0_0_0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.wRamRdEn_cascade_\ : std_logic;
signal \rUartRxStateZ0Z_0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rDataCount_c2\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rDataCount_0_sqmuxa\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_2\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rDataCount_axbxc3_1_1\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_1\ : std_logic;
signal \uart_inst0.wRxWrFull_0\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIK0HSZ0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_1\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_2\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_3\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_4\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_5\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_6\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_7\ : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_1\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_2\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIOAZ0Z54\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_6\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_5\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_7\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_4\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_5\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_8\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_4\ : std_logic;
signal \wUartRxEmpty\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_3\ : std_logic;
signal \P1A1_c\ : std_logic;
signal \uart_inst0.uart_inst0.rx_stateZ0Z_1\ : std_logic;
signal \wPllLocked_i\ : std_logic;
signal \uart_inst0.uart_inst0.rRxData_0_sqmuxa\ : std_logic;
signal \wPllLocked\ : std_logic;
signal \uart_inst0.uart_inst0.N_257_0\ : std_logic;
signal \uart_inst0.uart_inst0.N_273_cascade_\ : std_logic;
signal \uart_inst0.uart_inst0.rx_stateZ0Z_3\ : std_logic;
signal \uart_inst0.uart_inst0.rx_state_srsts_0_a5_0_0_3\ : std_logic;
signal \uart_inst0.uart_inst0.N_274_2\ : std_logic;
signal \uart_inst0.uart_inst0.un1_rx_bits_remaining_c3_cascade_\ : std_logic;
signal \uart_inst0.uart_inst0.rx_bits_remainingZ0Z_3\ : std_logic;
signal \uart_inst0.uart_inst0.tx_countdownZ0Z_3\ : std_logic;
signal \uart_inst0.uart_inst0.tx_N_2\ : std_logic;
signal \uart_inst0.uart_inst0.tx_countdownZ0Z_2\ : std_logic;
signal \N_292_g\ : std_logic;
signal \uart_inst0.uart_inst0.N_147_0_i\ : std_logic;
signal \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_2_s1_THRU_CO\ : std_logic;
signal \uart_inst0.uart_inst0.un1_rx_state49_i\ : std_logic;
signal \uart_inst0.uart_inst0.tx_countdownZ0Z_1\ : std_logic;
signal \uart_inst0.uart_inst0.tx_countdownZ0Z_0\ : std_logic;
signal \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_9\ : std_logic;
signal \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_11_3\ : std_logic;
signal \uart_inst0.uart_inst0.tx_m5_0_2_cascade_\ : std_logic;
signal \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_11_4\ : std_logic;
signal \uart_inst0.uart_inst0.tx_N_11_mux\ : std_logic;
signal \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_2\ : std_logic;
signal \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_0\ : std_logic;
signal \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_3\ : std_logic;
signal \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_1\ : std_logic;
signal \uart_inst0.uart_inst0.tx_m5_0\ : std_logic;
signal \ioFifoData_in_5\ : std_logic;
signal \fifo_inst.wRxWrData_5\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rRamWrAddr_5\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rRamWrAddr_4\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rRamWrAddr_2\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rRamWrAddr_7\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rRamWrAddr_6\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.m54_eZ0Z_5_cascade_\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.N_91_cascade_\ : std_logic;
signal \un1_rRamWrAddr_cry_2_c_RNIOTMG\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rRamWrAddr_3\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rRamWrAddr_1\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rRamWrAddr_8\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.m54_eZ0Z_6\ : std_logic;
signal \rRamWrAddr_RNI9D19_0\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.N_91\ : std_logic;
signal \fifo_inst_rx_fifo_inst_wRamWrEn\ : std_logic;
signal \fifo_inst_rx_fifo_inst_rRamWrAddr_0\ : std_logic;
signal \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_4\ : std_logic;
signal \wRxData_4\ : std_logic;
signal \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_3\ : std_logic;
signal \wRxData_3\ : std_logic;
signal \INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_4C_net\ : std_logic;
signal \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_7\ : std_logic;
signal \wRxData_7\ : std_logic;
signal \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_5\ : std_logic;
signal \wRxData_5\ : std_logic;
signal \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_1\ : std_logic;
signal \wRxData_1\ : std_logic;
signal \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_2\ : std_logic;
signal \wRxData_2\ : std_logic;
signal \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_6\ : std_logic;
signal \wRxData_6\ : std_logic;
signal \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_0\ : std_logic;
signal \P1A2_c\ : std_logic;
signal \wRxData_0\ : std_logic;
signal \INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7C_net\ : std_logic;
signal \N_84_mux_i\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_8\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_3\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_2\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_1\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_0_cascade_\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_6\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_6\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_5\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_7\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_4\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_5\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_5\ : std_logic;
signal \wUartRxData_5\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_6\ : std_logic;
signal \wUartRxData_6\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_7\ : std_logic;
signal \rUartRxEnZ0\ : std_logic;
signal \wUartRxData_7\ : std_logic;
signal \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_5C_net\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.wUartRxEmpty_i\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_0\ : std_logic;
signal \wUartRxData_0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_1\ : std_logic;
signal \wUartRxData_1\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_2\ : std_logic;
signal \wUartRxData_2\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_3\ : std_logic;
signal \wUartRxData_3\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_4\ : std_logic;
signal \wUartRxData_4\ : std_logic;
signal \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIUFMSZ0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_5_0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIQ9KSZ0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_3_0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNID4JC2Z0Z_0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_8\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNISCLSZ0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_4_0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.wRamRdEn\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNIO6JSZ0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_2_0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI0JNSZ0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_6_0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIM3ISZ0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_1_0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI2MOSZ0\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_7_0\ : std_logic;
signal \uart_inst0.uart_inst0.un1_rx_bits_remaining_c1\ : std_logic;
signal \uart_inst0.uart_inst0.rx_bits_remaining_2_sqmuxa\ : std_logic;
signal \uart_inst0.uart_inst0.rx_bits_remainingZ0Z_2\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIQDZ0Z64\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_1\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNI0NZ0Z94\ : std_logic;
signal \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_4\ : std_logic;
signal \uart_inst0.wRxWrData_4\ : std_logic;
signal \uart_inst0.wRxWrData_1\ : std_logic;
signal \uart_inst0.wRxWrData_0\ : std_logic;
signal \uart_inst0.wRxWrData_5\ : std_logic;
signal \uart_inst0.wRxWrData_7\ : std_logic;
signal \uart_inst0.wRxWrData_6\ : std_logic;
signal \uart_inst0.wRxWrData_3\ : std_logic;
signal \uart_inst0.wRxWrData_2\ : std_logic;
signal \uart_inst0.uart_inst0.rRxData_0_sqmuxa_0\ : std_logic;
signal \uart_inst0.uart_inst0.rx_stateZ0Z_2\ : std_logic;
signal \uart_inst0.uart_inst0.rx_bits_remainingZ0Z_0\ : std_logic;
signal \uart_inst0.uart_inst0.N_283\ : std_logic;
signal \uart_inst0.uart_inst0.rx_bits_remainingZ0Z_1\ : std_logic;
signal \uart_inst0.uart_inst0.rx_state_2_sqmuxa\ : std_logic;
signal \ioFifoData_in_2\ : std_logic;
signal \fifo_inst.wRxWrData_2\ : std_logic;
signal \ioFifoData_in_1\ : std_logic;
signal \fifo_inst.wRxWrData_1\ : std_logic;
signal \ioFifoData_in_3\ : std_logic;
signal \fifo_inst.wRxWrData_3\ : std_logic;
signal \ioFifoData_in_4\ : std_logic;
signal \fifo_inst.wRxWrData_4\ : std_logic;
signal \ioFifoData_in_0\ : std_logic;
signal \fifo_inst.wRxWrData_0\ : std_logic;
signal \ioFifoData_in_7\ : std_logic;
signal \fifo_inst.wRxWrData_7\ : std_logic;
signal \ioFifoData_in_6\ : std_logic;
signal \fifo_inst.ft2232h_inst.rFifoStateZ0Z_1\ : std_logic;
signal \fifo_inst.wRxWrData_6\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_48mhz : std_logic;
signal \wPllLocked_i_g\ : std_logic;

signal \iClk_wire\ : std_logic;
signal \P1A8_wire\ : std_logic;
signal \P1A4_wire\ : std_logic;
signal \oRx_n_wire\ : std_logic;
signal \iRxF_n_wire\ : std_logic;
signal \P1A7_wire\ : std_logic;
signal \BTN_N_wire\ : std_logic;
signal \oTx_n_wire\ : std_logic;
signal \iTxE_n_wire\ : std_logic;
signal \P1A1_wire\ : std_logic;
signal \P1A9_wire\ : std_logic;
signal \P1A2_wire\ : std_logic;
signal \P1A3_wire\ : std_logic;
signal \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \top_pll_inst.top_pll_inst_pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \iClk_wire\ <= iClk;
    P1A8 <= \P1A8_wire\;
    P1A4 <= \P1A4_wire\;
    oRx_n <= \oRx_n_wire\;
    \iRxF_n_wire\ <= iRxF_n;
    P1A7 <= \P1A7_wire\;
    \BTN_N_wire\ <= BTN_N;
    oTx_n <= \oTx_n_wire\;
    \iTxE_n_wire\ <= iTxE_n;
    \P1A1_wire\ <= P1A1;
    P1A9 <= \P1A9_wire\;
    P1A2 <= \P1A2_wire\;
    P1A3 <= \P1A3_wire\;
    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_7\ <= \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(14);
    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_6\ <= \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(12);
    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_5\ <= \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(10);
    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_4\ <= \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(8);
    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_3\ <= \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(6);
    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_2\ <= \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(4);
    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_1\ <= \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(2);
    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_0\ <= \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(0);
    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&\N__15677\&\N__15719\&\N__15500\&\N__15434\&\N__15479\&\N__15740\&\N__15698\&\N__11093\&\N__15455\;
    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&\N__15290\&\N__15083\&\N__15137\&\N__15110\&\N__15053\&\N__15263\&\N__15236\&\N__15209\&\N__15179\;
    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WDATA_wire\ <= '0'&\N__16147\&'0'&\N__16118\&'0'&\N__16166\&'0'&\N__16211\&'0'&\N__16100\&'0'&\N__16082\&'0'&\N__16196\&'0'&\N__16178\;
    \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_7\ <= \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(14);
    \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_6\ <= \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(12);
    \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_5\ <= \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(10);
    \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_4\ <= \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(8);
    \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_3\ <= \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(6);
    \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_2\ <= \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(4);
    \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_1\ <= \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(2);
    \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_0\ <= \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(0);
    \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&\N__9137\&\N__10802\&\N__9008\&\N__9332\&\N__10733\&\N__10748\&\N__9041\&\N__10781\&\N__10460\;
    \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&\N__14138\&\N__14255\&\N__14228\&\N__14342\&\N__14315\&\N__14189\&\N__14288\&\N__14165\&\N__14804\;
    \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WDATA_wire\ <= '0'&\N__17095\&'0'&\N__17006\&'0'&\N__14360\&'0'&\N__17155\&'0'&\N__17186\&'0'&\N__15835\&'0'&\N__17210\&'0'&\N__17128\;
    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_7\ <= \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(14);
    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_6\ <= \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(12);
    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_5\ <= \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(10);
    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_4\ <= \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(8);
    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_3\ <= \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(6);
    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_2\ <= \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(4);
    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_1\ <= \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(2);
    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_0\ <= \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(0);
    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&\N__9428\&\N__9440\&\N__9452\&\N__15581\&\N__9737\&\N__9365\&\N__15605\&\N__13469\&\N__9551\;
    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&\N__7577\&\N__8747\&\N__8696\&\N__8723\&\N__8669\&\N__7352\&\N__7382\&\N__7409\&\N__7445\;
    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WDATA_wire\ <= '0'&\N__10838\&'0'&\N__9116\&'0'&\N__9104\&'0'&\N__10859\&'0'&\N__10892\&'0'&\N__10817\&'0'&\N__9092\&'0'&\N__11198\;
    \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_0\ <= \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\(0);
    \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&\N__8879\&\N__8927\&\N__8951\&\N__8975\&\N__10313\&\N__10433\&\N__12803\&\N__8900\&\N__10376\;
    \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&\N__7052\&\N__7082\&\N__7109\&\N__7142\&\N__6850\&\N__6890\&\N__6920\&\N__6947\&\N__6983\;
    \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__10106\;
    \top_pll_inst.top_pll_inst_pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__16965\,
            RE => \N__12278\,
            WCLKE => \N__13155\,
            WCLK => \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net\,
            WE => \N__12257\
        );

    \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__16985\,
            RE => \N__12313\,
            WCLKE => \N__14836\,
            WCLK => \INVfifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net\,
            WE => \N__12256\
        );

    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__16950\,
            RE => \N__12267\,
            WCLKE => \N__8510\,
            WCLK => \INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net\,
            WE => \N__12316\
        );

    \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__16990\,
            RE => \N__12314\,
            WCLKE => \N__7928\,
            WCLK => \INVfifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net\,
            WE => \N__12315\
        );

    \top_pll_inst.top_pll_inst_pll\ : PLL40
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "0111111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            PLLOUTGLOBAL => clk_48mhz,
            SDI => \GNDG0\,
            BYPASS => \GNDG0\,
            RESETB => \N__6461\,
            PLLOUTCORE => OPEN,
            LOCK => \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO\,
            SDO => OPEN,
            SCLK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            EXTFEEDBACK => \GNDG0\,
            DYNAMICDELAY => \top_pll_inst.top_pll_inst_pll_DYNAMICDELAY_wire\,
            PLLIN => \N__17429\
        );

    \top_pll_inst.top_pll_inst_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \VCCG0\,
            DIN => '0',
            DOUT => \N__17429\,
            PACKAGEPIN => \iClk_wire\
        );

    \P1A8_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17415\,
            DIN => \N__17414\,
            DOUT => \N__17413\,
            PACKAGEPIN => \P1A8_wire\
        );

    \P1A8_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__17415\,
            PADOUT => \N__17414\,
            PADIN => \N__17413\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A4_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17406\,
            DIN => \N__17405\,
            DOUT => \N__17404\,
            PACKAGEPIN => \P1A4_wire\
        );

    \P1A4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__17406\,
            PADOUT => \N__17405\,
            PADIN => \N__17404\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8014\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \oRx_n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17397\,
            DIN => \N__17396\,
            DOUT => \N__17395\,
            PACKAGEPIN => \oRx_n_wire\
        );

    \oRx_n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__17397\,
            PADOUT => \N__17396\,
            PADIN => \N__17395\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6820\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \iRxF_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17388\,
            DIN => \N__17387\,
            DOUT => \N__17386\,
            PACKAGEPIN => \iRxF_n_wire\
        );

    \iRxF_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__17388\,
            PADOUT => \N__17387\,
            PADIN => \N__17386\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \iRxF_n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A7_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17379\,
            DIN => \N__17378\,
            DOUT => \N__17377\,
            PACKAGEPIN => \P1A7_wire\
        );

    \P1A7_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__17379\,
            PADOUT => \N__17378\,
            PADIN => \N__17377\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8615\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17370\,
            DIN => \N__17369\,
            DOUT => \N__17368\,
            PACKAGEPIN => ioFifoData(7)
        );

    \ioFifoData_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__17370\,
            PADOUT => \N__17369\,
            PADIN => \N__17368\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10088\,
            DIN0 => \ioFifoData_in_7\,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BTN_N_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17361\,
            DIN => \N__17360\,
            DOUT => \N__17359\,
            PACKAGEPIN => \BTN_N_wire\
        );

    \BTN_N_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__17361\,
            PADOUT => \N__17360\,
            PADIN => \N__17359\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \BTN_N_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17352\,
            DIN => \N__17351\,
            DOUT => \N__17350\,
            PACKAGEPIN => ioFifoData(4)
        );

    \ioFifoData_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__17352\,
            PADOUT => \N__17351\,
            PADIN => \N__17350\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10056\,
            DIN0 => \ioFifoData_in_4\,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17343\,
            DIN => \N__17342\,
            DOUT => \N__17341\,
            PACKAGEPIN => ioFifoData(1)
        );

    \ioFifoData_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__17343\,
            PADOUT => \N__17342\,
            PADIN => \N__17341\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10055\,
            DIN0 => \ioFifoData_in_1\,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17334\,
            DIN => \N__17333\,
            DOUT => \N__17332\,
            PACKAGEPIN => ioFifoData(5)
        );

    \ioFifoData_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__17334\,
            PADOUT => \N__17333\,
            PADIN => \N__17332\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10057\,
            DIN0 => \ioFifoData_in_5\,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \oTx_n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17325\,
            DIN => \N__17324\,
            DOUT => \N__17323\,
            PACKAGEPIN => \oTx_n_wire\
        );

    \oTx_n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__17325\,
            PADOUT => \N__17324\,
            PADIN => \N__17323\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8021\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \iTxE_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17316\,
            DIN => \N__17315\,
            DOUT => \N__17314\,
            PACKAGEPIN => \iTxE_n_wire\
        );

    \iTxE_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__17316\,
            PADOUT => \N__17315\,
            PADIN => \N__17314\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \iTxE_n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17307\,
            DIN => \N__17306\,
            DOUT => \N__17305\,
            PACKAGEPIN => \P1A1_wire\
        );

    \P1A1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__17307\,
            PADOUT => \N__17306\,
            PADIN => \N__17305\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \P1A1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17298\,
            DIN => \N__17297\,
            DOUT => \N__17296\,
            PACKAGEPIN => ioFifoData(2)
        );

    \ioFifoData_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__17298\,
            PADOUT => \N__17297\,
            PADIN => \N__17296\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10075\,
            DIN0 => \ioFifoData_in_2\,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A9_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17289\,
            DIN => \N__17288\,
            DOUT => \N__17287\,
            PACKAGEPIN => \P1A9_wire\
        );

    \P1A9_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__17289\,
            PADOUT => \N__17288\,
            PADIN => \N__17287\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17280\,
            DIN => \N__17279\,
            DOUT => \N__17278\,
            PACKAGEPIN => ioFifoData(6)
        );

    \ioFifoData_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__17280\,
            PADOUT => \N__17279\,
            PADIN => \N__17278\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10087\,
            DIN0 => \ioFifoData_in_6\,
            DOUT0 => \N__12470\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17271\,
            DIN => \N__17270\,
            DOUT => \N__17269\,
            PACKAGEPIN => ioFifoData(3)
        );

    \ioFifoData_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__17271\,
            PADOUT => \N__17270\,
            PADIN => \N__17269\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10068\,
            DIN0 => \ioFifoData_in_3\,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17262\,
            DIN => \N__17261\,
            DOUT => \N__17260\,
            PACKAGEPIN => \P1A2_wire\
        );

    \P1A2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__17262\,
            PADOUT => \N__17261\,
            PADIN => \N__17260\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__15419\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17253\,
            DIN => \N__17252\,
            DOUT => \N__17251\,
            PACKAGEPIN => ioFifoData(0)
        );

    \ioFifoData_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__17253\,
            PADOUT => \N__17252\,
            PADIN => \N__17251\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10064\,
            DIN0 => \ioFifoData_in_0\,
            DOUT0 => \N__8846\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__17244\,
            DIN => \N__17243\,
            DOUT => \N__17242\,
            PACKAGEPIN => \P1A3_wire\
        );

    \P1A3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__17244\,
            PADOUT => \N__17243\,
            PADIN => \N__17242\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6821\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__4123\ : InMux
    port map (
            O => \N__17225\,
            I => \N__17222\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__17222\,
            I => \N__17219\
        );

    \I__4121\ : Span4Mux_h
    port map (
            O => \N__17219\,
            I => \N__17216\
        );

    \I__4120\ : IoSpan4Mux
    port map (
            O => \N__17216\,
            I => \N__17213\
        );

    \I__4119\ : Odrv4
    port map (
            O => \N__17213\,
            I => \ioFifoData_in_1\
        );

    \I__4118\ : InMux
    port map (
            O => \N__17210\,
            I => \N__17206\
        );

    \I__4117\ : InMux
    port map (
            O => \N__17209\,
            I => \N__17203\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__17206\,
            I => \N__17200\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__17203\,
            I => \fifo_inst.wRxWrData_1\
        );

    \I__4114\ : Odrv4
    port map (
            O => \N__17200\,
            I => \fifo_inst.wRxWrData_1\
        );

    \I__4113\ : InMux
    port map (
            O => \N__17195\,
            I => \N__17192\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__17192\,
            I => \N__17189\
        );

    \I__4111\ : Odrv4
    port map (
            O => \N__17189\,
            I => \ioFifoData_in_3\
        );

    \I__4110\ : InMux
    port map (
            O => \N__17186\,
            I => \N__17183\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__17183\,
            I => \N__17179\
        );

    \I__4108\ : InMux
    port map (
            O => \N__17182\,
            I => \N__17176\
        );

    \I__4107\ : Span4Mux_h
    port map (
            O => \N__17179\,
            I => \N__17173\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__17176\,
            I => \fifo_inst.wRxWrData_3\
        );

    \I__4105\ : Odrv4
    port map (
            O => \N__17173\,
            I => \fifo_inst.wRxWrData_3\
        );

    \I__4104\ : InMux
    port map (
            O => \N__17168\,
            I => \N__17165\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__17165\,
            I => \N__17162\
        );

    \I__4102\ : IoSpan4Mux
    port map (
            O => \N__17162\,
            I => \N__17159\
        );

    \I__4101\ : Odrv4
    port map (
            O => \N__17159\,
            I => \ioFifoData_in_4\
        );

    \I__4100\ : InMux
    port map (
            O => \N__17156\,
            I => \N__17152\
        );

    \I__4099\ : InMux
    port map (
            O => \N__17155\,
            I => \N__17149\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__17152\,
            I => \fifo_inst.wRxWrData_4\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__17149\,
            I => \fifo_inst.wRxWrData_4\
        );

    \I__4096\ : InMux
    port map (
            O => \N__17144\,
            I => \N__17141\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__17141\,
            I => \N__17138\
        );

    \I__4094\ : Sp12to4
    port map (
            O => \N__17138\,
            I => \N__17135\
        );

    \I__4093\ : Span12Mux_h
    port map (
            O => \N__17135\,
            I => \N__17132\
        );

    \I__4092\ : Odrv12
    port map (
            O => \N__17132\,
            I => \ioFifoData_in_0\
        );

    \I__4091\ : InMux
    port map (
            O => \N__17129\,
            I => \N__17125\
        );

    \I__4090\ : InMux
    port map (
            O => \N__17128\,
            I => \N__17122\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__17125\,
            I => \fifo_inst.wRxWrData_0\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__17122\,
            I => \fifo_inst.wRxWrData_0\
        );

    \I__4087\ : InMux
    port map (
            O => \N__17117\,
            I => \N__17114\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__17114\,
            I => \N__17111\
        );

    \I__4085\ : Span4Mux_h
    port map (
            O => \N__17111\,
            I => \N__17108\
        );

    \I__4084\ : Sp12to4
    port map (
            O => \N__17108\,
            I => \N__17105\
        );

    \I__4083\ : Span12Mux_v
    port map (
            O => \N__17105\,
            I => \N__17102\
        );

    \I__4082\ : Span12Mux_v
    port map (
            O => \N__17102\,
            I => \N__17099\
        );

    \I__4081\ : Odrv12
    port map (
            O => \N__17099\,
            I => \ioFifoData_in_7\
        );

    \I__4080\ : InMux
    port map (
            O => \N__17096\,
            I => \N__17092\
        );

    \I__4079\ : InMux
    port map (
            O => \N__17095\,
            I => \N__17089\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__17092\,
            I => \fifo_inst.wRxWrData_7\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__17089\,
            I => \fifo_inst.wRxWrData_7\
        );

    \I__4076\ : InMux
    port map (
            O => \N__17084\,
            I => \N__17081\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__17081\,
            I => \N__17078\
        );

    \I__4074\ : Span4Mux_v
    port map (
            O => \N__17078\,
            I => \N__17075\
        );

    \I__4073\ : Sp12to4
    port map (
            O => \N__17075\,
            I => \N__17072\
        );

    \I__4072\ : Span12Mux_s6_h
    port map (
            O => \N__17072\,
            I => \N__17069\
        );

    \I__4071\ : Span12Mux_v
    port map (
            O => \N__17069\,
            I => \N__17066\
        );

    \I__4070\ : Odrv12
    port map (
            O => \N__17066\,
            I => \ioFifoData_in_6\
        );

    \I__4069\ : InMux
    port map (
            O => \N__17063\,
            I => \N__17044\
        );

    \I__4068\ : InMux
    port map (
            O => \N__17062\,
            I => \N__17044\
        );

    \I__4067\ : InMux
    port map (
            O => \N__17061\,
            I => \N__17044\
        );

    \I__4066\ : InMux
    port map (
            O => \N__17060\,
            I => \N__17044\
        );

    \I__4065\ : InMux
    port map (
            O => \N__17059\,
            I => \N__17044\
        );

    \I__4064\ : InMux
    port map (
            O => \N__17058\,
            I => \N__17044\
        );

    \I__4063\ : InMux
    port map (
            O => \N__17057\,
            I => \N__17041\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__17044\,
            I => \N__17035\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__17041\,
            I => \N__17035\
        );

    \I__4060\ : InMux
    port map (
            O => \N__17040\,
            I => \N__17032\
        );

    \I__4059\ : Span4Mux_v
    port map (
            O => \N__17035\,
            I => \N__17029\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__17032\,
            I => \N__17022\
        );

    \I__4057\ : Sp12to4
    port map (
            O => \N__17029\,
            I => \N__17022\
        );

    \I__4056\ : InMux
    port map (
            O => \N__17028\,
            I => \N__17019\
        );

    \I__4055\ : InMux
    port map (
            O => \N__17027\,
            I => \N__17016\
        );

    \I__4054\ : Span12Mux_s11_h
    port map (
            O => \N__17022\,
            I => \N__17011\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__17019\,
            I => \N__17011\
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__17016\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_1\
        );

    \I__4051\ : Odrv12
    port map (
            O => \N__17011\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_1\
        );

    \I__4050\ : InMux
    port map (
            O => \N__17006\,
            I => \N__17002\
        );

    \I__4049\ : InMux
    port map (
            O => \N__17005\,
            I => \N__16999\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__17002\,
            I => \N__16996\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__16999\,
            I => \fifo_inst.wRxWrData_6\
        );

    \I__4046\ : Odrv4
    port map (
            O => \N__16996\,
            I => \fifo_inst.wRxWrData_6\
        );

    \I__4045\ : ClkMux
    port map (
            O => \N__16991\,
            I => \N__16706\
        );

    \I__4044\ : ClkMux
    port map (
            O => \N__16990\,
            I => \N__16706\
        );

    \I__4043\ : ClkMux
    port map (
            O => \N__16989\,
            I => \N__16706\
        );

    \I__4042\ : ClkMux
    port map (
            O => \N__16988\,
            I => \N__16706\
        );

    \I__4041\ : ClkMux
    port map (
            O => \N__16987\,
            I => \N__16706\
        );

    \I__4040\ : ClkMux
    port map (
            O => \N__16986\,
            I => \N__16706\
        );

    \I__4039\ : ClkMux
    port map (
            O => \N__16985\,
            I => \N__16706\
        );

    \I__4038\ : ClkMux
    port map (
            O => \N__16984\,
            I => \N__16706\
        );

    \I__4037\ : ClkMux
    port map (
            O => \N__16983\,
            I => \N__16706\
        );

    \I__4036\ : ClkMux
    port map (
            O => \N__16982\,
            I => \N__16706\
        );

    \I__4035\ : ClkMux
    port map (
            O => \N__16981\,
            I => \N__16706\
        );

    \I__4034\ : ClkMux
    port map (
            O => \N__16980\,
            I => \N__16706\
        );

    \I__4033\ : ClkMux
    port map (
            O => \N__16979\,
            I => \N__16706\
        );

    \I__4032\ : ClkMux
    port map (
            O => \N__16978\,
            I => \N__16706\
        );

    \I__4031\ : ClkMux
    port map (
            O => \N__16977\,
            I => \N__16706\
        );

    \I__4030\ : ClkMux
    port map (
            O => \N__16976\,
            I => \N__16706\
        );

    \I__4029\ : ClkMux
    port map (
            O => \N__16975\,
            I => \N__16706\
        );

    \I__4028\ : ClkMux
    port map (
            O => \N__16974\,
            I => \N__16706\
        );

    \I__4027\ : ClkMux
    port map (
            O => \N__16973\,
            I => \N__16706\
        );

    \I__4026\ : ClkMux
    port map (
            O => \N__16972\,
            I => \N__16706\
        );

    \I__4025\ : ClkMux
    port map (
            O => \N__16971\,
            I => \N__16706\
        );

    \I__4024\ : ClkMux
    port map (
            O => \N__16970\,
            I => \N__16706\
        );

    \I__4023\ : ClkMux
    port map (
            O => \N__16969\,
            I => \N__16706\
        );

    \I__4022\ : ClkMux
    port map (
            O => \N__16968\,
            I => \N__16706\
        );

    \I__4021\ : ClkMux
    port map (
            O => \N__16967\,
            I => \N__16706\
        );

    \I__4020\ : ClkMux
    port map (
            O => \N__16966\,
            I => \N__16706\
        );

    \I__4019\ : ClkMux
    port map (
            O => \N__16965\,
            I => \N__16706\
        );

    \I__4018\ : ClkMux
    port map (
            O => \N__16964\,
            I => \N__16706\
        );

    \I__4017\ : ClkMux
    port map (
            O => \N__16963\,
            I => \N__16706\
        );

    \I__4016\ : ClkMux
    port map (
            O => \N__16962\,
            I => \N__16706\
        );

    \I__4015\ : ClkMux
    port map (
            O => \N__16961\,
            I => \N__16706\
        );

    \I__4014\ : ClkMux
    port map (
            O => \N__16960\,
            I => \N__16706\
        );

    \I__4013\ : ClkMux
    port map (
            O => \N__16959\,
            I => \N__16706\
        );

    \I__4012\ : ClkMux
    port map (
            O => \N__16958\,
            I => \N__16706\
        );

    \I__4011\ : ClkMux
    port map (
            O => \N__16957\,
            I => \N__16706\
        );

    \I__4010\ : ClkMux
    port map (
            O => \N__16956\,
            I => \N__16706\
        );

    \I__4009\ : ClkMux
    port map (
            O => \N__16955\,
            I => \N__16706\
        );

    \I__4008\ : ClkMux
    port map (
            O => \N__16954\,
            I => \N__16706\
        );

    \I__4007\ : ClkMux
    port map (
            O => \N__16953\,
            I => \N__16706\
        );

    \I__4006\ : ClkMux
    port map (
            O => \N__16952\,
            I => \N__16706\
        );

    \I__4005\ : ClkMux
    port map (
            O => \N__16951\,
            I => \N__16706\
        );

    \I__4004\ : ClkMux
    port map (
            O => \N__16950\,
            I => \N__16706\
        );

    \I__4003\ : ClkMux
    port map (
            O => \N__16949\,
            I => \N__16706\
        );

    \I__4002\ : ClkMux
    port map (
            O => \N__16948\,
            I => \N__16706\
        );

    \I__4001\ : ClkMux
    port map (
            O => \N__16947\,
            I => \N__16706\
        );

    \I__4000\ : ClkMux
    port map (
            O => \N__16946\,
            I => \N__16706\
        );

    \I__3999\ : ClkMux
    port map (
            O => \N__16945\,
            I => \N__16706\
        );

    \I__3998\ : ClkMux
    port map (
            O => \N__16944\,
            I => \N__16706\
        );

    \I__3997\ : ClkMux
    port map (
            O => \N__16943\,
            I => \N__16706\
        );

    \I__3996\ : ClkMux
    port map (
            O => \N__16942\,
            I => \N__16706\
        );

    \I__3995\ : ClkMux
    port map (
            O => \N__16941\,
            I => \N__16706\
        );

    \I__3994\ : ClkMux
    port map (
            O => \N__16940\,
            I => \N__16706\
        );

    \I__3993\ : ClkMux
    port map (
            O => \N__16939\,
            I => \N__16706\
        );

    \I__3992\ : ClkMux
    port map (
            O => \N__16938\,
            I => \N__16706\
        );

    \I__3991\ : ClkMux
    port map (
            O => \N__16937\,
            I => \N__16706\
        );

    \I__3990\ : ClkMux
    port map (
            O => \N__16936\,
            I => \N__16706\
        );

    \I__3989\ : ClkMux
    port map (
            O => \N__16935\,
            I => \N__16706\
        );

    \I__3988\ : ClkMux
    port map (
            O => \N__16934\,
            I => \N__16706\
        );

    \I__3987\ : ClkMux
    port map (
            O => \N__16933\,
            I => \N__16706\
        );

    \I__3986\ : ClkMux
    port map (
            O => \N__16932\,
            I => \N__16706\
        );

    \I__3985\ : ClkMux
    port map (
            O => \N__16931\,
            I => \N__16706\
        );

    \I__3984\ : ClkMux
    port map (
            O => \N__16930\,
            I => \N__16706\
        );

    \I__3983\ : ClkMux
    port map (
            O => \N__16929\,
            I => \N__16706\
        );

    \I__3982\ : ClkMux
    port map (
            O => \N__16928\,
            I => \N__16706\
        );

    \I__3981\ : ClkMux
    port map (
            O => \N__16927\,
            I => \N__16706\
        );

    \I__3980\ : ClkMux
    port map (
            O => \N__16926\,
            I => \N__16706\
        );

    \I__3979\ : ClkMux
    port map (
            O => \N__16925\,
            I => \N__16706\
        );

    \I__3978\ : ClkMux
    port map (
            O => \N__16924\,
            I => \N__16706\
        );

    \I__3977\ : ClkMux
    port map (
            O => \N__16923\,
            I => \N__16706\
        );

    \I__3976\ : ClkMux
    port map (
            O => \N__16922\,
            I => \N__16706\
        );

    \I__3975\ : ClkMux
    port map (
            O => \N__16921\,
            I => \N__16706\
        );

    \I__3974\ : ClkMux
    port map (
            O => \N__16920\,
            I => \N__16706\
        );

    \I__3973\ : ClkMux
    port map (
            O => \N__16919\,
            I => \N__16706\
        );

    \I__3972\ : ClkMux
    port map (
            O => \N__16918\,
            I => \N__16706\
        );

    \I__3971\ : ClkMux
    port map (
            O => \N__16917\,
            I => \N__16706\
        );

    \I__3970\ : ClkMux
    port map (
            O => \N__16916\,
            I => \N__16706\
        );

    \I__3969\ : ClkMux
    port map (
            O => \N__16915\,
            I => \N__16706\
        );

    \I__3968\ : ClkMux
    port map (
            O => \N__16914\,
            I => \N__16706\
        );

    \I__3967\ : ClkMux
    port map (
            O => \N__16913\,
            I => \N__16706\
        );

    \I__3966\ : ClkMux
    port map (
            O => \N__16912\,
            I => \N__16706\
        );

    \I__3965\ : ClkMux
    port map (
            O => \N__16911\,
            I => \N__16706\
        );

    \I__3964\ : ClkMux
    port map (
            O => \N__16910\,
            I => \N__16706\
        );

    \I__3963\ : ClkMux
    port map (
            O => \N__16909\,
            I => \N__16706\
        );

    \I__3962\ : ClkMux
    port map (
            O => \N__16908\,
            I => \N__16706\
        );

    \I__3961\ : ClkMux
    port map (
            O => \N__16907\,
            I => \N__16706\
        );

    \I__3960\ : ClkMux
    port map (
            O => \N__16906\,
            I => \N__16706\
        );

    \I__3959\ : ClkMux
    port map (
            O => \N__16905\,
            I => \N__16706\
        );

    \I__3958\ : ClkMux
    port map (
            O => \N__16904\,
            I => \N__16706\
        );

    \I__3957\ : ClkMux
    port map (
            O => \N__16903\,
            I => \N__16706\
        );

    \I__3956\ : ClkMux
    port map (
            O => \N__16902\,
            I => \N__16706\
        );

    \I__3955\ : ClkMux
    port map (
            O => \N__16901\,
            I => \N__16706\
        );

    \I__3954\ : ClkMux
    port map (
            O => \N__16900\,
            I => \N__16706\
        );

    \I__3953\ : ClkMux
    port map (
            O => \N__16899\,
            I => \N__16706\
        );

    \I__3952\ : ClkMux
    port map (
            O => \N__16898\,
            I => \N__16706\
        );

    \I__3951\ : ClkMux
    port map (
            O => \N__16897\,
            I => \N__16706\
        );

    \I__3950\ : GlobalMux
    port map (
            O => \N__16706\,
            I => clk_48mhz
        );

    \I__3949\ : CascadeMux
    port map (
            O => \N__16703\,
            I => \N__16690\
        );

    \I__3948\ : CascadeMux
    port map (
            O => \N__16702\,
            I => \N__16671\
        );

    \I__3947\ : CascadeMux
    port map (
            O => \N__16701\,
            I => \N__16667\
        );

    \I__3946\ : CascadeMux
    port map (
            O => \N__16700\,
            I => \N__16654\
        );

    \I__3945\ : CascadeMux
    port map (
            O => \N__16699\,
            I => \N__16650\
        );

    \I__3944\ : CascadeMux
    port map (
            O => \N__16698\,
            I => \N__16646\
        );

    \I__3943\ : CascadeMux
    port map (
            O => \N__16697\,
            I => \N__16641\
        );

    \I__3942\ : InMux
    port map (
            O => \N__16696\,
            I => \N__16615\
        );

    \I__3941\ : InMux
    port map (
            O => \N__16695\,
            I => \N__16610\
        );

    \I__3940\ : InMux
    port map (
            O => \N__16694\,
            I => \N__16610\
        );

    \I__3939\ : InMux
    port map (
            O => \N__16693\,
            I => \N__16607\
        );

    \I__3938\ : InMux
    port map (
            O => \N__16690\,
            I => \N__16594\
        );

    \I__3937\ : InMux
    port map (
            O => \N__16689\,
            I => \N__16594\
        );

    \I__3936\ : InMux
    port map (
            O => \N__16688\,
            I => \N__16594\
        );

    \I__3935\ : InMux
    port map (
            O => \N__16687\,
            I => \N__16594\
        );

    \I__3934\ : InMux
    port map (
            O => \N__16686\,
            I => \N__16594\
        );

    \I__3933\ : InMux
    port map (
            O => \N__16685\,
            I => \N__16594\
        );

    \I__3932\ : InMux
    port map (
            O => \N__16684\,
            I => \N__16589\
        );

    \I__3931\ : InMux
    port map (
            O => \N__16683\,
            I => \N__16589\
        );

    \I__3930\ : InMux
    port map (
            O => \N__16682\,
            I => \N__16580\
        );

    \I__3929\ : InMux
    port map (
            O => \N__16681\,
            I => \N__16580\
        );

    \I__3928\ : InMux
    port map (
            O => \N__16680\,
            I => \N__16580\
        );

    \I__3927\ : InMux
    port map (
            O => \N__16679\,
            I => \N__16580\
        );

    \I__3926\ : InMux
    port map (
            O => \N__16678\,
            I => \N__16577\
        );

    \I__3925\ : InMux
    port map (
            O => \N__16677\,
            I => \N__16572\
        );

    \I__3924\ : InMux
    port map (
            O => \N__16676\,
            I => \N__16572\
        );

    \I__3923\ : InMux
    port map (
            O => \N__16675\,
            I => \N__16569\
        );

    \I__3922\ : InMux
    port map (
            O => \N__16674\,
            I => \N__16566\
        );

    \I__3921\ : InMux
    port map (
            O => \N__16671\,
            I => \N__16563\
        );

    \I__3920\ : InMux
    port map (
            O => \N__16670\,
            I => \N__16560\
        );

    \I__3919\ : InMux
    port map (
            O => \N__16667\,
            I => \N__16555\
        );

    \I__3918\ : InMux
    port map (
            O => \N__16666\,
            I => \N__16555\
        );

    \I__3917\ : InMux
    port map (
            O => \N__16665\,
            I => \N__16548\
        );

    \I__3916\ : InMux
    port map (
            O => \N__16664\,
            I => \N__16548\
        );

    \I__3915\ : InMux
    port map (
            O => \N__16663\,
            I => \N__16548\
        );

    \I__3914\ : InMux
    port map (
            O => \N__16662\,
            I => \N__16541\
        );

    \I__3913\ : InMux
    port map (
            O => \N__16661\,
            I => \N__16541\
        );

    \I__3912\ : InMux
    port map (
            O => \N__16660\,
            I => \N__16541\
        );

    \I__3911\ : InMux
    port map (
            O => \N__16659\,
            I => \N__16538\
        );

    \I__3910\ : InMux
    port map (
            O => \N__16658\,
            I => \N__16531\
        );

    \I__3909\ : InMux
    port map (
            O => \N__16657\,
            I => \N__16531\
        );

    \I__3908\ : InMux
    port map (
            O => \N__16654\,
            I => \N__16531\
        );

    \I__3907\ : InMux
    port map (
            O => \N__16653\,
            I => \N__16526\
        );

    \I__3906\ : InMux
    port map (
            O => \N__16650\,
            I => \N__16526\
        );

    \I__3905\ : InMux
    port map (
            O => \N__16649\,
            I => \N__16523\
        );

    \I__3904\ : InMux
    port map (
            O => \N__16646\,
            I => \N__16518\
        );

    \I__3903\ : InMux
    port map (
            O => \N__16645\,
            I => \N__16518\
        );

    \I__3902\ : InMux
    port map (
            O => \N__16644\,
            I => \N__16511\
        );

    \I__3901\ : InMux
    port map (
            O => \N__16641\,
            I => \N__16511\
        );

    \I__3900\ : InMux
    port map (
            O => \N__16640\,
            I => \N__16511\
        );

    \I__3899\ : InMux
    port map (
            O => \N__16639\,
            I => \N__16504\
        );

    \I__3898\ : InMux
    port map (
            O => \N__16638\,
            I => \N__16504\
        );

    \I__3897\ : InMux
    port map (
            O => \N__16637\,
            I => \N__16504\
        );

    \I__3896\ : InMux
    port map (
            O => \N__16636\,
            I => \N__16497\
        );

    \I__3895\ : InMux
    port map (
            O => \N__16635\,
            I => \N__16497\
        );

    \I__3894\ : InMux
    port map (
            O => \N__16634\,
            I => \N__16497\
        );

    \I__3893\ : InMux
    port map (
            O => \N__16633\,
            I => \N__16490\
        );

    \I__3892\ : InMux
    port map (
            O => \N__16632\,
            I => \N__16490\
        );

    \I__3891\ : InMux
    port map (
            O => \N__16631\,
            I => \N__16490\
        );

    \I__3890\ : InMux
    port map (
            O => \N__16630\,
            I => \N__16483\
        );

    \I__3889\ : InMux
    port map (
            O => \N__16629\,
            I => \N__16483\
        );

    \I__3888\ : InMux
    port map (
            O => \N__16628\,
            I => \N__16483\
        );

    \I__3887\ : InMux
    port map (
            O => \N__16627\,
            I => \N__16480\
        );

    \I__3886\ : InMux
    port map (
            O => \N__16626\,
            I => \N__16473\
        );

    \I__3885\ : InMux
    port map (
            O => \N__16625\,
            I => \N__16473\
        );

    \I__3884\ : InMux
    port map (
            O => \N__16624\,
            I => \N__16473\
        );

    \I__3883\ : InMux
    port map (
            O => \N__16623\,
            I => \N__16466\
        );

    \I__3882\ : InMux
    port map (
            O => \N__16622\,
            I => \N__16466\
        );

    \I__3881\ : InMux
    port map (
            O => \N__16621\,
            I => \N__16466\
        );

    \I__3880\ : InMux
    port map (
            O => \N__16620\,
            I => \N__16459\
        );

    \I__3879\ : InMux
    port map (
            O => \N__16619\,
            I => \N__16459\
        );

    \I__3878\ : InMux
    port map (
            O => \N__16618\,
            I => \N__16459\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__16615\,
            I => \N__16456\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__16610\,
            I => \N__16450\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__16607\,
            I => \N__16445\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__16594\,
            I => \N__16442\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__16589\,
            I => \N__16439\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__16580\,
            I => \N__16433\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__16577\,
            I => \N__16430\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__16572\,
            I => \N__16426\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__16569\,
            I => \N__16422\
        );

    \I__3868\ : LocalMux
    port map (
            O => \N__16566\,
            I => \N__16410\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__16563\,
            I => \N__16407\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__16560\,
            I => \N__16404\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__16555\,
            I => \N__16401\
        );

    \I__3864\ : LocalMux
    port map (
            O => \N__16548\,
            I => \N__16398\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__16541\,
            I => \N__16395\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__16538\,
            I => \N__16392\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__16531\,
            I => \N__16389\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__16526\,
            I => \N__16386\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__16523\,
            I => \N__16381\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__16518\,
            I => \N__16378\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__16511\,
            I => \N__16375\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__16504\,
            I => \N__16372\
        );

    \I__3855\ : LocalMux
    port map (
            O => \N__16497\,
            I => \N__16369\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__16490\,
            I => \N__16363\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__16483\,
            I => \N__16360\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__16480\,
            I => \N__16352\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__16473\,
            I => \N__16347\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__16466\,
            I => \N__16344\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__16459\,
            I => \N__16341\
        );

    \I__3848\ : Glb2LocalMux
    port map (
            O => \N__16456\,
            I => \N__16217\
        );

    \I__3847\ : SRMux
    port map (
            O => \N__16455\,
            I => \N__16217\
        );

    \I__3846\ : SRMux
    port map (
            O => \N__16454\,
            I => \N__16217\
        );

    \I__3845\ : SRMux
    port map (
            O => \N__16453\,
            I => \N__16217\
        );

    \I__3844\ : Glb2LocalMux
    port map (
            O => \N__16450\,
            I => \N__16217\
        );

    \I__3843\ : SRMux
    port map (
            O => \N__16449\,
            I => \N__16217\
        );

    \I__3842\ : SRMux
    port map (
            O => \N__16448\,
            I => \N__16217\
        );

    \I__3841\ : Glb2LocalMux
    port map (
            O => \N__16445\,
            I => \N__16217\
        );

    \I__3840\ : Glb2LocalMux
    port map (
            O => \N__16442\,
            I => \N__16217\
        );

    \I__3839\ : Glb2LocalMux
    port map (
            O => \N__16439\,
            I => \N__16217\
        );

    \I__3838\ : SRMux
    port map (
            O => \N__16438\,
            I => \N__16217\
        );

    \I__3837\ : SRMux
    port map (
            O => \N__16437\,
            I => \N__16217\
        );

    \I__3836\ : SRMux
    port map (
            O => \N__16436\,
            I => \N__16217\
        );

    \I__3835\ : Glb2LocalMux
    port map (
            O => \N__16433\,
            I => \N__16217\
        );

    \I__3834\ : Glb2LocalMux
    port map (
            O => \N__16430\,
            I => \N__16217\
        );

    \I__3833\ : SRMux
    port map (
            O => \N__16429\,
            I => \N__16217\
        );

    \I__3832\ : Glb2LocalMux
    port map (
            O => \N__16426\,
            I => \N__16217\
        );

    \I__3831\ : SRMux
    port map (
            O => \N__16425\,
            I => \N__16217\
        );

    \I__3830\ : Glb2LocalMux
    port map (
            O => \N__16422\,
            I => \N__16217\
        );

    \I__3829\ : SRMux
    port map (
            O => \N__16421\,
            I => \N__16217\
        );

    \I__3828\ : SRMux
    port map (
            O => \N__16420\,
            I => \N__16217\
        );

    \I__3827\ : SRMux
    port map (
            O => \N__16419\,
            I => \N__16217\
        );

    \I__3826\ : SRMux
    port map (
            O => \N__16418\,
            I => \N__16217\
        );

    \I__3825\ : SRMux
    port map (
            O => \N__16417\,
            I => \N__16217\
        );

    \I__3824\ : SRMux
    port map (
            O => \N__16416\,
            I => \N__16217\
        );

    \I__3823\ : SRMux
    port map (
            O => \N__16415\,
            I => \N__16217\
        );

    \I__3822\ : SRMux
    port map (
            O => \N__16414\,
            I => \N__16217\
        );

    \I__3821\ : SRMux
    port map (
            O => \N__16413\,
            I => \N__16217\
        );

    \I__3820\ : Glb2LocalMux
    port map (
            O => \N__16410\,
            I => \N__16217\
        );

    \I__3819\ : Glb2LocalMux
    port map (
            O => \N__16407\,
            I => \N__16217\
        );

    \I__3818\ : Glb2LocalMux
    port map (
            O => \N__16404\,
            I => \N__16217\
        );

    \I__3817\ : Glb2LocalMux
    port map (
            O => \N__16401\,
            I => \N__16217\
        );

    \I__3816\ : Glb2LocalMux
    port map (
            O => \N__16398\,
            I => \N__16217\
        );

    \I__3815\ : Glb2LocalMux
    port map (
            O => \N__16395\,
            I => \N__16217\
        );

    \I__3814\ : Glb2LocalMux
    port map (
            O => \N__16392\,
            I => \N__16217\
        );

    \I__3813\ : Glb2LocalMux
    port map (
            O => \N__16389\,
            I => \N__16217\
        );

    \I__3812\ : Glb2LocalMux
    port map (
            O => \N__16386\,
            I => \N__16217\
        );

    \I__3811\ : SRMux
    port map (
            O => \N__16385\,
            I => \N__16217\
        );

    \I__3810\ : SRMux
    port map (
            O => \N__16384\,
            I => \N__16217\
        );

    \I__3809\ : Glb2LocalMux
    port map (
            O => \N__16381\,
            I => \N__16217\
        );

    \I__3808\ : Glb2LocalMux
    port map (
            O => \N__16378\,
            I => \N__16217\
        );

    \I__3807\ : Glb2LocalMux
    port map (
            O => \N__16375\,
            I => \N__16217\
        );

    \I__3806\ : Glb2LocalMux
    port map (
            O => \N__16372\,
            I => \N__16217\
        );

    \I__3805\ : Glb2LocalMux
    port map (
            O => \N__16369\,
            I => \N__16217\
        );

    \I__3804\ : SRMux
    port map (
            O => \N__16368\,
            I => \N__16217\
        );

    \I__3803\ : SRMux
    port map (
            O => \N__16367\,
            I => \N__16217\
        );

    \I__3802\ : SRMux
    port map (
            O => \N__16366\,
            I => \N__16217\
        );

    \I__3801\ : Glb2LocalMux
    port map (
            O => \N__16363\,
            I => \N__16217\
        );

    \I__3800\ : Glb2LocalMux
    port map (
            O => \N__16360\,
            I => \N__16217\
        );

    \I__3799\ : SRMux
    port map (
            O => \N__16359\,
            I => \N__16217\
        );

    \I__3798\ : SRMux
    port map (
            O => \N__16358\,
            I => \N__16217\
        );

    \I__3797\ : SRMux
    port map (
            O => \N__16357\,
            I => \N__16217\
        );

    \I__3796\ : SRMux
    port map (
            O => \N__16356\,
            I => \N__16217\
        );

    \I__3795\ : SRMux
    port map (
            O => \N__16355\,
            I => \N__16217\
        );

    \I__3794\ : Glb2LocalMux
    port map (
            O => \N__16352\,
            I => \N__16217\
        );

    \I__3793\ : SRMux
    port map (
            O => \N__16351\,
            I => \N__16217\
        );

    \I__3792\ : SRMux
    port map (
            O => \N__16350\,
            I => \N__16217\
        );

    \I__3791\ : Glb2LocalMux
    port map (
            O => \N__16347\,
            I => \N__16217\
        );

    \I__3790\ : Glb2LocalMux
    port map (
            O => \N__16344\,
            I => \N__16217\
        );

    \I__3789\ : Glb2LocalMux
    port map (
            O => \N__16341\,
            I => \N__16217\
        );

    \I__3788\ : SRMux
    port map (
            O => \N__16340\,
            I => \N__16217\
        );

    \I__3787\ : GlobalMux
    port map (
            O => \N__16217\,
            I => \N__16214\
        );

    \I__3786\ : gio2CtrlBuf
    port map (
            O => \N__16214\,
            I => \wPllLocked_i_g\
        );

    \I__3785\ : InMux
    port map (
            O => \N__16211\,
            I => \N__16207\
        );

    \I__3784\ : InMux
    port map (
            O => \N__16210\,
            I => \N__16204\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__16207\,
            I => \N__16201\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__16204\,
            I => \uart_inst0.wRxWrData_4\
        );

    \I__3781\ : Odrv4
    port map (
            O => \N__16201\,
            I => \uart_inst0.wRxWrData_4\
        );

    \I__3780\ : InMux
    port map (
            O => \N__16196\,
            I => \N__16193\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__16193\,
            I => \N__16189\
        );

    \I__3778\ : InMux
    port map (
            O => \N__16192\,
            I => \N__16186\
        );

    \I__3777\ : Span4Mux_h
    port map (
            O => \N__16189\,
            I => \N__16183\
        );

    \I__3776\ : LocalMux
    port map (
            O => \N__16186\,
            I => \uart_inst0.wRxWrData_1\
        );

    \I__3775\ : Odrv4
    port map (
            O => \N__16183\,
            I => \uart_inst0.wRxWrData_1\
        );

    \I__3774\ : InMux
    port map (
            O => \N__16178\,
            I => \N__16175\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__16175\,
            I => \N__16172\
        );

    \I__3772\ : Span4Mux_h
    port map (
            O => \N__16172\,
            I => \N__16169\
        );

    \I__3771\ : Odrv4
    port map (
            O => \N__16169\,
            I => \uart_inst0.wRxWrData_0\
        );

    \I__3770\ : InMux
    port map (
            O => \N__16166\,
            I => \N__16163\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__16163\,
            I => \N__16159\
        );

    \I__3768\ : InMux
    port map (
            O => \N__16162\,
            I => \N__16156\
        );

    \I__3767\ : Span4Mux_v
    port map (
            O => \N__16159\,
            I => \N__16153\
        );

    \I__3766\ : LocalMux
    port map (
            O => \N__16156\,
            I => \uart_inst0.wRxWrData_5\
        );

    \I__3765\ : Odrv4
    port map (
            O => \N__16153\,
            I => \uart_inst0.wRxWrData_5\
        );

    \I__3764\ : InMux
    port map (
            O => \N__16148\,
            I => \N__16144\
        );

    \I__3763\ : InMux
    port map (
            O => \N__16147\,
            I => \N__16141\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__16144\,
            I => \N__16138\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__16141\,
            I => \N__16134\
        );

    \I__3760\ : Span4Mux_v
    port map (
            O => \N__16138\,
            I => \N__16131\
        );

    \I__3759\ : InMux
    port map (
            O => \N__16137\,
            I => \N__16128\
        );

    \I__3758\ : Span4Mux_h
    port map (
            O => \N__16134\,
            I => \N__16125\
        );

    \I__3757\ : Odrv4
    port map (
            O => \N__16131\,
            I => \uart_inst0.wRxWrData_7\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__16128\,
            I => \uart_inst0.wRxWrData_7\
        );

    \I__3755\ : Odrv4
    port map (
            O => \N__16125\,
            I => \uart_inst0.wRxWrData_7\
        );

    \I__3754\ : InMux
    port map (
            O => \N__16118\,
            I => \N__16115\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__16115\,
            I => \N__16111\
        );

    \I__3752\ : InMux
    port map (
            O => \N__16114\,
            I => \N__16108\
        );

    \I__3751\ : Span4Mux_h
    port map (
            O => \N__16111\,
            I => \N__16105\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__16108\,
            I => \uart_inst0.wRxWrData_6\
        );

    \I__3749\ : Odrv4
    port map (
            O => \N__16105\,
            I => \uart_inst0.wRxWrData_6\
        );

    \I__3748\ : InMux
    port map (
            O => \N__16100\,
            I => \N__16097\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__16097\,
            I => \N__16093\
        );

    \I__3746\ : InMux
    port map (
            O => \N__16096\,
            I => \N__16090\
        );

    \I__3745\ : Span4Mux_v
    port map (
            O => \N__16093\,
            I => \N__16087\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__16090\,
            I => \uart_inst0.wRxWrData_3\
        );

    \I__3743\ : Odrv4
    port map (
            O => \N__16087\,
            I => \uart_inst0.wRxWrData_3\
        );

    \I__3742\ : InMux
    port map (
            O => \N__16082\,
            I => \N__16078\
        );

    \I__3741\ : InMux
    port map (
            O => \N__16081\,
            I => \N__16075\
        );

    \I__3740\ : LocalMux
    port map (
            O => \N__16078\,
            I => \N__16072\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__16075\,
            I => \uart_inst0.wRxWrData_2\
        );

    \I__3738\ : Odrv4
    port map (
            O => \N__16072\,
            I => \uart_inst0.wRxWrData_2\
        );

    \I__3737\ : CEMux
    port map (
            O => \N__16067\,
            I => \N__16063\
        );

    \I__3736\ : CEMux
    port map (
            O => \N__16066\,
            I => \N__16060\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__16063\,
            I => \N__16057\
        );

    \I__3734\ : LocalMux
    port map (
            O => \N__16060\,
            I => \N__16054\
        );

    \I__3733\ : Odrv4
    port map (
            O => \N__16057\,
            I => \uart_inst0.uart_inst0.rRxData_0_sqmuxa_0\
        );

    \I__3732\ : Odrv4
    port map (
            O => \N__16054\,
            I => \uart_inst0.uart_inst0.rRxData_0_sqmuxa_0\
        );

    \I__3731\ : InMux
    port map (
            O => \N__16049\,
            I => \N__16045\
        );

    \I__3730\ : InMux
    port map (
            O => \N__16048\,
            I => \N__16041\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__16045\,
            I => \N__16038\
        );

    \I__3728\ : CascadeMux
    port map (
            O => \N__16044\,
            I => \N__16029\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__16041\,
            I => \N__16026\
        );

    \I__3726\ : Span4Mux_h
    port map (
            O => \N__16038\,
            I => \N__16023\
        );

    \I__3725\ : InMux
    port map (
            O => \N__16037\,
            I => \N__16019\
        );

    \I__3724\ : InMux
    port map (
            O => \N__16036\,
            I => \N__16014\
        );

    \I__3723\ : InMux
    port map (
            O => \N__16035\,
            I => \N__16014\
        );

    \I__3722\ : InMux
    port map (
            O => \N__16034\,
            I => \N__16009\
        );

    \I__3721\ : InMux
    port map (
            O => \N__16033\,
            I => \N__16009\
        );

    \I__3720\ : InMux
    port map (
            O => \N__16032\,
            I => \N__16004\
        );

    \I__3719\ : InMux
    port map (
            O => \N__16029\,
            I => \N__16004\
        );

    \I__3718\ : Span4Mux_v
    port map (
            O => \N__16026\,
            I => \N__16001\
        );

    \I__3717\ : Span4Mux_v
    port map (
            O => \N__16023\,
            I => \N__15998\
        );

    \I__3716\ : InMux
    port map (
            O => \N__16022\,
            I => \N__15995\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__16019\,
            I => \N__15990\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__16014\,
            I => \N__15990\
        );

    \I__3713\ : LocalMux
    port map (
            O => \N__16009\,
            I => \N__15985\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__16004\,
            I => \N__15985\
        );

    \I__3711\ : Odrv4
    port map (
            O => \N__16001\,
            I => \uart_inst0.uart_inst0.rx_stateZ0Z_2\
        );

    \I__3710\ : Odrv4
    port map (
            O => \N__15998\,
            I => \uart_inst0.uart_inst0.rx_stateZ0Z_2\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__15995\,
            I => \uart_inst0.uart_inst0.rx_stateZ0Z_2\
        );

    \I__3708\ : Odrv4
    port map (
            O => \N__15990\,
            I => \uart_inst0.uart_inst0.rx_stateZ0Z_2\
        );

    \I__3707\ : Odrv4
    port map (
            O => \N__15985\,
            I => \uart_inst0.uart_inst0.rx_stateZ0Z_2\
        );

    \I__3706\ : CascadeMux
    port map (
            O => \N__15974\,
            I => \N__15970\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__15973\,
            I => \N__15966\
        );

    \I__3704\ : InMux
    port map (
            O => \N__15970\,
            I => \N__15961\
        );

    \I__3703\ : InMux
    port map (
            O => \N__15969\,
            I => \N__15958\
        );

    \I__3702\ : InMux
    port map (
            O => \N__15966\,
            I => \N__15953\
        );

    \I__3701\ : InMux
    port map (
            O => \N__15965\,
            I => \N__15953\
        );

    \I__3700\ : InMux
    port map (
            O => \N__15964\,
            I => \N__15950\
        );

    \I__3699\ : LocalMux
    port map (
            O => \N__15961\,
            I => \N__15943\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__15958\,
            I => \N__15943\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__15953\,
            I => \N__15943\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__15950\,
            I => \uart_inst0.uart_inst0.rx_bits_remainingZ0Z_0\
        );

    \I__3695\ : Odrv4
    port map (
            O => \N__15943\,
            I => \uart_inst0.uart_inst0.rx_bits_remainingZ0Z_0\
        );

    \I__3694\ : InMux
    port map (
            O => \N__15938\,
            I => \N__15934\
        );

    \I__3693\ : InMux
    port map (
            O => \N__15937\,
            I => \N__15930\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__15934\,
            I => \N__15927\
        );

    \I__3691\ : InMux
    port map (
            O => \N__15933\,
            I => \N__15924\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__15930\,
            I => \N__15913\
        );

    \I__3689\ : Span4Mux_v
    port map (
            O => \N__15927\,
            I => \N__15913\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__15924\,
            I => \N__15913\
        );

    \I__3687\ : InMux
    port map (
            O => \N__15923\,
            I => \N__15910\
        );

    \I__3686\ : InMux
    port map (
            O => \N__15922\,
            I => \N__15903\
        );

    \I__3685\ : InMux
    port map (
            O => \N__15921\,
            I => \N__15903\
        );

    \I__3684\ : InMux
    port map (
            O => \N__15920\,
            I => \N__15903\
        );

    \I__3683\ : Odrv4
    port map (
            O => \N__15913\,
            I => \uart_inst0.uart_inst0.N_283\
        );

    \I__3682\ : LocalMux
    port map (
            O => \N__15910\,
            I => \uart_inst0.uart_inst0.N_283\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__15903\,
            I => \uart_inst0.uart_inst0.N_283\
        );

    \I__3680\ : InMux
    port map (
            O => \N__15896\,
            I => \N__15892\
        );

    \I__3679\ : InMux
    port map (
            O => \N__15895\,
            I => \N__15888\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__15892\,
            I => \N__15885\
        );

    \I__3677\ : InMux
    port map (
            O => \N__15891\,
            I => \N__15882\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__15888\,
            I => \uart_inst0.uart_inst0.rx_bits_remainingZ0Z_1\
        );

    \I__3675\ : Odrv12
    port map (
            O => \N__15885\,
            I => \uart_inst0.uart_inst0.rx_bits_remainingZ0Z_1\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__15882\,
            I => \uart_inst0.uart_inst0.rx_bits_remainingZ0Z_1\
        );

    \I__3673\ : SRMux
    port map (
            O => \N__15875\,
            I => \N__15871\
        );

    \I__3672\ : SRMux
    port map (
            O => \N__15874\,
            I => \N__15868\
        );

    \I__3671\ : LocalMux
    port map (
            O => \N__15871\,
            I => \N__15865\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__15868\,
            I => \N__15861\
        );

    \I__3669\ : Span4Mux_h
    port map (
            O => \N__15865\,
            I => \N__15858\
        );

    \I__3668\ : InMux
    port map (
            O => \N__15864\,
            I => \N__15855\
        );

    \I__3667\ : Odrv4
    port map (
            O => \N__15861\,
            I => \uart_inst0.uart_inst0.rx_state_2_sqmuxa\
        );

    \I__3666\ : Odrv4
    port map (
            O => \N__15858\,
            I => \uart_inst0.uart_inst0.rx_state_2_sqmuxa\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__15855\,
            I => \uart_inst0.uart_inst0.rx_state_2_sqmuxa\
        );

    \I__3664\ : InMux
    port map (
            O => \N__15848\,
            I => \N__15845\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__15845\,
            I => \N__15842\
        );

    \I__3662\ : Span4Mux_h
    port map (
            O => \N__15842\,
            I => \N__15839\
        );

    \I__3661\ : Odrv4
    port map (
            O => \N__15839\,
            I => \ioFifoData_in_2\
        );

    \I__3660\ : InMux
    port map (
            O => \N__15836\,
            I => \N__15832\
        );

    \I__3659\ : InMux
    port map (
            O => \N__15835\,
            I => \N__15829\
        );

    \I__3658\ : LocalMux
    port map (
            O => \N__15832\,
            I => \fifo_inst.wRxWrData_2\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__15829\,
            I => \fifo_inst.wRxWrData_2\
        );

    \I__3656\ : InMux
    port map (
            O => \N__15824\,
            I => \N__15818\
        );

    \I__3655\ : InMux
    port map (
            O => \N__15823\,
            I => \N__15815\
        );

    \I__3654\ : InMux
    port map (
            O => \N__15822\,
            I => \N__15812\
        );

    \I__3653\ : InMux
    port map (
            O => \N__15821\,
            I => \N__15809\
        );

    \I__3652\ : LocalMux
    port map (
            O => \N__15818\,
            I => \uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7\
        );

    \I__3651\ : LocalMux
    port map (
            O => \N__15815\,
            I => \uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__15812\,
            I => \uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__15809\,
            I => \uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7\
        );

    \I__3648\ : InMux
    port map (
            O => \N__15800\,
            I => \N__15795\
        );

    \I__3647\ : CascadeMux
    port map (
            O => \N__15799\,
            I => \N__15791\
        );

    \I__3646\ : CascadeMux
    port map (
            O => \N__15798\,
            I => \N__15786\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__15795\,
            I => \N__15783\
        );

    \I__3644\ : InMux
    port map (
            O => \N__15794\,
            I => \N__15780\
        );

    \I__3643\ : InMux
    port map (
            O => \N__15791\,
            I => \N__15777\
        );

    \I__3642\ : InMux
    port map (
            O => \N__15790\,
            I => \N__15774\
        );

    \I__3641\ : CEMux
    port map (
            O => \N__15789\,
            I => \N__15771\
        );

    \I__3640\ : InMux
    port map (
            O => \N__15786\,
            I => \N__15768\
        );

    \I__3639\ : Odrv4
    port map (
            O => \N__15783\,
            I => \uart_inst0.rx_uart_fifo_inst.wRamRdEn\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__15780\,
            I => \uart_inst0.rx_uart_fifo_inst.wRamRdEn\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__15777\,
            I => \uart_inst0.rx_uart_fifo_inst.wRamRdEn\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__15774\,
            I => \uart_inst0.rx_uart_fifo_inst.wRamRdEn\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__15771\,
            I => \uart_inst0.rx_uart_fifo_inst.wRamRdEn\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__15768\,
            I => \uart_inst0.rx_uart_fifo_inst.wRamRdEn\
        );

    \I__3633\ : InMux
    port map (
            O => \N__15755\,
            I => \N__15752\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__15752\,
            I => \N__15748\
        );

    \I__3631\ : InMux
    port map (
            O => \N__15751\,
            I => \N__15745\
        );

    \I__3630\ : Odrv4
    port map (
            O => \N__15748\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNIO6JSZ0\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__15745\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNIO6JSZ0\
        );

    \I__3628\ : CascadeMux
    port map (
            O => \N__15740\,
            I => \N__15737\
        );

    \I__3627\ : InMux
    port map (
            O => \N__15737\,
            I => \N__15734\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__15734\,
            I => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_2_0\
        );

    \I__3625\ : InMux
    port map (
            O => \N__15731\,
            I => \N__15727\
        );

    \I__3624\ : InMux
    port map (
            O => \N__15730\,
            I => \N__15724\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__15727\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI0JNSZ0\
        );

    \I__3622\ : LocalMux
    port map (
            O => \N__15724\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI0JNSZ0\
        );

    \I__3621\ : CascadeMux
    port map (
            O => \N__15719\,
            I => \N__15716\
        );

    \I__3620\ : InMux
    port map (
            O => \N__15716\,
            I => \N__15713\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__15713\,
            I => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_6_0\
        );

    \I__3618\ : InMux
    port map (
            O => \N__15710\,
            I => \N__15706\
        );

    \I__3617\ : InMux
    port map (
            O => \N__15709\,
            I => \N__15703\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__15706\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIM3ISZ0\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__15703\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIM3ISZ0\
        );

    \I__3614\ : CascadeMux
    port map (
            O => \N__15698\,
            I => \N__15695\
        );

    \I__3613\ : InMux
    port map (
            O => \N__15695\,
            I => \N__15692\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__15692\,
            I => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_1_0\
        );

    \I__3611\ : InMux
    port map (
            O => \N__15689\,
            I => \N__15685\
        );

    \I__3610\ : InMux
    port map (
            O => \N__15688\,
            I => \N__15682\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__15685\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI2MOSZ0\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__15682\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI2MOSZ0\
        );

    \I__3607\ : CascadeMux
    port map (
            O => \N__15677\,
            I => \N__15674\
        );

    \I__3606\ : InMux
    port map (
            O => \N__15674\,
            I => \N__15671\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__15671\,
            I => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_7_0\
        );

    \I__3604\ : InMux
    port map (
            O => \N__15668\,
            I => \N__15665\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__15665\,
            I => \N__15662\
        );

    \I__3602\ : Odrv4
    port map (
            O => \N__15662\,
            I => \uart_inst0.uart_inst0.un1_rx_bits_remaining_c1\
        );

    \I__3601\ : InMux
    port map (
            O => \N__15659\,
            I => \N__15656\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__15656\,
            I => \N__15651\
        );

    \I__3599\ : InMux
    port map (
            O => \N__15655\,
            I => \N__15646\
        );

    \I__3598\ : InMux
    port map (
            O => \N__15654\,
            I => \N__15646\
        );

    \I__3597\ : Odrv4
    port map (
            O => \N__15651\,
            I => \uart_inst0.uart_inst0.rx_bits_remaining_2_sqmuxa\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__15646\,
            I => \uart_inst0.uart_inst0.rx_bits_remaining_2_sqmuxa\
        );

    \I__3595\ : CascadeMux
    port map (
            O => \N__15641\,
            I => \N__15638\
        );

    \I__3594\ : InMux
    port map (
            O => \N__15638\,
            I => \N__15634\
        );

    \I__3593\ : InMux
    port map (
            O => \N__15637\,
            I => \N__15631\
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__15634\,
            I => \N__15626\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__15631\,
            I => \N__15626\
        );

    \I__3590\ : Odrv4
    port map (
            O => \N__15626\,
            I => \uart_inst0.uart_inst0.rx_bits_remainingZ0Z_2\
        );

    \I__3589\ : InMux
    port map (
            O => \N__15623\,
            I => \N__15619\
        );

    \I__3588\ : InMux
    port map (
            O => \N__15622\,
            I => \N__15616\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__15619\,
            I => \N__15613\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__15616\,
            I => \N__15610\
        );

    \I__3585\ : Odrv4
    port map (
            O => \N__15613\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIQDZ0Z64\
        );

    \I__3584\ : Odrv12
    port map (
            O => \N__15610\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIQDZ0Z64\
        );

    \I__3583\ : CascadeMux
    port map (
            O => \N__15605\,
            I => \N__15602\
        );

    \I__3582\ : InMux
    port map (
            O => \N__15602\,
            I => \N__15599\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__15599\,
            I => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_1\
        );

    \I__3580\ : InMux
    port map (
            O => \N__15596\,
            I => \N__15592\
        );

    \I__3579\ : InMux
    port map (
            O => \N__15595\,
            I => \N__15589\
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__15592\,
            I => \N__15586\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__15589\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNI0NZ0Z94\
        );

    \I__3576\ : Odrv12
    port map (
            O => \N__15586\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNI0NZ0Z94\
        );

    \I__3575\ : CascadeMux
    port map (
            O => \N__15581\,
            I => \N__15578\
        );

    \I__3574\ : InMux
    port map (
            O => \N__15578\,
            I => \N__15575\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__15575\,
            I => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_4\
        );

    \I__3572\ : InMux
    port map (
            O => \N__15572\,
            I => \N__15569\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__15569\,
            I => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_1\
        );

    \I__3570\ : InMux
    port map (
            O => \N__15566\,
            I => \N__15563\
        );

    \I__3569\ : LocalMux
    port map (
            O => \N__15563\,
            I => \N__15560\
        );

    \I__3568\ : Odrv12
    port map (
            O => \N__15560\,
            I => \wUartRxData_1\
        );

    \I__3567\ : InMux
    port map (
            O => \N__15557\,
            I => \N__15554\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__15554\,
            I => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_2\
        );

    \I__3565\ : InMux
    port map (
            O => \N__15551\,
            I => \N__15548\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__15548\,
            I => \N__15545\
        );

    \I__3563\ : Odrv4
    port map (
            O => \N__15545\,
            I => \wUartRxData_2\
        );

    \I__3562\ : InMux
    port map (
            O => \N__15542\,
            I => \N__15539\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__15539\,
            I => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_3\
        );

    \I__3560\ : InMux
    port map (
            O => \N__15536\,
            I => \N__15533\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__15533\,
            I => \N__15530\
        );

    \I__3558\ : Odrv12
    port map (
            O => \N__15530\,
            I => \wUartRxData_3\
        );

    \I__3557\ : InMux
    port map (
            O => \N__15527\,
            I => \N__15524\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__15524\,
            I => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_4\
        );

    \I__3555\ : InMux
    port map (
            O => \N__15521\,
            I => \N__15518\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__15518\,
            I => \N__15515\
        );

    \I__3553\ : Odrv4
    port map (
            O => \N__15515\,
            I => \wUartRxData_4\
        );

    \I__3552\ : InMux
    port map (
            O => \N__15512\,
            I => \N__15508\
        );

    \I__3551\ : InMux
    port map (
            O => \N__15511\,
            I => \N__15505\
        );

    \I__3550\ : LocalMux
    port map (
            O => \N__15508\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIUFMSZ0\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__15505\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIUFMSZ0\
        );

    \I__3548\ : CascadeMux
    port map (
            O => \N__15500\,
            I => \N__15497\
        );

    \I__3547\ : InMux
    port map (
            O => \N__15497\,
            I => \N__15494\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__15494\,
            I => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_5_0\
        );

    \I__3545\ : InMux
    port map (
            O => \N__15491\,
            I => \N__15487\
        );

    \I__3544\ : InMux
    port map (
            O => \N__15490\,
            I => \N__15484\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__15487\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIQ9KSZ0\
        );

    \I__3542\ : LocalMux
    port map (
            O => \N__15484\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIQ9KSZ0\
        );

    \I__3541\ : CascadeMux
    port map (
            O => \N__15479\,
            I => \N__15476\
        );

    \I__3540\ : InMux
    port map (
            O => \N__15476\,
            I => \N__15473\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__15473\,
            I => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_3_0\
        );

    \I__3538\ : InMux
    port map (
            O => \N__15470\,
            I => \N__15467\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__15467\,
            I => \N__15463\
        );

    \I__3536\ : InMux
    port map (
            O => \N__15466\,
            I => \N__15460\
        );

    \I__3535\ : Odrv4
    port map (
            O => \N__15463\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNID4JC2Z0Z_0\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__15460\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNID4JC2Z0Z_0\
        );

    \I__3533\ : CascadeMux
    port map (
            O => \N__15455\,
            I => \N__15452\
        );

    \I__3532\ : InMux
    port map (
            O => \N__15452\,
            I => \N__15449\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__15449\,
            I => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_8\
        );

    \I__3530\ : InMux
    port map (
            O => \N__15446\,
            I => \N__15442\
        );

    \I__3529\ : InMux
    port map (
            O => \N__15445\,
            I => \N__15439\
        );

    \I__3528\ : LocalMux
    port map (
            O => \N__15442\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNISCLSZ0\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__15439\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNISCLSZ0\
        );

    \I__3526\ : CascadeMux
    port map (
            O => \N__15434\,
            I => \N__15431\
        );

    \I__3525\ : InMux
    port map (
            O => \N__15431\,
            I => \N__15428\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__15428\,
            I => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_4_0\
        );

    \I__3523\ : InMux
    port map (
            O => \N__15425\,
            I => \N__15422\
        );

    \I__3522\ : LocalMux
    port map (
            O => \N__15422\,
            I => \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_0\
        );

    \I__3521\ : IoInMux
    port map (
            O => \N__15419\,
            I => \N__15416\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__15416\,
            I => \N__15413\
        );

    \I__3519\ : IoSpan4Mux
    port map (
            O => \N__15413\,
            I => \N__15408\
        );

    \I__3518\ : InMux
    port map (
            O => \N__15412\,
            I => \N__15403\
        );

    \I__3517\ : InMux
    port map (
            O => \N__15411\,
            I => \N__15403\
        );

    \I__3516\ : Span4Mux_s3_v
    port map (
            O => \N__15408\,
            I => \N__15394\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__15403\,
            I => \N__15391\
        );

    \I__3514\ : InMux
    port map (
            O => \N__15402\,
            I => \N__15378\
        );

    \I__3513\ : InMux
    port map (
            O => \N__15401\,
            I => \N__15378\
        );

    \I__3512\ : InMux
    port map (
            O => \N__15400\,
            I => \N__15378\
        );

    \I__3511\ : InMux
    port map (
            O => \N__15399\,
            I => \N__15378\
        );

    \I__3510\ : InMux
    port map (
            O => \N__15398\,
            I => \N__15378\
        );

    \I__3509\ : InMux
    port map (
            O => \N__15397\,
            I => \N__15378\
        );

    \I__3508\ : Span4Mux_h
    port map (
            O => \N__15394\,
            I => \N__15369\
        );

    \I__3507\ : Span4Mux_s3_v
    port map (
            O => \N__15391\,
            I => \N__15369\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__15378\,
            I => \N__15369\
        );

    \I__3505\ : CascadeMux
    port map (
            O => \N__15377\,
            I => \N__15358\
        );

    \I__3504\ : InMux
    port map (
            O => \N__15376\,
            I => \N__15355\
        );

    \I__3503\ : Span4Mux_h
    port map (
            O => \N__15369\,
            I => \N__15352\
        );

    \I__3502\ : InMux
    port map (
            O => \N__15368\,
            I => \N__15349\
        );

    \I__3501\ : InMux
    port map (
            O => \N__15367\,
            I => \N__15338\
        );

    \I__3500\ : InMux
    port map (
            O => \N__15366\,
            I => \N__15338\
        );

    \I__3499\ : InMux
    port map (
            O => \N__15365\,
            I => \N__15338\
        );

    \I__3498\ : InMux
    port map (
            O => \N__15364\,
            I => \N__15338\
        );

    \I__3497\ : InMux
    port map (
            O => \N__15363\,
            I => \N__15338\
        );

    \I__3496\ : InMux
    port map (
            O => \N__15362\,
            I => \N__15331\
        );

    \I__3495\ : InMux
    port map (
            O => \N__15361\,
            I => \N__15331\
        );

    \I__3494\ : InMux
    port map (
            O => \N__15358\,
            I => \N__15331\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__15355\,
            I => \P1A2_c\
        );

    \I__3492\ : Odrv4
    port map (
            O => \N__15352\,
            I => \P1A2_c\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__15349\,
            I => \P1A2_c\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__15338\,
            I => \P1A2_c\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__15331\,
            I => \P1A2_c\
        );

    \I__3488\ : InMux
    port map (
            O => \N__15320\,
            I => \N__15316\
        );

    \I__3487\ : InMux
    port map (
            O => \N__15319\,
            I => \N__15313\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__15316\,
            I => \wRxData_0\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__15313\,
            I => \wRxData_0\
        );

    \I__3484\ : CEMux
    port map (
            O => \N__15308\,
            I => \N__15305\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__15305\,
            I => \N__15301\
        );

    \I__3482\ : CEMux
    port map (
            O => \N__15304\,
            I => \N__15298\
        );

    \I__3481\ : Span4Mux_s2_v
    port map (
            O => \N__15301\,
            I => \N__15293\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__15298\,
            I => \N__15293\
        );

    \I__3479\ : Odrv4
    port map (
            O => \N__15293\,
            I => \N_84_mux_i\
        );

    \I__3478\ : CascadeMux
    port map (
            O => \N__15290\,
            I => \N__15287\
        );

    \I__3477\ : InMux
    port map (
            O => \N__15287\,
            I => \N__15283\
        );

    \I__3476\ : InMux
    port map (
            O => \N__15286\,
            I => \N__15280\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__15283\,
            I => \N__15277\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__15280\,
            I => \N__15271\
        );

    \I__3473\ : Span4Mux_v
    port map (
            O => \N__15277\,
            I => \N__15271\
        );

    \I__3472\ : InMux
    port map (
            O => \N__15276\,
            I => \N__15268\
        );

    \I__3471\ : Odrv4
    port map (
            O => \N__15271\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_8\
        );

    \I__3470\ : LocalMux
    port map (
            O => \N__15268\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_8\
        );

    \I__3469\ : CascadeMux
    port map (
            O => \N__15263\,
            I => \N__15260\
        );

    \I__3468\ : InMux
    port map (
            O => \N__15260\,
            I => \N__15257\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__15257\,
            I => \N__15254\
        );

    \I__3466\ : Span4Mux_h
    port map (
            O => \N__15254\,
            I => \N__15249\
        );

    \I__3465\ : InMux
    port map (
            O => \N__15253\,
            I => \N__15246\
        );

    \I__3464\ : InMux
    port map (
            O => \N__15252\,
            I => \N__15243\
        );

    \I__3463\ : Odrv4
    port map (
            O => \N__15249\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_3\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__15246\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_3\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__15243\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_3\
        );

    \I__3460\ : CascadeMux
    port map (
            O => \N__15236\,
            I => \N__15233\
        );

    \I__3459\ : InMux
    port map (
            O => \N__15233\,
            I => \N__15230\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__15230\,
            I => \N__15226\
        );

    \I__3457\ : InMux
    port map (
            O => \N__15229\,
            I => \N__15222\
        );

    \I__3456\ : Span4Mux_v
    port map (
            O => \N__15226\,
            I => \N__15219\
        );

    \I__3455\ : InMux
    port map (
            O => \N__15225\,
            I => \N__15216\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__15222\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_2\
        );

    \I__3453\ : Odrv4
    port map (
            O => \N__15219\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_2\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__15216\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_2\
        );

    \I__3451\ : CascadeMux
    port map (
            O => \N__15209\,
            I => \N__15206\
        );

    \I__3450\ : InMux
    port map (
            O => \N__15206\,
            I => \N__15203\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__15203\,
            I => \N__15199\
        );

    \I__3448\ : InMux
    port map (
            O => \N__15202\,
            I => \N__15195\
        );

    \I__3447\ : Span4Mux_v
    port map (
            O => \N__15199\,
            I => \N__15192\
        );

    \I__3446\ : InMux
    port map (
            O => \N__15198\,
            I => \N__15189\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__15195\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_1\
        );

    \I__3444\ : Odrv4
    port map (
            O => \N__15192\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_1\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__15189\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_1\
        );

    \I__3442\ : CascadeMux
    port map (
            O => \N__15182\,
            I => \uart_inst0.rx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_0_cascade_\
        );

    \I__3441\ : CascadeMux
    port map (
            O => \N__15179\,
            I => \N__15176\
        );

    \I__3440\ : InMux
    port map (
            O => \N__15176\,
            I => \N__15173\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__15173\,
            I => \N__15169\
        );

    \I__3438\ : InMux
    port map (
            O => \N__15172\,
            I => \N__15165\
        );

    \I__3437\ : Span4Mux_h
    port map (
            O => \N__15169\,
            I => \N__15162\
        );

    \I__3436\ : InMux
    port map (
            O => \N__15168\,
            I => \N__15159\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__15165\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_0\
        );

    \I__3434\ : Odrv4
    port map (
            O => \N__15162\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_0\
        );

    \I__3433\ : LocalMux
    port map (
            O => \N__15159\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_0\
        );

    \I__3432\ : CascadeMux
    port map (
            O => \N__15152\,
            I => \N__15149\
        );

    \I__3431\ : InMux
    port map (
            O => \N__15149\,
            I => \N__15145\
        );

    \I__3430\ : InMux
    port map (
            O => \N__15148\,
            I => \N__15142\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__15145\,
            I => \uart_inst0.rx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_6\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__15142\,
            I => \uart_inst0.rx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_6\
        );

    \I__3427\ : CascadeMux
    port map (
            O => \N__15137\,
            I => \N__15134\
        );

    \I__3426\ : InMux
    port map (
            O => \N__15134\,
            I => \N__15131\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__15131\,
            I => \N__15128\
        );

    \I__3424\ : Span4Mux_v
    port map (
            O => \N__15128\,
            I => \N__15123\
        );

    \I__3423\ : InMux
    port map (
            O => \N__15127\,
            I => \N__15120\
        );

    \I__3422\ : InMux
    port map (
            O => \N__15126\,
            I => \N__15117\
        );

    \I__3421\ : Odrv4
    port map (
            O => \N__15123\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_6\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__15120\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_6\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__15117\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_6\
        );

    \I__3418\ : CascadeMux
    port map (
            O => \N__15110\,
            I => \N__15107\
        );

    \I__3417\ : InMux
    port map (
            O => \N__15107\,
            I => \N__15104\
        );

    \I__3416\ : LocalMux
    port map (
            O => \N__15104\,
            I => \N__15101\
        );

    \I__3415\ : Span4Mux_v
    port map (
            O => \N__15101\,
            I => \N__15096\
        );

    \I__3414\ : InMux
    port map (
            O => \N__15100\,
            I => \N__15093\
        );

    \I__3413\ : InMux
    port map (
            O => \N__15099\,
            I => \N__15090\
        );

    \I__3412\ : Odrv4
    port map (
            O => \N__15096\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_5\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__15093\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_5\
        );

    \I__3410\ : LocalMux
    port map (
            O => \N__15090\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_5\
        );

    \I__3409\ : CascadeMux
    port map (
            O => \N__15083\,
            I => \N__15080\
        );

    \I__3408\ : InMux
    port map (
            O => \N__15080\,
            I => \N__15076\
        );

    \I__3407\ : CascadeMux
    port map (
            O => \N__15079\,
            I => \N__15073\
        );

    \I__3406\ : LocalMux
    port map (
            O => \N__15076\,
            I => \N__15069\
        );

    \I__3405\ : InMux
    port map (
            O => \N__15073\,
            I => \N__15066\
        );

    \I__3404\ : InMux
    port map (
            O => \N__15072\,
            I => \N__15063\
        );

    \I__3403\ : Span4Mux_v
    port map (
            O => \N__15069\,
            I => \N__15060\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__15066\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_7\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__15063\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_7\
        );

    \I__3400\ : Odrv4
    port map (
            O => \N__15060\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_7\
        );

    \I__3399\ : CascadeMux
    port map (
            O => \N__15053\,
            I => \N__15050\
        );

    \I__3398\ : InMux
    port map (
            O => \N__15050\,
            I => \N__15047\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__15047\,
            I => \N__15044\
        );

    \I__3396\ : Span4Mux_v
    port map (
            O => \N__15044\,
            I => \N__15039\
        );

    \I__3395\ : InMux
    port map (
            O => \N__15043\,
            I => \N__15036\
        );

    \I__3394\ : InMux
    port map (
            O => \N__15042\,
            I => \N__15033\
        );

    \I__3393\ : Odrv4
    port map (
            O => \N__15039\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_4\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__15036\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_4\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__15033\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_4\
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__15026\,
            I => \N__15022\
        );

    \I__3389\ : InMux
    port map (
            O => \N__15025\,
            I => \N__15017\
        );

    \I__3388\ : InMux
    port map (
            O => \N__15022\,
            I => \N__15017\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__15017\,
            I => \uart_inst0.rx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_5\
        );

    \I__3386\ : InMux
    port map (
            O => \N__15014\,
            I => \N__15011\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__15011\,
            I => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_5\
        );

    \I__3384\ : InMux
    port map (
            O => \N__15008\,
            I => \N__15004\
        );

    \I__3383\ : InMux
    port map (
            O => \N__15007\,
            I => \N__15001\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__15004\,
            I => \N__14998\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__15001\,
            I => \wUartRxData_5\
        );

    \I__3380\ : Odrv12
    port map (
            O => \N__14998\,
            I => \wUartRxData_5\
        );

    \I__3379\ : CascadeMux
    port map (
            O => \N__14993\,
            I => \N__14990\
        );

    \I__3378\ : InMux
    port map (
            O => \N__14990\,
            I => \N__14987\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__14987\,
            I => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_6\
        );

    \I__3376\ : InMux
    port map (
            O => \N__14984\,
            I => \N__14980\
        );

    \I__3375\ : InMux
    port map (
            O => \N__14983\,
            I => \N__14977\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__14980\,
            I => \N__14974\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__14977\,
            I => \wUartRxData_6\
        );

    \I__3372\ : Odrv12
    port map (
            O => \N__14974\,
            I => \wUartRxData_6\
        );

    \I__3371\ : InMux
    port map (
            O => \N__14969\,
            I => \N__14966\
        );

    \I__3370\ : LocalMux
    port map (
            O => \N__14966\,
            I => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_7\
        );

    \I__3369\ : InMux
    port map (
            O => \N__14963\,
            I => \N__14957\
        );

    \I__3368\ : CascadeMux
    port map (
            O => \N__14962\,
            I => \N__14954\
        );

    \I__3367\ : CascadeMux
    port map (
            O => \N__14961\,
            I => \N__14951\
        );

    \I__3366\ : InMux
    port map (
            O => \N__14960\,
            I => \N__14940\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__14957\,
            I => \N__14937\
        );

    \I__3364\ : InMux
    port map (
            O => \N__14954\,
            I => \N__14934\
        );

    \I__3363\ : InMux
    port map (
            O => \N__14951\,
            I => \N__14931\
        );

    \I__3362\ : InMux
    port map (
            O => \N__14950\,
            I => \N__14928\
        );

    \I__3361\ : InMux
    port map (
            O => \N__14949\,
            I => \N__14925\
        );

    \I__3360\ : InMux
    port map (
            O => \N__14948\,
            I => \N__14918\
        );

    \I__3359\ : InMux
    port map (
            O => \N__14947\,
            I => \N__14918\
        );

    \I__3358\ : InMux
    port map (
            O => \N__14946\,
            I => \N__14918\
        );

    \I__3357\ : InMux
    port map (
            O => \N__14945\,
            I => \N__14911\
        );

    \I__3356\ : InMux
    port map (
            O => \N__14944\,
            I => \N__14911\
        );

    \I__3355\ : InMux
    port map (
            O => \N__14943\,
            I => \N__14911\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__14940\,
            I => \rUartRxEnZ0\
        );

    \I__3353\ : Odrv4
    port map (
            O => \N__14937\,
            I => \rUartRxEnZ0\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__14934\,
            I => \rUartRxEnZ0\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__14931\,
            I => \rUartRxEnZ0\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__14928\,
            I => \rUartRxEnZ0\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__14925\,
            I => \rUartRxEnZ0\
        );

    \I__3348\ : LocalMux
    port map (
            O => \N__14918\,
            I => \rUartRxEnZ0\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__14911\,
            I => \rUartRxEnZ0\
        );

    \I__3346\ : InMux
    port map (
            O => \N__14894\,
            I => \N__14890\
        );

    \I__3345\ : InMux
    port map (
            O => \N__14893\,
            I => \N__14887\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__14890\,
            I => \N__14884\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__14887\,
            I => \wUartRxData_7\
        );

    \I__3342\ : Odrv4
    port map (
            O => \N__14884\,
            I => \wUartRxData_7\
        );

    \I__3341\ : CEMux
    port map (
            O => \N__14879\,
            I => \N__14876\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__14876\,
            I => \N__14873\
        );

    \I__3339\ : Odrv4
    port map (
            O => \N__14873\,
            I => \uart_inst0.rx_uart_fifo_inst.wUartRxEmpty_i\
        );

    \I__3338\ : InMux
    port map (
            O => \N__14870\,
            I => \N__14867\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__14867\,
            I => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_0\
        );

    \I__3336\ : InMux
    port map (
            O => \N__14864\,
            I => \N__14861\
        );

    \I__3335\ : LocalMux
    port map (
            O => \N__14861\,
            I => \N__14858\
        );

    \I__3334\ : Odrv12
    port map (
            O => \N__14858\,
            I => \wUartRxData_0\
        );

    \I__3333\ : InMux
    port map (
            O => \N__14855\,
            I => \N__14852\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__14852\,
            I => \rRamWrAddr_RNI9D19_0\
        );

    \I__3331\ : InMux
    port map (
            O => \N__14849\,
            I => \N__14846\
        );

    \I__3330\ : LocalMux
    port map (
            O => \N__14846\,
            I => \uart_inst0.tx_uart_fifo_inst.N_91\
        );

    \I__3329\ : CascadeMux
    port map (
            O => \N__14843\,
            I => \N__14837\
        );

    \I__3328\ : InMux
    port map (
            O => \N__14842\,
            I => \N__14831\
        );

    \I__3327\ : InMux
    port map (
            O => \N__14841\,
            I => \N__14831\
        );

    \I__3326\ : InMux
    port map (
            O => \N__14840\,
            I => \N__14828\
        );

    \I__3325\ : InMux
    port map (
            O => \N__14837\,
            I => \N__14825\
        );

    \I__3324\ : CEMux
    port map (
            O => \N__14836\,
            I => \N__14822\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__14831\,
            I => \N__14815\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__14828\,
            I => \N__14815\
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__14825\,
            I => \N__14815\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__14822\,
            I => \N__14812\
        );

    \I__3319\ : Span4Mux_s3_v
    port map (
            O => \N__14815\,
            I => \N__14807\
        );

    \I__3318\ : Span4Mux_h
    port map (
            O => \N__14812\,
            I => \N__14807\
        );

    \I__3317\ : Odrv4
    port map (
            O => \N__14807\,
            I => \fifo_inst_rx_fifo_inst_wRamWrEn\
        );

    \I__3316\ : CascadeMux
    port map (
            O => \N__14804\,
            I => \N__14801\
        );

    \I__3315\ : InMux
    port map (
            O => \N__14801\,
            I => \N__14798\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__14798\,
            I => \N__14793\
        );

    \I__3313\ : InMux
    port map (
            O => \N__14797\,
            I => \N__14790\
        );

    \I__3312\ : InMux
    port map (
            O => \N__14796\,
            I => \N__14787\
        );

    \I__3311\ : Odrv4
    port map (
            O => \N__14793\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_0\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__14790\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_0\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__14787\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_0\
        );

    \I__3308\ : InMux
    port map (
            O => \N__14780\,
            I => \N__14777\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__14777\,
            I => \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_4\
        );

    \I__3306\ : InMux
    port map (
            O => \N__14774\,
            I => \N__14771\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__14771\,
            I => \N__14767\
        );

    \I__3304\ : InMux
    port map (
            O => \N__14770\,
            I => \N__14764\
        );

    \I__3303\ : Span4Mux_v
    port map (
            O => \N__14767\,
            I => \N__14761\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__14764\,
            I => \wRxData_4\
        );

    \I__3301\ : Odrv4
    port map (
            O => \N__14761\,
            I => \wRxData_4\
        );

    \I__3300\ : InMux
    port map (
            O => \N__14756\,
            I => \N__14753\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__14753\,
            I => \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_3\
        );

    \I__3298\ : InMux
    port map (
            O => \N__14750\,
            I => \N__14746\
        );

    \I__3297\ : InMux
    port map (
            O => \N__14749\,
            I => \N__14743\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__14746\,
            I => \N__14740\
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__14743\,
            I => \wRxData_3\
        );

    \I__3294\ : Odrv4
    port map (
            O => \N__14740\,
            I => \wRxData_3\
        );

    \I__3293\ : InMux
    port map (
            O => \N__14735\,
            I => \N__14732\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__14732\,
            I => \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_7\
        );

    \I__3291\ : InMux
    port map (
            O => \N__14729\,
            I => \N__14725\
        );

    \I__3290\ : InMux
    port map (
            O => \N__14728\,
            I => \N__14722\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__14725\,
            I => \wRxData_7\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__14722\,
            I => \wRxData_7\
        );

    \I__3287\ : InMux
    port map (
            O => \N__14717\,
            I => \N__14714\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__14714\,
            I => \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_5\
        );

    \I__3285\ : InMux
    port map (
            O => \N__14711\,
            I => \N__14707\
        );

    \I__3284\ : InMux
    port map (
            O => \N__14710\,
            I => \N__14704\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__14707\,
            I => \wRxData_5\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__14704\,
            I => \wRxData_5\
        );

    \I__3281\ : InMux
    port map (
            O => \N__14699\,
            I => \N__14696\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__14696\,
            I => \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_1\
        );

    \I__3279\ : InMux
    port map (
            O => \N__14693\,
            I => \N__14690\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__14690\,
            I => \N__14686\
        );

    \I__3277\ : InMux
    port map (
            O => \N__14689\,
            I => \N__14683\
        );

    \I__3276\ : Odrv4
    port map (
            O => \N__14686\,
            I => \wRxData_1\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__14683\,
            I => \wRxData_1\
        );

    \I__3274\ : InMux
    port map (
            O => \N__14678\,
            I => \N__14675\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__14675\,
            I => \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_2\
        );

    \I__3272\ : InMux
    port map (
            O => \N__14672\,
            I => \N__14668\
        );

    \I__3271\ : InMux
    port map (
            O => \N__14671\,
            I => \N__14665\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__14668\,
            I => \wRxData_2\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__14665\,
            I => \wRxData_2\
        );

    \I__3268\ : InMux
    port map (
            O => \N__14660\,
            I => \N__14657\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__14657\,
            I => \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_6\
        );

    \I__3266\ : InMux
    port map (
            O => \N__14654\,
            I => \N__14650\
        );

    \I__3265\ : InMux
    port map (
            O => \N__14653\,
            I => \N__14647\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__14650\,
            I => \wRxData_6\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__14647\,
            I => \wRxData_6\
        );

    \I__3262\ : SRMux
    port map (
            O => \N__14642\,
            I => \N__14639\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__14639\,
            I => \N__14632\
        );

    \I__3260\ : SRMux
    port map (
            O => \N__14638\,
            I => \N__14629\
        );

    \I__3259\ : SRMux
    port map (
            O => \N__14637\,
            I => \N__14626\
        );

    \I__3258\ : SRMux
    port map (
            O => \N__14636\,
            I => \N__14623\
        );

    \I__3257\ : SRMux
    port map (
            O => \N__14635\,
            I => \N__14620\
        );

    \I__3256\ : Span4Mux_v
    port map (
            O => \N__14632\,
            I => \N__14617\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__14629\,
            I => \N__14614\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__14626\,
            I => \N__14607\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__14623\,
            I => \N__14607\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__14620\,
            I => \N__14607\
        );

    \I__3251\ : Odrv4
    port map (
            O => \N__14617\,
            I => \uart_inst0.uart_inst0.un1_rx_state49_i\
        );

    \I__3250\ : Odrv4
    port map (
            O => \N__14614\,
            I => \uart_inst0.uart_inst0.un1_rx_state49_i\
        );

    \I__3249\ : Odrv4
    port map (
            O => \N__14607\,
            I => \uart_inst0.uart_inst0.un1_rx_state49_i\
        );

    \I__3248\ : InMux
    port map (
            O => \N__14600\,
            I => \N__14594\
        );

    \I__3247\ : InMux
    port map (
            O => \N__14599\,
            I => \N__14594\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__14594\,
            I => \N__14587\
        );

    \I__3245\ : InMux
    port map (
            O => \N__14593\,
            I => \N__14584\
        );

    \I__3244\ : InMux
    port map (
            O => \N__14592\,
            I => \N__14581\
        );

    \I__3243\ : InMux
    port map (
            O => \N__14591\,
            I => \N__14578\
        );

    \I__3242\ : InMux
    port map (
            O => \N__14590\,
            I => \N__14575\
        );

    \I__3241\ : Span4Mux_h
    port map (
            O => \N__14587\,
            I => \N__14572\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__14584\,
            I => \N__14569\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__14581\,
            I => \N__14566\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__14578\,
            I => \uart_inst0.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__14575\,
            I => \uart_inst0.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__3236\ : Odrv4
    port map (
            O => \N__14572\,
            I => \uart_inst0.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__3235\ : Odrv12
    port map (
            O => \N__14569\,
            I => \uart_inst0.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__3234\ : Odrv4
    port map (
            O => \N__14566\,
            I => \uart_inst0.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__3233\ : InMux
    port map (
            O => \N__14555\,
            I => \N__14552\
        );

    \I__3232\ : LocalMux
    port map (
            O => \N__14552\,
            I => \N__14544\
        );

    \I__3231\ : InMux
    port map (
            O => \N__14551\,
            I => \N__14540\
        );

    \I__3230\ : InMux
    port map (
            O => \N__14550\,
            I => \N__14537\
        );

    \I__3229\ : InMux
    port map (
            O => \N__14549\,
            I => \N__14532\
        );

    \I__3228\ : InMux
    port map (
            O => \N__14548\,
            I => \N__14532\
        );

    \I__3227\ : InMux
    port map (
            O => \N__14547\,
            I => \N__14529\
        );

    \I__3226\ : Span4Mux_h
    port map (
            O => \N__14544\,
            I => \N__14526\
        );

    \I__3225\ : InMux
    port map (
            O => \N__14543\,
            I => \N__14523\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__14540\,
            I => \N__14520\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__14537\,
            I => \N__14517\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__14532\,
            I => \uart_inst0.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__14529\,
            I => \uart_inst0.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__3220\ : Odrv4
    port map (
            O => \N__14526\,
            I => \uart_inst0.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__14523\,
            I => \uart_inst0.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__3218\ : Odrv4
    port map (
            O => \N__14520\,
            I => \uart_inst0.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__3217\ : Odrv4
    port map (
            O => \N__14517\,
            I => \uart_inst0.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__3216\ : InMux
    port map (
            O => \N__14504\,
            I => \N__14501\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__14501\,
            I => \N__14497\
        );

    \I__3214\ : InMux
    port map (
            O => \N__14500\,
            I => \N__14494\
        );

    \I__3213\ : Odrv4
    port map (
            O => \N__14497\,
            I => \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_9\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__14494\,
            I => \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_9\
        );

    \I__3211\ : InMux
    port map (
            O => \N__14489\,
            I => \N__14486\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__14486\,
            I => \N__14483\
        );

    \I__3209\ : Odrv4
    port map (
            O => \N__14483\,
            I => \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_11_3\
        );

    \I__3208\ : CascadeMux
    port map (
            O => \N__14480\,
            I => \uart_inst0.uart_inst0.tx_m5_0_2_cascade_\
        );

    \I__3207\ : InMux
    port map (
            O => \N__14477\,
            I => \N__14474\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__14474\,
            I => \N__14471\
        );

    \I__3205\ : Span4Mux_v
    port map (
            O => \N__14471\,
            I => \N__14467\
        );

    \I__3204\ : InMux
    port map (
            O => \N__14470\,
            I => \N__14464\
        );

    \I__3203\ : Odrv4
    port map (
            O => \N__14467\,
            I => \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_11_4\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__14464\,
            I => \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_11_4\
        );

    \I__3201\ : InMux
    port map (
            O => \N__14459\,
            I => \N__14456\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__14456\,
            I => \N__14453\
        );

    \I__3199\ : Odrv4
    port map (
            O => \N__14453\,
            I => \uart_inst0.uart_inst0.tx_N_11_mux\
        );

    \I__3198\ : InMux
    port map (
            O => \N__14450\,
            I => \N__14445\
        );

    \I__3197\ : InMux
    port map (
            O => \N__14449\,
            I => \N__14442\
        );

    \I__3196\ : InMux
    port map (
            O => \N__14448\,
            I => \N__14439\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__14445\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_2\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__14442\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_2\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__14439\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_2\
        );

    \I__3192\ : InMux
    port map (
            O => \N__14432\,
            I => \N__14428\
        );

    \I__3191\ : InMux
    port map (
            O => \N__14431\,
            I => \N__14425\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__14428\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_0\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__14425\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_0\
        );

    \I__3188\ : CascadeMux
    port map (
            O => \N__14420\,
            I => \N__14415\
        );

    \I__3187\ : InMux
    port map (
            O => \N__14419\,
            I => \N__14412\
        );

    \I__3186\ : InMux
    port map (
            O => \N__14418\,
            I => \N__14409\
        );

    \I__3185\ : InMux
    port map (
            O => \N__14415\,
            I => \N__14406\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__14412\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_3\
        );

    \I__3183\ : LocalMux
    port map (
            O => \N__14409\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_3\
        );

    \I__3182\ : LocalMux
    port map (
            O => \N__14406\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_3\
        );

    \I__3181\ : InMux
    port map (
            O => \N__14399\,
            I => \N__14394\
        );

    \I__3180\ : InMux
    port map (
            O => \N__14398\,
            I => \N__14391\
        );

    \I__3179\ : InMux
    port map (
            O => \N__14397\,
            I => \N__14388\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__14394\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_1\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__14391\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_1\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__14388\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_1\
        );

    \I__3175\ : InMux
    port map (
            O => \N__14381\,
            I => \N__14377\
        );

    \I__3174\ : InMux
    port map (
            O => \N__14380\,
            I => \N__14374\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__14377\,
            I => \N__14371\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__14374\,
            I => \uart_inst0.uart_inst0.tx_m5_0\
        );

    \I__3171\ : Odrv4
    port map (
            O => \N__14371\,
            I => \uart_inst0.uart_inst0.tx_m5_0\
        );

    \I__3170\ : InMux
    port map (
            O => \N__14366\,
            I => \N__14363\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__14363\,
            I => \ioFifoData_in_5\
        );

    \I__3168\ : InMux
    port map (
            O => \N__14360\,
            I => \N__14357\
        );

    \I__3167\ : LocalMux
    port map (
            O => \N__14357\,
            I => \N__14353\
        );

    \I__3166\ : InMux
    port map (
            O => \N__14356\,
            I => \N__14350\
        );

    \I__3165\ : Span4Mux_h
    port map (
            O => \N__14353\,
            I => \N__14347\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__14350\,
            I => \fifo_inst.wRxWrData_5\
        );

    \I__3163\ : Odrv4
    port map (
            O => \N__14347\,
            I => \fifo_inst.wRxWrData_5\
        );

    \I__3162\ : CascadeMux
    port map (
            O => \N__14342\,
            I => \N__14339\
        );

    \I__3161\ : InMux
    port map (
            O => \N__14339\,
            I => \N__14336\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__14336\,
            I => \N__14333\
        );

    \I__3159\ : Span4Mux_h
    port map (
            O => \N__14333\,
            I => \N__14328\
        );

    \I__3158\ : InMux
    port map (
            O => \N__14332\,
            I => \N__14325\
        );

    \I__3157\ : InMux
    port map (
            O => \N__14331\,
            I => \N__14322\
        );

    \I__3156\ : Odrv4
    port map (
            O => \N__14328\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_5\
        );

    \I__3155\ : LocalMux
    port map (
            O => \N__14325\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_5\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__14322\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_5\
        );

    \I__3153\ : CascadeMux
    port map (
            O => \N__14315\,
            I => \N__14312\
        );

    \I__3152\ : InMux
    port map (
            O => \N__14312\,
            I => \N__14309\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__14309\,
            I => \N__14304\
        );

    \I__3150\ : InMux
    port map (
            O => \N__14308\,
            I => \N__14301\
        );

    \I__3149\ : InMux
    port map (
            O => \N__14307\,
            I => \N__14298\
        );

    \I__3148\ : Span4Mux_h
    port map (
            O => \N__14304\,
            I => \N__14295\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__14301\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_4\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__14298\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_4\
        );

    \I__3145\ : Odrv4
    port map (
            O => \N__14295\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_4\
        );

    \I__3144\ : CascadeMux
    port map (
            O => \N__14288\,
            I => \N__14284\
        );

    \I__3143\ : CascadeMux
    port map (
            O => \N__14287\,
            I => \N__14281\
        );

    \I__3142\ : InMux
    port map (
            O => \N__14284\,
            I => \N__14278\
        );

    \I__3141\ : InMux
    port map (
            O => \N__14281\,
            I => \N__14275\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__14278\,
            I => \N__14271\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__14275\,
            I => \N__14268\
        );

    \I__3138\ : InMux
    port map (
            O => \N__14274\,
            I => \N__14265\
        );

    \I__3137\ : Span4Mux_v
    port map (
            O => \N__14271\,
            I => \N__14262\
        );

    \I__3136\ : Odrv4
    port map (
            O => \N__14268\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_2\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__14265\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_2\
        );

    \I__3134\ : Odrv4
    port map (
            O => \N__14262\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_2\
        );

    \I__3133\ : CascadeMux
    port map (
            O => \N__14255\,
            I => \N__14252\
        );

    \I__3132\ : InMux
    port map (
            O => \N__14252\,
            I => \N__14249\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__14249\,
            I => \N__14245\
        );

    \I__3130\ : InMux
    port map (
            O => \N__14248\,
            I => \N__14241\
        );

    \I__3129\ : Span4Mux_h
    port map (
            O => \N__14245\,
            I => \N__14238\
        );

    \I__3128\ : InMux
    port map (
            O => \N__14244\,
            I => \N__14235\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__14241\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_7\
        );

    \I__3126\ : Odrv4
    port map (
            O => \N__14238\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_7\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__14235\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_7\
        );

    \I__3124\ : CascadeMux
    port map (
            O => \N__14228\,
            I => \N__14225\
        );

    \I__3123\ : InMux
    port map (
            O => \N__14225\,
            I => \N__14222\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__14222\,
            I => \N__14219\
        );

    \I__3121\ : Span4Mux_h
    port map (
            O => \N__14219\,
            I => \N__14214\
        );

    \I__3120\ : InMux
    port map (
            O => \N__14218\,
            I => \N__14211\
        );

    \I__3119\ : InMux
    port map (
            O => \N__14217\,
            I => \N__14208\
        );

    \I__3118\ : Odrv4
    port map (
            O => \N__14214\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_6\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__14211\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_6\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__14208\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_6\
        );

    \I__3115\ : CascadeMux
    port map (
            O => \N__14201\,
            I => \uart_inst0.tx_uart_fifo_inst.m54_eZ0Z_5_cascade_\
        );

    \I__3114\ : CascadeMux
    port map (
            O => \N__14198\,
            I => \uart_inst0.tx_uart_fifo_inst.N_91_cascade_\
        );

    \I__3113\ : InMux
    port map (
            O => \N__14195\,
            I => \N__14192\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__14192\,
            I => \un1_rRamWrAddr_cry_2_c_RNIOTMG\
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__14189\,
            I => \N__14186\
        );

    \I__3110\ : InMux
    port map (
            O => \N__14186\,
            I => \N__14183\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__14183\,
            I => \N__14178\
        );

    \I__3108\ : InMux
    port map (
            O => \N__14182\,
            I => \N__14175\
        );

    \I__3107\ : InMux
    port map (
            O => \N__14181\,
            I => \N__14172\
        );

    \I__3106\ : Odrv4
    port map (
            O => \N__14178\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_3\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__14175\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_3\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__14172\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_3\
        );

    \I__3103\ : CascadeMux
    port map (
            O => \N__14165\,
            I => \N__14162\
        );

    \I__3102\ : InMux
    port map (
            O => \N__14162\,
            I => \N__14159\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__14159\,
            I => \N__14156\
        );

    \I__3100\ : Span4Mux_h
    port map (
            O => \N__14156\,
            I => \N__14151\
        );

    \I__3099\ : InMux
    port map (
            O => \N__14155\,
            I => \N__14148\
        );

    \I__3098\ : InMux
    port map (
            O => \N__14154\,
            I => \N__14145\
        );

    \I__3097\ : Odrv4
    port map (
            O => \N__14151\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_1\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__14148\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_1\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__14145\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_1\
        );

    \I__3094\ : CascadeMux
    port map (
            O => \N__14138\,
            I => \N__14135\
        );

    \I__3093\ : InMux
    port map (
            O => \N__14135\,
            I => \N__14132\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__14132\,
            I => \N__14127\
        );

    \I__3091\ : CascadeMux
    port map (
            O => \N__14131\,
            I => \N__14124\
        );

    \I__3090\ : InMux
    port map (
            O => \N__14130\,
            I => \N__14121\
        );

    \I__3089\ : Span4Mux_h
    port map (
            O => \N__14127\,
            I => \N__14118\
        );

    \I__3088\ : InMux
    port map (
            O => \N__14124\,
            I => \N__14115\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__14121\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_8\
        );

    \I__3086\ : Odrv4
    port map (
            O => \N__14118\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_8\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__14115\,
            I => \fifo_inst_rx_fifo_inst_rRamWrAddr_8\
        );

    \I__3084\ : InMux
    port map (
            O => \N__14108\,
            I => \N__14105\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__14105\,
            I => \uart_inst0.tx_uart_fifo_inst.m54_eZ0Z_6\
        );

    \I__3082\ : InMux
    port map (
            O => \N__14102\,
            I => \N__14097\
        );

    \I__3081\ : IoInMux
    port map (
            O => \N__14101\,
            I => \N__14094\
        );

    \I__3080\ : InMux
    port map (
            O => \N__14100\,
            I => \N__14091\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__14097\,
            I => \N__14088\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__14094\,
            I => \N__14085\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__14091\,
            I => \N__14082\
        );

    \I__3076\ : Span4Mux_h
    port map (
            O => \N__14088\,
            I => \N__14078\
        );

    \I__3075\ : IoSpan4Mux
    port map (
            O => \N__14085\,
            I => \N__14075\
        );

    \I__3074\ : Span4Mux_v
    port map (
            O => \N__14082\,
            I => \N__14072\
        );

    \I__3073\ : InMux
    port map (
            O => \N__14081\,
            I => \N__14069\
        );

    \I__3072\ : Span4Mux_h
    port map (
            O => \N__14078\,
            I => \N__14063\
        );

    \I__3071\ : Span4Mux_s2_v
    port map (
            O => \N__14075\,
            I => \N__14063\
        );

    \I__3070\ : Span4Mux_v
    port map (
            O => \N__14072\,
            I => \N__14058\
        );

    \I__3069\ : LocalMux
    port map (
            O => \N__14069\,
            I => \N__14058\
        );

    \I__3068\ : InMux
    port map (
            O => \N__14068\,
            I => \N__14055\
        );

    \I__3067\ : Sp12to4
    port map (
            O => \N__14063\,
            I => \N__14052\
        );

    \I__3066\ : Span4Mux_v
    port map (
            O => \N__14058\,
            I => \N__14049\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__14055\,
            I => \N__14046\
        );

    \I__3064\ : Span12Mux_v
    port map (
            O => \N__14052\,
            I => \N__14039\
        );

    \I__3063\ : Sp12to4
    port map (
            O => \N__14049\,
            I => \N__14039\
        );

    \I__3062\ : Sp12to4
    port map (
            O => \N__14046\,
            I => \N__14039\
        );

    \I__3061\ : Odrv12
    port map (
            O => \N__14039\,
            I => \wPllLocked_i\
        );

    \I__3060\ : InMux
    port map (
            O => \N__14036\,
            I => \N__14032\
        );

    \I__3059\ : InMux
    port map (
            O => \N__14035\,
            I => \N__14029\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__14032\,
            I => \uart_inst0.uart_inst0.rRxData_0_sqmuxa\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__14029\,
            I => \uart_inst0.uart_inst0.rRxData_0_sqmuxa\
        );

    \I__3056\ : InMux
    port map (
            O => \N__14024\,
            I => \N__14017\
        );

    \I__3055\ : InMux
    port map (
            O => \N__14023\,
            I => \N__14006\
        );

    \I__3054\ : InMux
    port map (
            O => \N__14022\,
            I => \N__14006\
        );

    \I__3053\ : CascadeMux
    port map (
            O => \N__14021\,
            I => \N__14000\
        );

    \I__3052\ : InMux
    port map (
            O => \N__14020\,
            I => \N__13995\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__14017\,
            I => \N__13992\
        );

    \I__3050\ : InMux
    port map (
            O => \N__14016\,
            I => \N__13987\
        );

    \I__3049\ : InMux
    port map (
            O => \N__14015\,
            I => \N__13987\
        );

    \I__3048\ : InMux
    port map (
            O => \N__14014\,
            I => \N__13983\
        );

    \I__3047\ : CascadeMux
    port map (
            O => \N__14013\,
            I => \N__13980\
        );

    \I__3046\ : CascadeMux
    port map (
            O => \N__14012\,
            I => \N__13977\
        );

    \I__3045\ : CascadeMux
    port map (
            O => \N__14011\,
            I => \N__13974\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__14006\,
            I => \N__13971\
        );

    \I__3043\ : InMux
    port map (
            O => \N__14005\,
            I => \N__13968\
        );

    \I__3042\ : InMux
    port map (
            O => \N__14004\,
            I => \N__13963\
        );

    \I__3041\ : InMux
    port map (
            O => \N__14003\,
            I => \N__13963\
        );

    \I__3040\ : InMux
    port map (
            O => \N__14000\,
            I => \N__13956\
        );

    \I__3039\ : InMux
    port map (
            O => \N__13999\,
            I => \N__13956\
        );

    \I__3038\ : InMux
    port map (
            O => \N__13998\,
            I => \N__13956\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__13995\,
            I => \N__13953\
        );

    \I__3036\ : Span4Mux_v
    port map (
            O => \N__13992\,
            I => \N__13950\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__13987\,
            I => \N__13947\
        );

    \I__3034\ : CascadeMux
    port map (
            O => \N__13986\,
            I => \N__13943\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__13983\,
            I => \N__13940\
        );

    \I__3032\ : InMux
    port map (
            O => \N__13980\,
            I => \N__13937\
        );

    \I__3031\ : InMux
    port map (
            O => \N__13977\,
            I => \N__13932\
        );

    \I__3030\ : InMux
    port map (
            O => \N__13974\,
            I => \N__13932\
        );

    \I__3029\ : Span4Mux_v
    port map (
            O => \N__13971\,
            I => \N__13929\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__13968\,
            I => \N__13922\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__13963\,
            I => \N__13922\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__13956\,
            I => \N__13922\
        );

    \I__3025\ : Span4Mux_s3_v
    port map (
            O => \N__13953\,
            I => \N__13918\
        );

    \I__3024\ : Span4Mux_h
    port map (
            O => \N__13950\,
            I => \N__13913\
        );

    \I__3023\ : Span4Mux_v
    port map (
            O => \N__13947\,
            I => \N__13913\
        );

    \I__3022\ : InMux
    port map (
            O => \N__13946\,
            I => \N__13910\
        );

    \I__3021\ : InMux
    port map (
            O => \N__13943\,
            I => \N__13907\
        );

    \I__3020\ : Span4Mux_v
    port map (
            O => \N__13940\,
            I => \N__13904\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__13937\,
            I => \N__13895\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__13932\,
            I => \N__13895\
        );

    \I__3017\ : Span4Mux_h
    port map (
            O => \N__13929\,
            I => \N__13895\
        );

    \I__3016\ : Span4Mux_v
    port map (
            O => \N__13922\,
            I => \N__13895\
        );

    \I__3015\ : InMux
    port map (
            O => \N__13921\,
            I => \N__13891\
        );

    \I__3014\ : Span4Mux_h
    port map (
            O => \N__13918\,
            I => \N__13888\
        );

    \I__3013\ : Span4Mux_v
    port map (
            O => \N__13913\,
            I => \N__13885\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__13910\,
            I => \N__13880\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__13907\,
            I => \N__13880\
        );

    \I__3010\ : Span4Mux_h
    port map (
            O => \N__13904\,
            I => \N__13875\
        );

    \I__3009\ : Span4Mux_h
    port map (
            O => \N__13895\,
            I => \N__13875\
        );

    \I__3008\ : InMux
    port map (
            O => \N__13894\,
            I => \N__13872\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__13891\,
            I => \N__13869\
        );

    \I__3006\ : Sp12to4
    port map (
            O => \N__13888\,
            I => \N__13866\
        );

    \I__3005\ : Sp12to4
    port map (
            O => \N__13885\,
            I => \N__13857\
        );

    \I__3004\ : Span12Mux_h
    port map (
            O => \N__13880\,
            I => \N__13857\
        );

    \I__3003\ : Sp12to4
    port map (
            O => \N__13875\,
            I => \N__13857\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__13872\,
            I => \N__13857\
        );

    \I__3001\ : Span4Mux_v
    port map (
            O => \N__13869\,
            I => \N__13854\
        );

    \I__3000\ : Span12Mux_v
    port map (
            O => \N__13866\,
            I => \N__13851\
        );

    \I__2999\ : Span12Mux_h
    port map (
            O => \N__13857\,
            I => \N__13848\
        );

    \I__2998\ : Sp12to4
    port map (
            O => \N__13854\,
            I => \N__13845\
        );

    \I__2997\ : Span12Mux_h
    port map (
            O => \N__13851\,
            I => \N__13842\
        );

    \I__2996\ : Span12Mux_v
    port map (
            O => \N__13848\,
            I => \N__13839\
        );

    \I__2995\ : Span12Mux_v
    port map (
            O => \N__13845\,
            I => \N__13836\
        );

    \I__2994\ : Odrv12
    port map (
            O => \N__13842\,
            I => \wPllLocked\
        );

    \I__2993\ : Odrv12
    port map (
            O => \N__13839\,
            I => \wPllLocked\
        );

    \I__2992\ : Odrv12
    port map (
            O => \N__13836\,
            I => \wPllLocked\
        );

    \I__2991\ : InMux
    port map (
            O => \N__13829\,
            I => \N__13826\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__13826\,
            I => \N__13819\
        );

    \I__2989\ : InMux
    port map (
            O => \N__13825\,
            I => \N__13814\
        );

    \I__2988\ : InMux
    port map (
            O => \N__13824\,
            I => \N__13807\
        );

    \I__2987\ : InMux
    port map (
            O => \N__13823\,
            I => \N__13807\
        );

    \I__2986\ : InMux
    port map (
            O => \N__13822\,
            I => \N__13807\
        );

    \I__2985\ : Span4Mux_h
    port map (
            O => \N__13819\,
            I => \N__13804\
        );

    \I__2984\ : InMux
    port map (
            O => \N__13818\,
            I => \N__13799\
        );

    \I__2983\ : InMux
    port map (
            O => \N__13817\,
            I => \N__13799\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__13814\,
            I => \uart_inst0.uart_inst0.N_257_0\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__13807\,
            I => \uart_inst0.uart_inst0.N_257_0\
        );

    \I__2980\ : Odrv4
    port map (
            O => \N__13804\,
            I => \uart_inst0.uart_inst0.N_257_0\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__13799\,
            I => \uart_inst0.uart_inst0.N_257_0\
        );

    \I__2978\ : CascadeMux
    port map (
            O => \N__13790\,
            I => \uart_inst0.uart_inst0.N_273_cascade_\
        );

    \I__2977\ : CascadeMux
    port map (
            O => \N__13787\,
            I => \N__13784\
        );

    \I__2976\ : InMux
    port map (
            O => \N__13784\,
            I => \N__13781\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__13781\,
            I => \N__13775\
        );

    \I__2974\ : InMux
    port map (
            O => \N__13780\,
            I => \N__13772\
        );

    \I__2973\ : InMux
    port map (
            O => \N__13779\,
            I => \N__13768\
        );

    \I__2972\ : InMux
    port map (
            O => \N__13778\,
            I => \N__13765\
        );

    \I__2971\ : Span4Mux_v
    port map (
            O => \N__13775\,
            I => \N__13762\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__13772\,
            I => \N__13759\
        );

    \I__2969\ : InMux
    port map (
            O => \N__13771\,
            I => \N__13756\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__13768\,
            I => \N__13749\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__13765\,
            I => \N__13749\
        );

    \I__2966\ : Span4Mux_h
    port map (
            O => \N__13762\,
            I => \N__13749\
        );

    \I__2965\ : Span4Mux_h
    port map (
            O => \N__13759\,
            I => \N__13746\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__13756\,
            I => \uart_inst0.uart_inst0.rx_stateZ0Z_3\
        );

    \I__2963\ : Odrv4
    port map (
            O => \N__13749\,
            I => \uart_inst0.uart_inst0.rx_stateZ0Z_3\
        );

    \I__2962\ : Odrv4
    port map (
            O => \N__13746\,
            I => \uart_inst0.uart_inst0.rx_stateZ0Z_3\
        );

    \I__2961\ : InMux
    port map (
            O => \N__13739\,
            I => \N__13735\
        );

    \I__2960\ : InMux
    port map (
            O => \N__13738\,
            I => \N__13732\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__13735\,
            I => \N__13729\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__13732\,
            I => \uart_inst0.uart_inst0.rx_state_srsts_0_a5_0_0_3\
        );

    \I__2957\ : Odrv4
    port map (
            O => \N__13729\,
            I => \uart_inst0.uart_inst0.rx_state_srsts_0_a5_0_0_3\
        );

    \I__2956\ : InMux
    port map (
            O => \N__13724\,
            I => \N__13721\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__13721\,
            I => \N__13716\
        );

    \I__2954\ : InMux
    port map (
            O => \N__13720\,
            I => \N__13713\
        );

    \I__2953\ : InMux
    port map (
            O => \N__13719\,
            I => \N__13710\
        );

    \I__2952\ : Span4Mux_v
    port map (
            O => \N__13716\,
            I => \N__13707\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__13713\,
            I => \uart_inst0.uart_inst0.N_274_2\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__13710\,
            I => \uart_inst0.uart_inst0.N_274_2\
        );

    \I__2949\ : Odrv4
    port map (
            O => \N__13707\,
            I => \uart_inst0.uart_inst0.N_274_2\
        );

    \I__2948\ : CascadeMux
    port map (
            O => \N__13700\,
            I => \uart_inst0.uart_inst0.un1_rx_bits_remaining_c3_cascade_\
        );

    \I__2947\ : InMux
    port map (
            O => \N__13697\,
            I => \N__13693\
        );

    \I__2946\ : InMux
    port map (
            O => \N__13696\,
            I => \N__13690\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__13693\,
            I => \uart_inst0.uart_inst0.rx_bits_remainingZ0Z_3\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__13690\,
            I => \uart_inst0.uart_inst0.rx_bits_remainingZ0Z_3\
        );

    \I__2943\ : InMux
    port map (
            O => \N__13685\,
            I => \N__13681\
        );

    \I__2942\ : CascadeMux
    port map (
            O => \N__13684\,
            I => \N__13676\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__13681\,
            I => \N__13673\
        );

    \I__2940\ : CascadeMux
    port map (
            O => \N__13680\,
            I => \N__13670\
        );

    \I__2939\ : CascadeMux
    port map (
            O => \N__13679\,
            I => \N__13667\
        );

    \I__2938\ : InMux
    port map (
            O => \N__13676\,
            I => \N__13664\
        );

    \I__2937\ : Span4Mux_h
    port map (
            O => \N__13673\,
            I => \N__13661\
        );

    \I__2936\ : InMux
    port map (
            O => \N__13670\,
            I => \N__13658\
        );

    \I__2935\ : InMux
    port map (
            O => \N__13667\,
            I => \N__13655\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__13664\,
            I => \N__13652\
        );

    \I__2933\ : Odrv4
    port map (
            O => \N__13661\,
            I => \uart_inst0.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__13658\,
            I => \uart_inst0.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__13655\,
            I => \uart_inst0.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__2930\ : Odrv4
    port map (
            O => \N__13652\,
            I => \uart_inst0.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__2929\ : CascadeMux
    port map (
            O => \N__13643\,
            I => \N__13640\
        );

    \I__2928\ : InMux
    port map (
            O => \N__13640\,
            I => \N__13637\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__13637\,
            I => \uart_inst0.uart_inst0.tx_N_2\
        );

    \I__2926\ : InMux
    port map (
            O => \N__13634\,
            I => \N__13631\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__13631\,
            I => \N__13625\
        );

    \I__2924\ : InMux
    port map (
            O => \N__13630\,
            I => \N__13622\
        );

    \I__2923\ : InMux
    port map (
            O => \N__13629\,
            I => \N__13619\
        );

    \I__2922\ : InMux
    port map (
            O => \N__13628\,
            I => \N__13616\
        );

    \I__2921\ : Span4Mux_v
    port map (
            O => \N__13625\,
            I => \N__13611\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__13622\,
            I => \N__13611\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__13619\,
            I => \uart_inst0.uart_inst0.tx_countdownZ0Z_2\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__13616\,
            I => \uart_inst0.uart_inst0.tx_countdownZ0Z_2\
        );

    \I__2917\ : Odrv4
    port map (
            O => \N__13611\,
            I => \uart_inst0.uart_inst0.tx_countdownZ0Z_2\
        );

    \I__2916\ : SRMux
    port map (
            O => \N__13604\,
            I => \N__13562\
        );

    \I__2915\ : SRMux
    port map (
            O => \N__13603\,
            I => \N__13562\
        );

    \I__2914\ : SRMux
    port map (
            O => \N__13602\,
            I => \N__13562\
        );

    \I__2913\ : SRMux
    port map (
            O => \N__13601\,
            I => \N__13562\
        );

    \I__2912\ : SRMux
    port map (
            O => \N__13600\,
            I => \N__13562\
        );

    \I__2911\ : SRMux
    port map (
            O => \N__13599\,
            I => \N__13562\
        );

    \I__2910\ : SRMux
    port map (
            O => \N__13598\,
            I => \N__13562\
        );

    \I__2909\ : SRMux
    port map (
            O => \N__13597\,
            I => \N__13562\
        );

    \I__2908\ : SRMux
    port map (
            O => \N__13596\,
            I => \N__13562\
        );

    \I__2907\ : SRMux
    port map (
            O => \N__13595\,
            I => \N__13562\
        );

    \I__2906\ : SRMux
    port map (
            O => \N__13594\,
            I => \N__13562\
        );

    \I__2905\ : SRMux
    port map (
            O => \N__13593\,
            I => \N__13562\
        );

    \I__2904\ : SRMux
    port map (
            O => \N__13592\,
            I => \N__13562\
        );

    \I__2903\ : SRMux
    port map (
            O => \N__13591\,
            I => \N__13562\
        );

    \I__2902\ : GlobalMux
    port map (
            O => \N__13562\,
            I => \N__13559\
        );

    \I__2901\ : gio2CtrlBuf
    port map (
            O => \N__13559\,
            I => \N_292_g\
        );

    \I__2900\ : CascadeMux
    port map (
            O => \N__13556\,
            I => \N__13551\
        );

    \I__2899\ : InMux
    port map (
            O => \N__13555\,
            I => \N__13538\
        );

    \I__2898\ : InMux
    port map (
            O => \N__13554\,
            I => \N__13529\
        );

    \I__2897\ : InMux
    port map (
            O => \N__13551\,
            I => \N__13529\
        );

    \I__2896\ : InMux
    port map (
            O => \N__13550\,
            I => \N__13529\
        );

    \I__2895\ : InMux
    port map (
            O => \N__13549\,
            I => \N__13529\
        );

    \I__2894\ : InMux
    port map (
            O => \N__13548\,
            I => \N__13526\
        );

    \I__2893\ : InMux
    port map (
            O => \N__13547\,
            I => \N__13511\
        );

    \I__2892\ : InMux
    port map (
            O => \N__13546\,
            I => \N__13511\
        );

    \I__2891\ : InMux
    port map (
            O => \N__13545\,
            I => \N__13511\
        );

    \I__2890\ : InMux
    port map (
            O => \N__13544\,
            I => \N__13511\
        );

    \I__2889\ : InMux
    port map (
            O => \N__13543\,
            I => \N__13511\
        );

    \I__2888\ : InMux
    port map (
            O => \N__13542\,
            I => \N__13511\
        );

    \I__2887\ : InMux
    port map (
            O => \N__13541\,
            I => \N__13511\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__13538\,
            I => \N__13505\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__13529\,
            I => \N__13505\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__13526\,
            I => \N__13500\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__13511\,
            I => \N__13500\
        );

    \I__2882\ : InMux
    port map (
            O => \N__13510\,
            I => \N__13497\
        );

    \I__2881\ : Odrv4
    port map (
            O => \N__13505\,
            I => \uart_inst0.uart_inst0.N_147_0_i\
        );

    \I__2880\ : Odrv4
    port map (
            O => \N__13500\,
            I => \uart_inst0.uart_inst0.N_147_0_i\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__13497\,
            I => \uart_inst0.uart_inst0.N_147_0_i\
        );

    \I__2878\ : InMux
    port map (
            O => \N__13490\,
            I => \N__13487\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__13487\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_2_s1_THRU_CO\
        );

    \I__2876\ : InMux
    port map (
            O => \N__13484\,
            I => \N__13480\
        );

    \I__2875\ : InMux
    port map (
            O => \N__13483\,
            I => \N__13477\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__13480\,
            I => \N__13472\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__13477\,
            I => \N__13472\
        );

    \I__2872\ : Odrv4
    port map (
            O => \N__13472\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIOAZ0Z54\
        );

    \I__2871\ : CascadeMux
    port map (
            O => \N__13469\,
            I => \N__13466\
        );

    \I__2870\ : InMux
    port map (
            O => \N__13466\,
            I => \N__13463\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__13463\,
            I => \N__13460\
        );

    \I__2868\ : Odrv4
    port map (
            O => \N__13460\,
            I => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_0\
        );

    \I__2867\ : CascadeMux
    port map (
            O => \N__13457\,
            I => \N__13453\
        );

    \I__2866\ : InMux
    port map (
            O => \N__13456\,
            I => \N__13450\
        );

    \I__2865\ : InMux
    port map (
            O => \N__13453\,
            I => \N__13447\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__13450\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_6\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__13447\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_6\
        );

    \I__2862\ : InMux
    port map (
            O => \N__13442\,
            I => \N__13438\
        );

    \I__2861\ : InMux
    port map (
            O => \N__13441\,
            I => \N__13435\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__13438\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_5\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__13435\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_5\
        );

    \I__2858\ : CascadeMux
    port map (
            O => \N__13430\,
            I => \N__13427\
        );

    \I__2857\ : InMux
    port map (
            O => \N__13427\,
            I => \N__13423\
        );

    \I__2856\ : InMux
    port map (
            O => \N__13426\,
            I => \N__13420\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__13423\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_7\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__13420\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_7\
        );

    \I__2853\ : InMux
    port map (
            O => \N__13415\,
            I => \N__13411\
        );

    \I__2852\ : InMux
    port map (
            O => \N__13414\,
            I => \N__13408\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__13411\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_4\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__13408\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_4\
        );

    \I__2849\ : CascadeMux
    port map (
            O => \N__13403\,
            I => \N__13400\
        );

    \I__2848\ : InMux
    port map (
            O => \N__13400\,
            I => \N__13397\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__13397\,
            I => \uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_5\
        );

    \I__2846\ : InMux
    port map (
            O => \N__13394\,
            I => \N__13388\
        );

    \I__2845\ : InMux
    port map (
            O => \N__13393\,
            I => \N__13388\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__13388\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_8\
        );

    \I__2843\ : InMux
    port map (
            O => \N__13385\,
            I => \N__13382\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__13382\,
            I => \uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_4\
        );

    \I__2841\ : CascadeMux
    port map (
            O => \N__13379\,
            I => \N__13376\
        );

    \I__2840\ : InMux
    port map (
            O => \N__13376\,
            I => \N__13373\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__13373\,
            I => \N__13367\
        );

    \I__2838\ : InMux
    port map (
            O => \N__13372\,
            I => \N__13364\
        );

    \I__2837\ : InMux
    port map (
            O => \N__13371\,
            I => \N__13359\
        );

    \I__2836\ : InMux
    port map (
            O => \N__13370\,
            I => \N__13359\
        );

    \I__2835\ : Odrv12
    port map (
            O => \N__13367\,
            I => \wUartRxEmpty\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__13364\,
            I => \wUartRxEmpty\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__13359\,
            I => \wUartRxEmpty\
        );

    \I__2832\ : InMux
    port map (
            O => \N__13352\,
            I => \N__13348\
        );

    \I__2831\ : InMux
    port map (
            O => \N__13351\,
            I => \N__13345\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__13348\,
            I => \N__13342\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__13345\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_0\
        );

    \I__2828\ : Odrv4
    port map (
            O => \N__13342\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_0\
        );

    \I__2827\ : CascadeMux
    port map (
            O => \N__13337\,
            I => \N__13334\
        );

    \I__2826\ : InMux
    port map (
            O => \N__13334\,
            I => \N__13330\
        );

    \I__2825\ : InMux
    port map (
            O => \N__13333\,
            I => \N__13327\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__13330\,
            I => \N__13324\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__13327\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_3\
        );

    \I__2822\ : Odrv4
    port map (
            O => \N__13324\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_3\
        );

    \I__2821\ : CascadeMux
    port map (
            O => \N__13319\,
            I => \N__13312\
        );

    \I__2820\ : InMux
    port map (
            O => \N__13318\,
            I => \N__13309\
        );

    \I__2819\ : InMux
    port map (
            O => \N__13317\,
            I => \N__13304\
        );

    \I__2818\ : InMux
    port map (
            O => \N__13316\,
            I => \N__13304\
        );

    \I__2817\ : InMux
    port map (
            O => \N__13315\,
            I => \N__13299\
        );

    \I__2816\ : InMux
    port map (
            O => \N__13312\,
            I => \N__13299\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__13309\,
            I => \N__13291\
        );

    \I__2814\ : LocalMux
    port map (
            O => \N__13304\,
            I => \N__13291\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__13299\,
            I => \N__13291\
        );

    \I__2812\ : InMux
    port map (
            O => \N__13298\,
            I => \N__13287\
        );

    \I__2811\ : Span4Mux_v
    port map (
            O => \N__13291\,
            I => \N__13284\
        );

    \I__2810\ : InMux
    port map (
            O => \N__13290\,
            I => \N__13281\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__13287\,
            I => \N__13274\
        );

    \I__2808\ : Sp12to4
    port map (
            O => \N__13284\,
            I => \N__13274\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__13281\,
            I => \N__13274\
        );

    \I__2806\ : Span12Mux_h
    port map (
            O => \N__13274\,
            I => \N__13271\
        );

    \I__2805\ : Span12Mux_v
    port map (
            O => \N__13271\,
            I => \N__13268\
        );

    \I__2804\ : Odrv12
    port map (
            O => \N__13268\,
            I => \P1A1_c\
        );

    \I__2803\ : InMux
    port map (
            O => \N__13265\,
            I => \N__13260\
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__13264\,
            I => \N__13255\
        );

    \I__2801\ : CascadeMux
    port map (
            O => \N__13263\,
            I => \N__13251\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__13260\,
            I => \N__13247\
        );

    \I__2799\ : InMux
    port map (
            O => \N__13259\,
            I => \N__13242\
        );

    \I__2798\ : InMux
    port map (
            O => \N__13258\,
            I => \N__13242\
        );

    \I__2797\ : InMux
    port map (
            O => \N__13255\,
            I => \N__13239\
        );

    \I__2796\ : InMux
    port map (
            O => \N__13254\,
            I => \N__13236\
        );

    \I__2795\ : InMux
    port map (
            O => \N__13251\,
            I => \N__13231\
        );

    \I__2794\ : InMux
    port map (
            O => \N__13250\,
            I => \N__13231\
        );

    \I__2793\ : Span4Mux_h
    port map (
            O => \N__13247\,
            I => \N__13226\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__13242\,
            I => \N__13226\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__13239\,
            I => \uart_inst0.uart_inst0.rx_stateZ0Z_1\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__13236\,
            I => \uart_inst0.uart_inst0.rx_stateZ0Z_1\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__13231\,
            I => \uart_inst0.uart_inst0.rx_stateZ0Z_1\
        );

    \I__2788\ : Odrv4
    port map (
            O => \N__13226\,
            I => \uart_inst0.uart_inst0.rx_stateZ0Z_1\
        );

    \I__2787\ : InMux
    port map (
            O => \N__13217\,
            I => \N__13213\
        );

    \I__2786\ : InMux
    port map (
            O => \N__13216\,
            I => \N__13210\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__13213\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIK0HSZ0\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__13210\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIK0HSZ0\
        );

    \I__2783\ : InMux
    port map (
            O => \N__13205\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_0\
        );

    \I__2782\ : InMux
    port map (
            O => \N__13202\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_1\
        );

    \I__2781\ : InMux
    port map (
            O => \N__13199\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_2\
        );

    \I__2780\ : InMux
    port map (
            O => \N__13196\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_3\
        );

    \I__2779\ : InMux
    port map (
            O => \N__13193\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_4\
        );

    \I__2778\ : InMux
    port map (
            O => \N__13190\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_5\
        );

    \I__2777\ : InMux
    port map (
            O => \N__13187\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_6\
        );

    \I__2776\ : InMux
    port map (
            O => \N__13184\,
            I => \bfn_17_11_0_\
        );

    \I__2775\ : InMux
    port map (
            O => \N__13181\,
            I => \N__13177\
        );

    \I__2774\ : InMux
    port map (
            O => \N__13180\,
            I => \N__13174\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__13177\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_1\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__13174\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_1\
        );

    \I__2771\ : InMux
    port map (
            O => \N__13169\,
            I => \N__13165\
        );

    \I__2770\ : InMux
    port map (
            O => \N__13168\,
            I => \N__13162\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__13165\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_2\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__13162\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_2\
        );

    \I__2767\ : CascadeMux
    port map (
            O => \N__13157\,
            I => \N__13151\
        );

    \I__2766\ : CascadeMux
    port map (
            O => \N__13156\,
            I => \N__13148\
        );

    \I__2765\ : CEMux
    port map (
            O => \N__13155\,
            I => \N__13143\
        );

    \I__2764\ : InMux
    port map (
            O => \N__13154\,
            I => \N__13137\
        );

    \I__2763\ : InMux
    port map (
            O => \N__13151\,
            I => \N__13134\
        );

    \I__2762\ : InMux
    port map (
            O => \N__13148\,
            I => \N__13131\
        );

    \I__2761\ : InMux
    port map (
            O => \N__13147\,
            I => \N__13126\
        );

    \I__2760\ : InMux
    port map (
            O => \N__13146\,
            I => \N__13126\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__13143\,
            I => \N__13123\
        );

    \I__2758\ : InMux
    port map (
            O => \N__13142\,
            I => \N__13118\
        );

    \I__2757\ : InMux
    port map (
            O => \N__13141\,
            I => \N__13118\
        );

    \I__2756\ : InMux
    port map (
            O => \N__13140\,
            I => \N__13115\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__13137\,
            I => \N__13110\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__13134\,
            I => \N__13110\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__13131\,
            I => \N__13103\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__13126\,
            I => \N__13103\
        );

    \I__2751\ : Span4Mux_h
    port map (
            O => \N__13123\,
            I => \N__13103\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__13118\,
            I => \uart_inst0.rx_uart_fifo_inst.wRamWrEn\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__13115\,
            I => \uart_inst0.rx_uart_fifo_inst.wRamWrEn\
        );

    \I__2748\ : Odrv4
    port map (
            O => \N__13110\,
            I => \uart_inst0.rx_uart_fifo_inst.wRamWrEn\
        );

    \I__2747\ : Odrv4
    port map (
            O => \N__13103\,
            I => \uart_inst0.rx_uart_fifo_inst.wRamWrEn\
        );

    \I__2746\ : InMux
    port map (
            O => \N__13094\,
            I => \N__13085\
        );

    \I__2745\ : InMux
    port map (
            O => \N__13093\,
            I => \N__13082\
        );

    \I__2744\ : InMux
    port map (
            O => \N__13092\,
            I => \N__13075\
        );

    \I__2743\ : InMux
    port map (
            O => \N__13091\,
            I => \N__13075\
        );

    \I__2742\ : InMux
    port map (
            O => \N__13090\,
            I => \N__13075\
        );

    \I__2741\ : InMux
    port map (
            O => \N__13089\,
            I => \N__13070\
        );

    \I__2740\ : InMux
    port map (
            O => \N__13088\,
            I => \N__13070\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__13085\,
            I => \uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_0\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__13082\,
            I => \uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_0\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__13075\,
            I => \uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_0\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__13070\,
            I => \uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_0\
        );

    \I__2735\ : CascadeMux
    port map (
            O => \N__13061\,
            I => \uart_inst0.rx_uart_fifo_inst.rDataCount_RNI3V391Z0Z_2_cascade_\
        );

    \I__2734\ : InMux
    port map (
            O => \N__13058\,
            I => \N__13055\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__13055\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rDataCount15_2_0_0_0\
        );

    \I__2732\ : CascadeMux
    port map (
            O => \N__13052\,
            I => \uart_inst0.rx_uart_fifo_inst.wRamRdEn_cascade_\
        );

    \I__2731\ : InMux
    port map (
            O => \N__13049\,
            I => \N__13046\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__13046\,
            I => \N__13043\
        );

    \I__2729\ : Span12Mux_s7_v
    port map (
            O => \N__13043\,
            I => \N__13037\
        );

    \I__2728\ : InMux
    port map (
            O => \N__13042\,
            I => \N__13034\
        );

    \I__2727\ : InMux
    port map (
            O => \N__13041\,
            I => \N__13031\
        );

    \I__2726\ : InMux
    port map (
            O => \N__13040\,
            I => \N__13028\
        );

    \I__2725\ : Odrv12
    port map (
            O => \N__13037\,
            I => \rUartRxStateZ0Z_0\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__13034\,
            I => \rUartRxStateZ0Z_0\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__13031\,
            I => \rUartRxStateZ0Z_0\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__13028\,
            I => \rUartRxStateZ0Z_0\
        );

    \I__2721\ : InMux
    port map (
            O => \N__13019\,
            I => \N__13016\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__13016\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rDataCount_c2\
        );

    \I__2719\ : InMux
    port map (
            O => \N__13013\,
            I => \N__13007\
        );

    \I__2718\ : InMux
    port map (
            O => \N__13012\,
            I => \N__13007\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__13007\,
            I => \uart_inst0.rx_uart_fifo_inst.rDataCount_0_sqmuxa\
        );

    \I__2716\ : CascadeMux
    port map (
            O => \N__13004\,
            I => \N__12997\
        );

    \I__2715\ : CascadeMux
    port map (
            O => \N__13003\,
            I => \N__12994\
        );

    \I__2714\ : InMux
    port map (
            O => \N__13002\,
            I => \N__12991\
        );

    \I__2713\ : InMux
    port map (
            O => \N__13001\,
            I => \N__12986\
        );

    \I__2712\ : InMux
    port map (
            O => \N__13000\,
            I => \N__12986\
        );

    \I__2711\ : InMux
    port map (
            O => \N__12997\,
            I => \N__12981\
        );

    \I__2710\ : InMux
    port map (
            O => \N__12994\,
            I => \N__12981\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__12991\,
            I => \uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_2\
        );

    \I__2708\ : LocalMux
    port map (
            O => \N__12986\,
            I => \uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_2\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__12981\,
            I => \uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_2\
        );

    \I__2706\ : InMux
    port map (
            O => \N__12974\,
            I => \N__12971\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__12971\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rDataCount_axbxc3_1_1\
        );

    \I__2704\ : CascadeMux
    port map (
            O => \N__12968\,
            I => \N__12963\
        );

    \I__2703\ : CascadeMux
    port map (
            O => \N__12967\,
            I => \N__12959\
        );

    \I__2702\ : InMux
    port map (
            O => \N__12966\,
            I => \N__12954\
        );

    \I__2701\ : InMux
    port map (
            O => \N__12963\,
            I => \N__12949\
        );

    \I__2700\ : InMux
    port map (
            O => \N__12962\,
            I => \N__12949\
        );

    \I__2699\ : InMux
    port map (
            O => \N__12959\,
            I => \N__12942\
        );

    \I__2698\ : InMux
    port map (
            O => \N__12958\,
            I => \N__12942\
        );

    \I__2697\ : InMux
    port map (
            O => \N__12957\,
            I => \N__12942\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__12954\,
            I => \uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_1\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__12949\,
            I => \uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_1\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__12942\,
            I => \uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_1\
        );

    \I__2693\ : CascadeMux
    port map (
            O => \N__12935\,
            I => \N__12931\
        );

    \I__2692\ : InMux
    port map (
            O => \N__12934\,
            I => \N__12922\
        );

    \I__2691\ : InMux
    port map (
            O => \N__12931\,
            I => \N__12922\
        );

    \I__2690\ : InMux
    port map (
            O => \N__12930\,
            I => \N__12917\
        );

    \I__2689\ : InMux
    port map (
            O => \N__12929\,
            I => \N__12917\
        );

    \I__2688\ : InMux
    port map (
            O => \N__12928\,
            I => \N__12912\
        );

    \I__2687\ : InMux
    port map (
            O => \N__12927\,
            I => \N__12912\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__12922\,
            I => \uart_inst0.wRxWrFull_0\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__12917\,
            I => \uart_inst0.wRxWrFull_0\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__12912\,
            I => \uart_inst0.wRxWrFull_0\
        );

    \I__2683\ : InMux
    port map (
            O => \N__12905\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_5\
        );

    \I__2682\ : InMux
    port map (
            O => \N__12902\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_6\
        );

    \I__2681\ : InMux
    port map (
            O => \N__12899\,
            I => \bfn_17_7_0_\
        );

    \I__2680\ : InMux
    port map (
            O => \N__12896\,
            I => \N__12893\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__12893\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNO_0_0_3\
        );

    \I__2678\ : InMux
    port map (
            O => \N__12890\,
            I => \N__12887\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__12887\,
            I => \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNO_0_0_0\
        );

    \I__2676\ : CascadeMux
    port map (
            O => \N__12884\,
            I => \wUartRxEmpty_cascade_\
        );

    \I__2675\ : InMux
    port map (
            O => \N__12881\,
            I => \N__12878\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__12878\,
            I => \N__12875\
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__12875\,
            I => \rRxDataZ0Z_0\
        );

    \I__2672\ : InMux
    port map (
            O => \N__12872\,
            I => \N__12869\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__12869\,
            I => \N__12866\
        );

    \I__2670\ : Span4Mux_h
    port map (
            O => \N__12866\,
            I => \N__12863\
        );

    \I__2669\ : Odrv4
    port map (
            O => \N__12863\,
            I => \rRxDataZ0Z_5\
        );

    \I__2668\ : InMux
    port map (
            O => \N__12860\,
            I => \N__12857\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__12857\,
            I => \N__12854\
        );

    \I__2666\ : Odrv4
    port map (
            O => \N__12854\,
            I => \rRxDataZ0Z_7\
        );

    \I__2665\ : CEMux
    port map (
            O => \N__12851\,
            I => \N__12847\
        );

    \I__2664\ : CEMux
    port map (
            O => \N__12850\,
            I => \N__12844\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__12847\,
            I => \N__12841\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__12844\,
            I => \N__12838\
        );

    \I__2661\ : Span4Mux_h
    port map (
            O => \N__12841\,
            I => \N__12835\
        );

    \I__2660\ : Span4Mux_h
    port map (
            O => \N__12838\,
            I => \N__12832\
        );

    \I__2659\ : Odrv4
    port map (
            O => \N__12835\,
            I => \N_27_0\
        );

    \I__2658\ : Odrv4
    port map (
            O => \N__12832\,
            I => \N_27_0\
        );

    \I__2657\ : InMux
    port map (
            O => \N__12827\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_0\
        );

    \I__2656\ : InMux
    port map (
            O => \N__12824\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_1\
        );

    \I__2655\ : InMux
    port map (
            O => \N__12821\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_2\
        );

    \I__2654\ : InMux
    port map (
            O => \N__12818\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_3\
        );

    \I__2653\ : InMux
    port map (
            O => \N__12815\,
            I => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_4\
        );

    \I__2652\ : InMux
    port map (
            O => \N__12812\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_5\
        );

    \I__2651\ : InMux
    port map (
            O => \N__12809\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_6\
        );

    \I__2650\ : InMux
    port map (
            O => \N__12806\,
            I => \bfn_17_3_0_\
        );

    \I__2649\ : CascadeMux
    port map (
            O => \N__12803\,
            I => \N__12800\
        );

    \I__2648\ : InMux
    port map (
            O => \N__12800\,
            I => \N__12797\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__12797\,
            I => \N__12793\
        );

    \I__2646\ : InMux
    port map (
            O => \N__12796\,
            I => \N__12790\
        );

    \I__2645\ : Span4Mux_s2_v
    port map (
            O => \N__12793\,
            I => \N__12787\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__12790\,
            I => \N__12784\
        );

    \I__2643\ : Odrv4
    port map (
            O => \N__12787\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIGAUPZ0\
        );

    \I__2642\ : Odrv4
    port map (
            O => \N__12784\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIGAUPZ0\
        );

    \I__2641\ : InMux
    port map (
            O => \N__12779\,
            I => \N__12776\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__12776\,
            I => \N__12772\
        );

    \I__2639\ : InMux
    port map (
            O => \N__12775\,
            I => \N__12769\
        );

    \I__2638\ : Odrv4
    port map (
            O => \N__12772\,
            I => \fifo_inst_tx_fifo_inst_rRamRdAddr_2\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__12769\,
            I => \fifo_inst_tx_fifo_inst_rRamRdAddr_2\
        );

    \I__2636\ : InMux
    port map (
            O => \N__12764\,
            I => \N__12759\
        );

    \I__2635\ : InMux
    port map (
            O => \N__12763\,
            I => \N__12751\
        );

    \I__2634\ : InMux
    port map (
            O => \N__12762\,
            I => \N__12746\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__12759\,
            I => \N__12743\
        );

    \I__2632\ : InMux
    port map (
            O => \N__12758\,
            I => \N__12732\
        );

    \I__2631\ : InMux
    port map (
            O => \N__12757\,
            I => \N__12732\
        );

    \I__2630\ : InMux
    port map (
            O => \N__12756\,
            I => \N__12732\
        );

    \I__2629\ : InMux
    port map (
            O => \N__12755\,
            I => \N__12732\
        );

    \I__2628\ : InMux
    port map (
            O => \N__12754\,
            I => \N__12732\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__12751\,
            I => \N__12729\
        );

    \I__2626\ : InMux
    port map (
            O => \N__12750\,
            I => \N__12726\
        );

    \I__2625\ : InMux
    port map (
            O => \N__12749\,
            I => \N__12722\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__12746\,
            I => \N__12719\
        );

    \I__2623\ : Span4Mux_h
    port map (
            O => \N__12743\,
            I => \N__12712\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__12732\,
            I => \N__12712\
        );

    \I__2621\ : Span4Mux_v
    port map (
            O => \N__12729\,
            I => \N__12712\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__12726\,
            I => \N__12709\
        );

    \I__2619\ : InMux
    port map (
            O => \N__12725\,
            I => \N__12706\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__12722\,
            I => \fifo_inst_wRxWrFull\
        );

    \I__2617\ : Odrv12
    port map (
            O => \N__12719\,
            I => \fifo_inst_wRxWrFull\
        );

    \I__2616\ : Odrv4
    port map (
            O => \N__12712\,
            I => \fifo_inst_wRxWrFull\
        );

    \I__2615\ : Odrv4
    port map (
            O => \N__12709\,
            I => \fifo_inst_wRxWrFull\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__12706\,
            I => \fifo_inst_wRxWrFull\
        );

    \I__2613\ : InMux
    port map (
            O => \N__12695\,
            I => \N__12692\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__12692\,
            I => \N__12683\
        );

    \I__2611\ : InMux
    port map (
            O => \N__12691\,
            I => \N__12680\
        );

    \I__2610\ : InMux
    port map (
            O => \N__12690\,
            I => \N__12675\
        );

    \I__2609\ : InMux
    port map (
            O => \N__12689\,
            I => \N__12675\
        );

    \I__2608\ : InMux
    port map (
            O => \N__12688\,
            I => \N__12668\
        );

    \I__2607\ : InMux
    port map (
            O => \N__12687\,
            I => \N__12668\
        );

    \I__2606\ : InMux
    port map (
            O => \N__12686\,
            I => \N__12668\
        );

    \I__2605\ : Span4Mux_h
    port map (
            O => \N__12683\,
            I => \N__12665\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__12680\,
            I => \fifo_inst_rx_fifo_inst_rDataCount_2\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__12675\,
            I => \fifo_inst_rx_fifo_inst_rDataCount_2\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__12668\,
            I => \fifo_inst_rx_fifo_inst_rDataCount_2\
        );

    \I__2601\ : Odrv4
    port map (
            O => \N__12665\,
            I => \fifo_inst_rx_fifo_inst_rDataCount_2\
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__12656\,
            I => \N__12653\
        );

    \I__2599\ : InMux
    port map (
            O => \N__12653\,
            I => \N__12647\
        );

    \I__2598\ : CascadeMux
    port map (
            O => \N__12652\,
            I => \N__12642\
        );

    \I__2597\ : CascadeMux
    port map (
            O => \N__12651\,
            I => \N__12638\
        );

    \I__2596\ : CascadeMux
    port map (
            O => \N__12650\,
            I => \N__12634\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__12647\,
            I => \N__12631\
        );

    \I__2594\ : InMux
    port map (
            O => \N__12646\,
            I => \N__12628\
        );

    \I__2593\ : InMux
    port map (
            O => \N__12645\,
            I => \N__12625\
        );

    \I__2592\ : InMux
    port map (
            O => \N__12642\,
            I => \N__12618\
        );

    \I__2591\ : InMux
    port map (
            O => \N__12641\,
            I => \N__12618\
        );

    \I__2590\ : InMux
    port map (
            O => \N__12638\,
            I => \N__12618\
        );

    \I__2589\ : InMux
    port map (
            O => \N__12637\,
            I => \N__12613\
        );

    \I__2588\ : InMux
    port map (
            O => \N__12634\,
            I => \N__12613\
        );

    \I__2587\ : Span4Mux_h
    port map (
            O => \N__12631\,
            I => \N__12610\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__12628\,
            I => \fifo_inst_rx_fifo_inst_rDataCount_0\
        );

    \I__2585\ : LocalMux
    port map (
            O => \N__12625\,
            I => \fifo_inst_rx_fifo_inst_rDataCount_0\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__12618\,
            I => \fifo_inst_rx_fifo_inst_rDataCount_0\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__12613\,
            I => \fifo_inst_rx_fifo_inst_rDataCount_0\
        );

    \I__2582\ : Odrv4
    port map (
            O => \N__12610\,
            I => \fifo_inst_rx_fifo_inst_rDataCount_0\
        );

    \I__2581\ : InMux
    port map (
            O => \N__12599\,
            I => \N__12595\
        );

    \I__2580\ : CascadeMux
    port map (
            O => \N__12598\,
            I => \N__12589\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__12595\,
            I => \N__12583\
        );

    \I__2578\ : InMux
    port map (
            O => \N__12594\,
            I => \N__12580\
        );

    \I__2577\ : InMux
    port map (
            O => \N__12593\,
            I => \N__12577\
        );

    \I__2576\ : InMux
    port map (
            O => \N__12592\,
            I => \N__12574\
        );

    \I__2575\ : InMux
    port map (
            O => \N__12589\,
            I => \N__12567\
        );

    \I__2574\ : InMux
    port map (
            O => \N__12588\,
            I => \N__12567\
        );

    \I__2573\ : InMux
    port map (
            O => \N__12587\,
            I => \N__12567\
        );

    \I__2572\ : InMux
    port map (
            O => \N__12586\,
            I => \N__12564\
        );

    \I__2571\ : Span4Mux_v
    port map (
            O => \N__12583\,
            I => \N__12561\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__12580\,
            I => \fifo_inst_rx_fifo_inst_rDataCount_1\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__12577\,
            I => \fifo_inst_rx_fifo_inst_rDataCount_1\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__12574\,
            I => \fifo_inst_rx_fifo_inst_rDataCount_1\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__12567\,
            I => \fifo_inst_rx_fifo_inst_rDataCount_1\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__12564\,
            I => \fifo_inst_rx_fifo_inst_rDataCount_1\
        );

    \I__2565\ : Odrv4
    port map (
            O => \N__12561\,
            I => \fifo_inst_rx_fifo_inst_rDataCount_1\
        );

    \I__2564\ : InMux
    port map (
            O => \N__12548\,
            I => \N__12545\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__12545\,
            I => \N__12542\
        );

    \I__2562\ : Span4Mux_h
    port map (
            O => \N__12542\,
            I => \N__12539\
        );

    \I__2561\ : Odrv4
    port map (
            O => \N__12539\,
            I => \rRxDataZ0Z_6\
        );

    \I__2560\ : InMux
    port map (
            O => \N__12536\,
            I => \N__12533\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__12533\,
            I => \N__12530\
        );

    \I__2558\ : Span4Mux_h
    port map (
            O => \N__12530\,
            I => \N__12527\
        );

    \I__2557\ : Odrv4
    port map (
            O => \N__12527\,
            I => \rRxDataZ0Z_1\
        );

    \I__2556\ : CascadeMux
    port map (
            O => \N__12524\,
            I => \N__12521\
        );

    \I__2555\ : InMux
    port map (
            O => \N__12521\,
            I => \N__12518\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__12518\,
            I => \N__12515\
        );

    \I__2553\ : Odrv4
    port map (
            O => \N__12515\,
            I => \rRxDataZ0Z_2\
        );

    \I__2552\ : InMux
    port map (
            O => \N__12512\,
            I => \N__12509\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__12509\,
            I => \N__12506\
        );

    \I__2550\ : Odrv4
    port map (
            O => \N__12506\,
            I => \rRxDataZ0Z_3\
        );

    \I__2549\ : InMux
    port map (
            O => \N__12503\,
            I => \N__12498\
        );

    \I__2548\ : InMux
    port map (
            O => \N__12502\,
            I => \N__12495\
        );

    \I__2547\ : InMux
    port map (
            O => \N__12501\,
            I => \N__12492\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__12498\,
            I => \N__12487\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__12495\,
            I => \N__12487\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__12492\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_12\
        );

    \I__2543\ : Odrv4
    port map (
            O => \N__12487\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_12\
        );

    \I__2542\ : InMux
    port map (
            O => \N__12482\,
            I => \N__12479\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__12479\,
            I => \N__12476\
        );

    \I__2540\ : Odrv4
    port map (
            O => \N__12476\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_11_s1_THRU_CO\
        );

    \I__2539\ : InMux
    port map (
            O => \N__12473\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_11_s1\
        );

    \I__2538\ : IoInMux
    port map (
            O => \N__12470\,
            I => \N__12467\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__12467\,
            I => \N__12464\
        );

    \I__2536\ : IoSpan4Mux
    port map (
            O => \N__12464\,
            I => \N__12461\
        );

    \I__2535\ : Span4Mux_s2_v
    port map (
            O => \N__12461\,
            I => \N__12446\
        );

    \I__2534\ : CascadeMux
    port map (
            O => \N__12460\,
            I => \N__12443\
        );

    \I__2533\ : CascadeMux
    port map (
            O => \N__12459\,
            I => \N__12440\
        );

    \I__2532\ : CascadeMux
    port map (
            O => \N__12458\,
            I => \N__12436\
        );

    \I__2531\ : CascadeMux
    port map (
            O => \N__12457\,
            I => \N__12433\
        );

    \I__2530\ : CascadeMux
    port map (
            O => \N__12456\,
            I => \N__12430\
        );

    \I__2529\ : CascadeMux
    port map (
            O => \N__12455\,
            I => \N__12427\
        );

    \I__2528\ : CascadeMux
    port map (
            O => \N__12454\,
            I => \N__12424\
        );

    \I__2527\ : CascadeMux
    port map (
            O => \N__12453\,
            I => \N__12421\
        );

    \I__2526\ : CascadeMux
    port map (
            O => \N__12452\,
            I => \N__12418\
        );

    \I__2525\ : CascadeMux
    port map (
            O => \N__12451\,
            I => \N__12415\
        );

    \I__2524\ : CascadeMux
    port map (
            O => \N__12450\,
            I => \N__12412\
        );

    \I__2523\ : CascadeMux
    port map (
            O => \N__12449\,
            I => \N__12409\
        );

    \I__2522\ : Span4Mux_v
    port map (
            O => \N__12446\,
            I => \N__12399\
        );

    \I__2521\ : InMux
    port map (
            O => \N__12443\,
            I => \N__12390\
        );

    \I__2520\ : InMux
    port map (
            O => \N__12440\,
            I => \N__12390\
        );

    \I__2519\ : InMux
    port map (
            O => \N__12439\,
            I => \N__12390\
        );

    \I__2518\ : InMux
    port map (
            O => \N__12436\,
            I => \N__12390\
        );

    \I__2517\ : InMux
    port map (
            O => \N__12433\,
            I => \N__12385\
        );

    \I__2516\ : InMux
    port map (
            O => \N__12430\,
            I => \N__12385\
        );

    \I__2515\ : InMux
    port map (
            O => \N__12427\,
            I => \N__12378\
        );

    \I__2514\ : InMux
    port map (
            O => \N__12424\,
            I => \N__12378\
        );

    \I__2513\ : InMux
    port map (
            O => \N__12421\,
            I => \N__12378\
        );

    \I__2512\ : InMux
    port map (
            O => \N__12418\,
            I => \N__12369\
        );

    \I__2511\ : InMux
    port map (
            O => \N__12415\,
            I => \N__12369\
        );

    \I__2510\ : InMux
    port map (
            O => \N__12412\,
            I => \N__12369\
        );

    \I__2509\ : InMux
    port map (
            O => \N__12409\,
            I => \N__12369\
        );

    \I__2508\ : CascadeMux
    port map (
            O => \N__12408\,
            I => \N__12366\
        );

    \I__2507\ : CascadeMux
    port map (
            O => \N__12407\,
            I => \N__12363\
        );

    \I__2506\ : CascadeMux
    port map (
            O => \N__12406\,
            I => \N__12360\
        );

    \I__2505\ : CascadeMux
    port map (
            O => \N__12405\,
            I => \N__12357\
        );

    \I__2504\ : CascadeMux
    port map (
            O => \N__12404\,
            I => \N__12353\
        );

    \I__2503\ : CascadeMux
    port map (
            O => \N__12403\,
            I => \N__12349\
        );

    \I__2502\ : CascadeMux
    port map (
            O => \N__12402\,
            I => \N__12345\
        );

    \I__2501\ : Span4Mux_v
    port map (
            O => \N__12399\,
            I => \N__12327\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__12390\,
            I => \N__12327\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__12385\,
            I => \N__12327\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__12378\,
            I => \N__12327\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__12369\,
            I => \N__12327\
        );

    \I__2496\ : InMux
    port map (
            O => \N__12366\,
            I => \N__12322\
        );

    \I__2495\ : InMux
    port map (
            O => \N__12363\,
            I => \N__12322\
        );

    \I__2494\ : InMux
    port map (
            O => \N__12360\,
            I => \N__12317\
        );

    \I__2493\ : InMux
    port map (
            O => \N__12357\,
            I => \N__12317\
        );

    \I__2492\ : InMux
    port map (
            O => \N__12356\,
            I => \N__12300\
        );

    \I__2491\ : InMux
    port map (
            O => \N__12353\,
            I => \N__12300\
        );

    \I__2490\ : InMux
    port map (
            O => \N__12352\,
            I => \N__12300\
        );

    \I__2489\ : InMux
    port map (
            O => \N__12349\,
            I => \N__12300\
        );

    \I__2488\ : InMux
    port map (
            O => \N__12348\,
            I => \N__12300\
        );

    \I__2487\ : InMux
    port map (
            O => \N__12345\,
            I => \N__12300\
        );

    \I__2486\ : CascadeMux
    port map (
            O => \N__12344\,
            I => \N__12297\
        );

    \I__2485\ : CascadeMux
    port map (
            O => \N__12343\,
            I => \N__12294\
        );

    \I__2484\ : CascadeMux
    port map (
            O => \N__12342\,
            I => \N__12291\
        );

    \I__2483\ : CascadeMux
    port map (
            O => \N__12341\,
            I => \N__12288\
        );

    \I__2482\ : CascadeMux
    port map (
            O => \N__12340\,
            I => \N__12285\
        );

    \I__2481\ : CascadeMux
    port map (
            O => \N__12339\,
            I => \N__12282\
        );

    \I__2480\ : CascadeMux
    port map (
            O => \N__12338\,
            I => \N__12279\
        );

    \I__2479\ : Span4Mux_v
    port map (
            O => \N__12327\,
            I => \N__12271\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__12322\,
            I => \N__12271\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__12317\,
            I => \N__12271\
        );

    \I__2476\ : SRMux
    port map (
            O => \N__12316\,
            I => \N__12268\
        );

    \I__2475\ : SRMux
    port map (
            O => \N__12315\,
            I => \N__12264\
        );

    \I__2474\ : SRMux
    port map (
            O => \N__12314\,
            I => \N__12261\
        );

    \I__2473\ : SRMux
    port map (
            O => \N__12313\,
            I => \N__12258\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__12300\,
            I => \N__12253\
        );

    \I__2471\ : InMux
    port map (
            O => \N__12297\,
            I => \N__12246\
        );

    \I__2470\ : InMux
    port map (
            O => \N__12294\,
            I => \N__12246\
        );

    \I__2469\ : InMux
    port map (
            O => \N__12291\,
            I => \N__12246\
        );

    \I__2468\ : InMux
    port map (
            O => \N__12288\,
            I => \N__12237\
        );

    \I__2467\ : InMux
    port map (
            O => \N__12285\,
            I => \N__12237\
        );

    \I__2466\ : InMux
    port map (
            O => \N__12282\,
            I => \N__12237\
        );

    \I__2465\ : InMux
    port map (
            O => \N__12279\,
            I => \N__12237\
        );

    \I__2464\ : SRMux
    port map (
            O => \N__12278\,
            I => \N__12234\
        );

    \I__2463\ : Span4Mux_v
    port map (
            O => \N__12271\,
            I => \N__12229\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__12268\,
            I => \N__12229\
        );

    \I__2461\ : SRMux
    port map (
            O => \N__12267\,
            I => \N__12226\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__12264\,
            I => \N__12223\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__12261\,
            I => \N__12218\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__12258\,
            I => \N__12218\
        );

    \I__2457\ : SRMux
    port map (
            O => \N__12257\,
            I => \N__12215\
        );

    \I__2456\ : SRMux
    port map (
            O => \N__12256\,
            I => \N__12212\
        );

    \I__2455\ : Span4Mux_v
    port map (
            O => \N__12253\,
            I => \N__12205\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__12246\,
            I => \N__12205\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__12237\,
            I => \N__12205\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__12234\,
            I => \N__12202\
        );

    \I__2451\ : Span4Mux_h
    port map (
            O => \N__12229\,
            I => \N__12197\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__12226\,
            I => \N__12197\
        );

    \I__2449\ : Span4Mux_s3_v
    port map (
            O => \N__12223\,
            I => \N__12192\
        );

    \I__2448\ : Span4Mux_s3_v
    port map (
            O => \N__12218\,
            I => \N__12192\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__12215\,
            I => \N__12189\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__12212\,
            I => \N__12186\
        );

    \I__2445\ : Span4Mux_h
    port map (
            O => \N__12205\,
            I => \N__12183\
        );

    \I__2444\ : Span4Mux_h
    port map (
            O => \N__12202\,
            I => \N__12180\
        );

    \I__2443\ : Span4Mux_v
    port map (
            O => \N__12197\,
            I => \N__12177\
        );

    \I__2442\ : Span4Mux_v
    port map (
            O => \N__12192\,
            I => \N__12172\
        );

    \I__2441\ : Span4Mux_v
    port map (
            O => \N__12189\,
            I => \N__12172\
        );

    \I__2440\ : Span12Mux_h
    port map (
            O => \N__12186\,
            I => \N__12169\
        );

    \I__2439\ : Span4Mux_v
    port map (
            O => \N__12183\,
            I => \N__12166\
        );

    \I__2438\ : Span4Mux_h
    port map (
            O => \N__12180\,
            I => \N__12163\
        );

    \I__2437\ : Span4Mux_h
    port map (
            O => \N__12177\,
            I => \N__12158\
        );

    \I__2436\ : Span4Mux_h
    port map (
            O => \N__12172\,
            I => \N__12158\
        );

    \I__2435\ : Odrv12
    port map (
            O => \N__12169\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2434\ : Odrv4
    port map (
            O => \N__12166\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2433\ : Odrv4
    port map (
            O => \N__12163\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2432\ : Odrv4
    port map (
            O => \N__12158\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2431\ : CascadeMux
    port map (
            O => \N__12149\,
            I => \N__12145\
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__12148\,
            I => \N__12141\
        );

    \I__2429\ : InMux
    port map (
            O => \N__12145\,
            I => \N__12138\
        );

    \I__2428\ : InMux
    port map (
            O => \N__12144\,
            I => \N__12133\
        );

    \I__2427\ : InMux
    port map (
            O => \N__12141\,
            I => \N__12133\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__12138\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_13\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__12133\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_13\
        );

    \I__2424\ : InMux
    port map (
            O => \N__12128\,
            I => \N__12125\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__12125\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_12_s1_THRU_CO\
        );

    \I__2422\ : InMux
    port map (
            O => \N__12122\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_12_s1\
        );

    \I__2421\ : InMux
    port map (
            O => \N__12119\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_13_s1\
        );

    \I__2420\ : InMux
    port map (
            O => \N__12116\,
            I => \N__12112\
        );

    \I__2419\ : InMux
    port map (
            O => \N__12115\,
            I => \N__12109\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__12112\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_14\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__12109\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_14\
        );

    \I__2416\ : CEMux
    port map (
            O => \N__12104\,
            I => \N__12101\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__12101\,
            I => \N__12098\
        );

    \I__2414\ : Span4Mux_h
    port map (
            O => \N__12098\,
            I => \N__12095\
        );

    \I__2413\ : Odrv4
    port map (
            O => \N__12095\,
            I => \uart_inst0.uart_inst0.N_147_0_i_0\
        );

    \I__2412\ : InMux
    port map (
            O => \N__12092\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_0\
        );

    \I__2411\ : InMux
    port map (
            O => \N__12089\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_1\
        );

    \I__2410\ : InMux
    port map (
            O => \N__12086\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_2\
        );

    \I__2409\ : InMux
    port map (
            O => \N__12083\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_3\
        );

    \I__2408\ : InMux
    port map (
            O => \N__12080\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_4\
        );

    \I__2407\ : CascadeMux
    port map (
            O => \N__12077\,
            I => \N__12072\
        );

    \I__2406\ : InMux
    port map (
            O => \N__12076\,
            I => \N__12069\
        );

    \I__2405\ : InMux
    port map (
            O => \N__12075\,
            I => \N__12066\
        );

    \I__2404\ : InMux
    port map (
            O => \N__12072\,
            I => \N__12063\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__12069\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_5\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__12066\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_5\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__12063\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_5\
        );

    \I__2400\ : InMux
    port map (
            O => \N__12056\,
            I => \N__12053\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__12053\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_4_s1_THRU_CO\
        );

    \I__2398\ : InMux
    port map (
            O => \N__12050\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_4_s1\
        );

    \I__2397\ : InMux
    port map (
            O => \N__12047\,
            I => \N__12042\
        );

    \I__2396\ : InMux
    port map (
            O => \N__12046\,
            I => \N__12039\
        );

    \I__2395\ : InMux
    port map (
            O => \N__12045\,
            I => \N__12036\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__12042\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_6\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__12039\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_6\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__12036\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_6\
        );

    \I__2391\ : InMux
    port map (
            O => \N__12029\,
            I => \N__12026\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__12026\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_5_s1_THRU_CO\
        );

    \I__2389\ : InMux
    port map (
            O => \N__12023\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_5_s1\
        );

    \I__2388\ : InMux
    port map (
            O => \N__12020\,
            I => \N__12015\
        );

    \I__2387\ : InMux
    port map (
            O => \N__12019\,
            I => \N__12012\
        );

    \I__2386\ : InMux
    port map (
            O => \N__12018\,
            I => \N__12009\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__12015\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_7\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__12012\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_7\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__12009\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_7\
        );

    \I__2382\ : InMux
    port map (
            O => \N__12002\,
            I => \N__11999\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__11999\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_6_s1_THRU_CO\
        );

    \I__2380\ : InMux
    port map (
            O => \N__11996\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_6_s1\
        );

    \I__2379\ : InMux
    port map (
            O => \N__11993\,
            I => \N__11989\
        );

    \I__2378\ : InMux
    port map (
            O => \N__11992\,
            I => \N__11985\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__11989\,
            I => \N__11982\
        );

    \I__2376\ : InMux
    port map (
            O => \N__11988\,
            I => \N__11979\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__11985\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_8\
        );

    \I__2374\ : Odrv4
    port map (
            O => \N__11982\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_8\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__11979\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_8\
        );

    \I__2372\ : InMux
    port map (
            O => \N__11972\,
            I => \N__11969\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__11969\,
            I => \N__11966\
        );

    \I__2370\ : Odrv4
    port map (
            O => \N__11966\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_7_s1_THRU_CO\
        );

    \I__2369\ : InMux
    port map (
            O => \N__11963\,
            I => \bfn_16_19_0_\
        );

    \I__2368\ : InMux
    port map (
            O => \N__11960\,
            I => \N__11956\
        );

    \I__2367\ : InMux
    port map (
            O => \N__11959\,
            I => \N__11952\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__11956\,
            I => \N__11949\
        );

    \I__2365\ : InMux
    port map (
            O => \N__11955\,
            I => \N__11946\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__11952\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_9\
        );

    \I__2363\ : Odrv4
    port map (
            O => \N__11949\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_9\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__11946\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_9\
        );

    \I__2361\ : InMux
    port map (
            O => \N__11939\,
            I => \N__11936\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__11936\,
            I => \N__11933\
        );

    \I__2359\ : Odrv4
    port map (
            O => \N__11933\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_8_s1_THRU_CO\
        );

    \I__2358\ : InMux
    port map (
            O => \N__11930\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_8_s1\
        );

    \I__2357\ : InMux
    port map (
            O => \N__11927\,
            I => \N__11922\
        );

    \I__2356\ : InMux
    port map (
            O => \N__11926\,
            I => \N__11917\
        );

    \I__2355\ : InMux
    port map (
            O => \N__11925\,
            I => \N__11917\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__11922\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_10\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__11917\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_10\
        );

    \I__2352\ : InMux
    port map (
            O => \N__11912\,
            I => \N__11909\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__11909\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_9_s1_THRU_CO\
        );

    \I__2350\ : InMux
    port map (
            O => \N__11906\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_9_s1\
        );

    \I__2349\ : InMux
    port map (
            O => \N__11903\,
            I => \N__11898\
        );

    \I__2348\ : InMux
    port map (
            O => \N__11902\,
            I => \N__11893\
        );

    \I__2347\ : InMux
    port map (
            O => \N__11901\,
            I => \N__11893\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__11898\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_11\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__11893\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_11\
        );

    \I__2344\ : InMux
    port map (
            O => \N__11888\,
            I => \N__11885\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__11885\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_10_s1_THRU_CO\
        );

    \I__2342\ : InMux
    port map (
            O => \N__11882\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_10_s1\
        );

    \I__2341\ : CascadeMux
    port map (
            O => \N__11879\,
            I => \N__11876\
        );

    \I__2340\ : InMux
    port map (
            O => \N__11876\,
            I => \N__11868\
        );

    \I__2339\ : InMux
    port map (
            O => \N__11875\,
            I => \N__11868\
        );

    \I__2338\ : InMux
    port map (
            O => \N__11874\,
            I => \N__11865\
        );

    \I__2337\ : InMux
    port map (
            O => \N__11873\,
            I => \N__11862\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__11868\,
            I => \N__11850\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__11865\,
            I => \N__11845\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__11862\,
            I => \N__11845\
        );

    \I__2333\ : InMux
    port map (
            O => \N__11861\,
            I => \N__11840\
        );

    \I__2332\ : InMux
    port map (
            O => \N__11860\,
            I => \N__11840\
        );

    \I__2331\ : InMux
    port map (
            O => \N__11859\,
            I => \N__11831\
        );

    \I__2330\ : InMux
    port map (
            O => \N__11858\,
            I => \N__11831\
        );

    \I__2329\ : InMux
    port map (
            O => \N__11857\,
            I => \N__11831\
        );

    \I__2328\ : InMux
    port map (
            O => \N__11856\,
            I => \N__11831\
        );

    \I__2327\ : InMux
    port map (
            O => \N__11855\,
            I => \N__11824\
        );

    \I__2326\ : InMux
    port map (
            O => \N__11854\,
            I => \N__11824\
        );

    \I__2325\ : InMux
    port map (
            O => \N__11853\,
            I => \N__11824\
        );

    \I__2324\ : Odrv4
    port map (
            O => \N__11850\,
            I => \uart_inst0.uart_inst0.N_147_0\
        );

    \I__2323\ : Odrv4
    port map (
            O => \N__11845\,
            I => \uart_inst0.uart_inst0.N_147_0\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__11840\,
            I => \uart_inst0.uart_inst0.N_147_0\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__11831\,
            I => \uart_inst0.uart_inst0.N_147_0\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__11824\,
            I => \uart_inst0.uart_inst0.N_147_0\
        );

    \I__2319\ : CascadeMux
    port map (
            O => \N__11813\,
            I => \N__11810\
        );

    \I__2318\ : InMux
    port map (
            O => \N__11810\,
            I => \N__11807\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__11807\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_0_s1_THRU_CO\
        );

    \I__2316\ : InMux
    port map (
            O => \N__11804\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_0_s1\
        );

    \I__2315\ : InMux
    port map (
            O => \N__11801\,
            I => \N__11798\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__11798\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_1_s1_THRU_CO\
        );

    \I__2313\ : InMux
    port map (
            O => \N__11795\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_1_s1\
        );

    \I__2312\ : InMux
    port map (
            O => \N__11792\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_2_s1\
        );

    \I__2311\ : InMux
    port map (
            O => \N__11789\,
            I => \N__11784\
        );

    \I__2310\ : InMux
    port map (
            O => \N__11788\,
            I => \N__11781\
        );

    \I__2309\ : InMux
    port map (
            O => \N__11787\,
            I => \N__11778\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__11784\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_4\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__11781\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_4\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__11778\,
            I => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_4\
        );

    \I__2305\ : InMux
    port map (
            O => \N__11771\,
            I => \N__11768\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__11768\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_3_s1_THRU_CO\
        );

    \I__2303\ : InMux
    port map (
            O => \N__11765\,
            I => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_3_s1\
        );

    \I__2302\ : InMux
    port map (
            O => \N__11762\,
            I => \N__11759\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__11759\,
            I => \uart_inst0.uart_inst0.rx_countdown_cry_3_THRU_CO\
        );

    \I__2300\ : InMux
    port map (
            O => \N__11756\,
            I => \uart_inst0.uart_inst0.rx_countdown_cry_3\
        );

    \I__2299\ : InMux
    port map (
            O => \N__11753\,
            I => \N__11745\
        );

    \I__2298\ : InMux
    port map (
            O => \N__11752\,
            I => \N__11734\
        );

    \I__2297\ : InMux
    port map (
            O => \N__11751\,
            I => \N__11734\
        );

    \I__2296\ : InMux
    port map (
            O => \N__11750\,
            I => \N__11734\
        );

    \I__2295\ : InMux
    port map (
            O => \N__11749\,
            I => \N__11734\
        );

    \I__2294\ : InMux
    port map (
            O => \N__11748\,
            I => \N__11734\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__11745\,
            I => \uart_inst0.uart_inst0.N_252_0_i\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__11734\,
            I => \uart_inst0.uart_inst0.N_252_0_i\
        );

    \I__2291\ : InMux
    port map (
            O => \N__11729\,
            I => \uart_inst0.uart_inst0.rx_countdown_cry_4\
        );

    \I__2290\ : CascadeMux
    port map (
            O => \N__11726\,
            I => \N__11722\
        );

    \I__2289\ : InMux
    port map (
            O => \N__11725\,
            I => \N__11719\
        );

    \I__2288\ : InMux
    port map (
            O => \N__11722\,
            I => \N__11716\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__11719\,
            I => \uart_inst0.uart_inst0.rx_countdownZ0Z_5\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__11716\,
            I => \uart_inst0.uart_inst0.rx_countdownZ0Z_5\
        );

    \I__2285\ : CEMux
    port map (
            O => \N__11711\,
            I => \N__11707\
        );

    \I__2284\ : CEMux
    port map (
            O => \N__11710\,
            I => \N__11704\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__11707\,
            I => \N__11701\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__11704\,
            I => \N__11698\
        );

    \I__2281\ : Odrv4
    port map (
            O => \N__11701\,
            I => \uart_inst0.uart_inst0.rx_countdowne_0_i\
        );

    \I__2280\ : Odrv4
    port map (
            O => \N__11698\,
            I => \uart_inst0.uart_inst0.rx_countdowne_0_i\
        );

    \I__2279\ : InMux
    port map (
            O => \N__11693\,
            I => \N__11688\
        );

    \I__2278\ : InMux
    port map (
            O => \N__11692\,
            I => \N__11685\
        );

    \I__2277\ : InMux
    port map (
            O => \N__11691\,
            I => \N__11682\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__11688\,
            I => \N__11675\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__11685\,
            I => \N__11675\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__11682\,
            I => \N__11675\
        );

    \I__2273\ : Odrv4
    port map (
            O => \N__11675\,
            I => \uart_inst0.uart_inst0.N_258_0\
        );

    \I__2272\ : CascadeMux
    port map (
            O => \N__11672\,
            I => \uart_inst0.uart_inst0.N_276_cascade_\
        );

    \I__2271\ : InMux
    port map (
            O => \N__11669\,
            I => \N__11666\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__11666\,
            I => \N__11662\
        );

    \I__2269\ : InMux
    port map (
            O => \N__11665\,
            I => \N__11655\
        );

    \I__2268\ : Span4Mux_h
    port map (
            O => \N__11662\,
            I => \N__11645\
        );

    \I__2267\ : InMux
    port map (
            O => \N__11661\,
            I => \N__11640\
        );

    \I__2266\ : InMux
    port map (
            O => \N__11660\,
            I => \N__11640\
        );

    \I__2265\ : InMux
    port map (
            O => \N__11659\,
            I => \N__11637\
        );

    \I__2264\ : InMux
    port map (
            O => \N__11658\,
            I => \N__11634\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__11655\,
            I => \N__11631\
        );

    \I__2262\ : InMux
    port map (
            O => \N__11654\,
            I => \N__11628\
        );

    \I__2261\ : InMux
    port map (
            O => \N__11653\,
            I => \N__11625\
        );

    \I__2260\ : InMux
    port map (
            O => \N__11652\,
            I => \N__11620\
        );

    \I__2259\ : InMux
    port map (
            O => \N__11651\,
            I => \N__11620\
        );

    \I__2258\ : InMux
    port map (
            O => \N__11650\,
            I => \N__11613\
        );

    \I__2257\ : InMux
    port map (
            O => \N__11649\,
            I => \N__11613\
        );

    \I__2256\ : InMux
    port map (
            O => \N__11648\,
            I => \N__11613\
        );

    \I__2255\ : Span4Mux_v
    port map (
            O => \N__11645\,
            I => \N__11606\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__11640\,
            I => \N__11606\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__11637\,
            I => \N__11606\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__11634\,
            I => \uart_inst0.uart_inst0.tx_stateZ0Z_0\
        );

    \I__2251\ : Odrv4
    port map (
            O => \N__11631\,
            I => \uart_inst0.uart_inst0.tx_stateZ0Z_0\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__11628\,
            I => \uart_inst0.uart_inst0.tx_stateZ0Z_0\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__11625\,
            I => \uart_inst0.uart_inst0.tx_stateZ0Z_0\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__11620\,
            I => \uart_inst0.uart_inst0.tx_stateZ0Z_0\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__11613\,
            I => \uart_inst0.uart_inst0.tx_stateZ0Z_0\
        );

    \I__2246\ : Odrv4
    port map (
            O => \N__11606\,
            I => \uart_inst0.uart_inst0.tx_stateZ0Z_0\
        );

    \I__2245\ : InMux
    port map (
            O => \N__11591\,
            I => \N__11588\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__11588\,
            I => \N__11584\
        );

    \I__2243\ : InMux
    port map (
            O => \N__11587\,
            I => \N__11576\
        );

    \I__2242\ : Span4Mux_h
    port map (
            O => \N__11584\,
            I => \N__11572\
        );

    \I__2241\ : CascadeMux
    port map (
            O => \N__11583\,
            I => \N__11569\
        );

    \I__2240\ : CascadeMux
    port map (
            O => \N__11582\,
            I => \N__11566\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__11581\,
            I => \N__11562\
        );

    \I__2238\ : CascadeMux
    port map (
            O => \N__11580\,
            I => \N__11557\
        );

    \I__2237\ : CascadeMux
    port map (
            O => \N__11579\,
            I => \N__11553\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__11576\,
            I => \N__11549\
        );

    \I__2235\ : InMux
    port map (
            O => \N__11575\,
            I => \N__11546\
        );

    \I__2234\ : Span4Mux_v
    port map (
            O => \N__11572\,
            I => \N__11543\
        );

    \I__2233\ : InMux
    port map (
            O => \N__11569\,
            I => \N__11540\
        );

    \I__2232\ : InMux
    port map (
            O => \N__11566\,
            I => \N__11535\
        );

    \I__2231\ : InMux
    port map (
            O => \N__11565\,
            I => \N__11535\
        );

    \I__2230\ : InMux
    port map (
            O => \N__11562\,
            I => \N__11528\
        );

    \I__2229\ : InMux
    port map (
            O => \N__11561\,
            I => \N__11528\
        );

    \I__2228\ : InMux
    port map (
            O => \N__11560\,
            I => \N__11528\
        );

    \I__2227\ : InMux
    port map (
            O => \N__11557\,
            I => \N__11521\
        );

    \I__2226\ : InMux
    port map (
            O => \N__11556\,
            I => \N__11521\
        );

    \I__2225\ : InMux
    port map (
            O => \N__11553\,
            I => \N__11521\
        );

    \I__2224\ : InMux
    port map (
            O => \N__11552\,
            I => \N__11518\
        );

    \I__2223\ : Odrv12
    port map (
            O => \N__11549\,
            I => \uart_inst0.uart_inst0.tx_stateZ0Z_1\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__11546\,
            I => \uart_inst0.uart_inst0.tx_stateZ0Z_1\
        );

    \I__2221\ : Odrv4
    port map (
            O => \N__11543\,
            I => \uart_inst0.uart_inst0.tx_stateZ0Z_1\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__11540\,
            I => \uart_inst0.uart_inst0.tx_stateZ0Z_1\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__11535\,
            I => \uart_inst0.uart_inst0.tx_stateZ0Z_1\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__11528\,
            I => \uart_inst0.uart_inst0.tx_stateZ0Z_1\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__11521\,
            I => \uart_inst0.uart_inst0.tx_stateZ0Z_1\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__11518\,
            I => \uart_inst0.uart_inst0.tx_stateZ0Z_1\
        );

    \I__2215\ : InMux
    port map (
            O => \N__11501\,
            I => \N__11498\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__11498\,
            I => \N__11495\
        );

    \I__2213\ : Odrv4
    port map (
            O => \N__11495\,
            I => \uart_inst0.uart_inst0.un1_m3_0_a2_0\
        );

    \I__2212\ : InMux
    port map (
            O => \N__11492\,
            I => \N__11489\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__11489\,
            I => \uart_inst0.uart_inst0.N_275\
        );

    \I__2210\ : CascadeMux
    port map (
            O => \N__11486\,
            I => \uart_inst0.uart_inst0.N_283_cascade_\
        );

    \I__2209\ : InMux
    port map (
            O => \N__11483\,
            I => \N__11479\
        );

    \I__2208\ : InMux
    port map (
            O => \N__11482\,
            I => \N__11476\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__11479\,
            I => \N__11473\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__11476\,
            I => \N__11470\
        );

    \I__2205\ : Odrv12
    port map (
            O => \N__11473\,
            I => \uart_inst0.uart_inst0.rx_stateZ0Z_6\
        );

    \I__2204\ : Odrv4
    port map (
            O => \N__11470\,
            I => \uart_inst0.uart_inst0.rx_stateZ0Z_6\
        );

    \I__2203\ : InMux
    port map (
            O => \N__11465\,
            I => \N__11459\
        );

    \I__2202\ : InMux
    port map (
            O => \N__11464\,
            I => \N__11459\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__11459\,
            I => \uart_inst0.uart_inst0.rx_state_srsts_0_o2_3_3\
        );

    \I__2200\ : InMux
    port map (
            O => \N__11456\,
            I => \N__11452\
        );

    \I__2199\ : InMux
    port map (
            O => \N__11455\,
            I => \N__11449\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__11452\,
            I => \uart_inst0.uart_inst0.rx_countdown_2_sqmuxa_i_1\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__11449\,
            I => \uart_inst0.uart_inst0.rx_countdown_2_sqmuxa_i_1\
        );

    \I__2196\ : InMux
    port map (
            O => \N__11444\,
            I => \N__11441\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__11441\,
            I => \N__11438\
        );

    \I__2194\ : Odrv12
    port map (
            O => \N__11438\,
            I => \uart_inst0.uart_inst0.un1_rx_clk_divider_0\
        );

    \I__2193\ : CascadeMux
    port map (
            O => \N__11435\,
            I => \uart_inst0.uart_inst0.N_258_0_cascade_\
        );

    \I__2192\ : InMux
    port map (
            O => \N__11432\,
            I => \N__11425\
        );

    \I__2191\ : InMux
    port map (
            O => \N__11431\,
            I => \N__11422\
        );

    \I__2190\ : InMux
    port map (
            O => \N__11430\,
            I => \N__11419\
        );

    \I__2189\ : InMux
    port map (
            O => \N__11429\,
            I => \N__11414\
        );

    \I__2188\ : InMux
    port map (
            O => \N__11428\,
            I => \N__11414\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__11425\,
            I => \uart_inst0.uart_inst0.rx_countdownZ0Z_0\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__11422\,
            I => \uart_inst0.uart_inst0.rx_countdownZ0Z_0\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__11419\,
            I => \uart_inst0.uart_inst0.rx_countdownZ0Z_0\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__11414\,
            I => \uart_inst0.uart_inst0.rx_countdownZ0Z_0\
        );

    \I__2183\ : InMux
    port map (
            O => \N__11405\,
            I => \N__11399\
        );

    \I__2182\ : InMux
    port map (
            O => \N__11404\,
            I => \N__11396\
        );

    \I__2181\ : InMux
    port map (
            O => \N__11403\,
            I => \N__11391\
        );

    \I__2180\ : InMux
    port map (
            O => \N__11402\,
            I => \N__11391\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__11399\,
            I => \uart_inst0.uart_inst0.rx_countdownZ0Z_1\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__11396\,
            I => \uart_inst0.uart_inst0.rx_countdownZ0Z_1\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__11391\,
            I => \uart_inst0.uart_inst0.rx_countdownZ0Z_1\
        );

    \I__2176\ : InMux
    port map (
            O => \N__11384\,
            I => \N__11381\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__11381\,
            I => \uart_inst0.uart_inst0.rx_countdown_s_1\
        );

    \I__2174\ : InMux
    port map (
            O => \N__11378\,
            I => \uart_inst0.uart_inst0.rx_countdown_cry_0\
        );

    \I__2173\ : InMux
    port map (
            O => \N__11375\,
            I => \N__11371\
        );

    \I__2172\ : InMux
    port map (
            O => \N__11374\,
            I => \N__11368\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__11371\,
            I => \uart_inst0.uart_inst0.rx_countdownZ0Z_2\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__11368\,
            I => \uart_inst0.uart_inst0.rx_countdownZ0Z_2\
        );

    \I__2169\ : InMux
    port map (
            O => \N__11363\,
            I => \N__11360\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__11360\,
            I => \uart_inst0.uart_inst0.rx_countdown_s_2\
        );

    \I__2167\ : InMux
    port map (
            O => \N__11357\,
            I => \uart_inst0.uart_inst0.rx_countdown_cry_1\
        );

    \I__2166\ : InMux
    port map (
            O => \N__11354\,
            I => \N__11350\
        );

    \I__2165\ : InMux
    port map (
            O => \N__11353\,
            I => \N__11347\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__11350\,
            I => \uart_inst0.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__11347\,
            I => \uart_inst0.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__2162\ : InMux
    port map (
            O => \N__11342\,
            I => \N__11339\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__11339\,
            I => \uart_inst0.uart_inst0.rx_countdown_s_3\
        );

    \I__2160\ : InMux
    port map (
            O => \N__11336\,
            I => \uart_inst0.uart_inst0.rx_countdown_cry_2\
        );

    \I__2159\ : InMux
    port map (
            O => \N__11333\,
            I => \N__11328\
        );

    \I__2158\ : InMux
    port map (
            O => \N__11332\,
            I => \N__11325\
        );

    \I__2157\ : InMux
    port map (
            O => \N__11331\,
            I => \N__11322\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__11328\,
            I => \uart_inst0.uart_inst0.rx_countdownZ0Z_4\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__11325\,
            I => \uart_inst0.uart_inst0.rx_countdownZ0Z_4\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__11322\,
            I => \uart_inst0.uart_inst0.rx_countdownZ0Z_4\
        );

    \I__2153\ : InMux
    port map (
            O => \N__11315\,
            I => \N__11311\
        );

    \I__2152\ : InMux
    port map (
            O => \N__11314\,
            I => \N__11308\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__11311\,
            I => \N__11305\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__11308\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ1Z_1\
        );

    \I__2149\ : Odrv4
    port map (
            O => \N__11305\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ1Z_1\
        );

    \I__2148\ : CascadeMux
    port map (
            O => \N__11300\,
            I => \N__11297\
        );

    \I__2147\ : InMux
    port map (
            O => \N__11297\,
            I => \N__11293\
        );

    \I__2146\ : InMux
    port map (
            O => \N__11296\,
            I => \N__11290\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__11293\,
            I => \N__11287\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__11290\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ0Z_2\
        );

    \I__2143\ : Odrv4
    port map (
            O => \N__11287\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ0Z_2\
        );

    \I__2142\ : CascadeMux
    port map (
            O => \N__11282\,
            I => \N__11279\
        );

    \I__2141\ : InMux
    port map (
            O => \N__11279\,
            I => \N__11276\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__11276\,
            I => \N__11270\
        );

    \I__2139\ : InMux
    port map (
            O => \N__11275\,
            I => \N__11267\
        );

    \I__2138\ : InMux
    port map (
            O => \N__11274\,
            I => \N__11262\
        );

    \I__2137\ : InMux
    port map (
            O => \N__11273\,
            I => \N__11262\
        );

    \I__2136\ : Odrv4
    port map (
            O => \N__11270\,
            I => \uart_inst0.uart_inst0.rx_stateZ0Z_5\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__11267\,
            I => \uart_inst0.uart_inst0.rx_stateZ0Z_5\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__11262\,
            I => \uart_inst0.uart_inst0.rx_stateZ0Z_5\
        );

    \I__2133\ : InMux
    port map (
            O => \N__11255\,
            I => \N__11252\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__11252\,
            I => \N__11249\
        );

    \I__2131\ : Odrv4
    port map (
            O => \N__11249\,
            I => \rUartRxDataZ0Z_0\
        );

    \I__2130\ : InMux
    port map (
            O => \N__11246\,
            I => \N__11231\
        );

    \I__2129\ : InMux
    port map (
            O => \N__11245\,
            I => \N__11231\
        );

    \I__2128\ : InMux
    port map (
            O => \N__11244\,
            I => \N__11231\
        );

    \I__2127\ : InMux
    port map (
            O => \N__11243\,
            I => \N__11231\
        );

    \I__2126\ : InMux
    port map (
            O => \N__11242\,
            I => \N__11231\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__11231\,
            I => \N__11225\
        );

    \I__2124\ : InMux
    port map (
            O => \N__11230\,
            I => \N__11218\
        );

    \I__2123\ : InMux
    port map (
            O => \N__11229\,
            I => \N__11218\
        );

    \I__2122\ : InMux
    port map (
            O => \N__11228\,
            I => \N__11218\
        );

    \I__2121\ : Span4Mux_h
    port map (
            O => \N__11225\,
            I => \N__11211\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__11218\,
            I => \N__11211\
        );

    \I__2119\ : InMux
    port map (
            O => \N__11217\,
            I => \N__11208\
        );

    \I__2118\ : InMux
    port map (
            O => \N__11216\,
            I => \N__11205\
        );

    \I__2117\ : Odrv4
    port map (
            O => \N__11211\,
            I => \rUartRxFlagZ0\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__11208\,
            I => \rUartRxFlagZ0\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__11205\,
            I => \rUartRxFlagZ0\
        );

    \I__2114\ : InMux
    port map (
            O => \N__11198\,
            I => \N__11195\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__11195\,
            I => \N__11192\
        );

    \I__2112\ : Span4Mux_v
    port map (
            O => \N__11192\,
            I => \N__11189\
        );

    \I__2111\ : Span4Mux_h
    port map (
            O => \N__11189\,
            I => \N__11186\
        );

    \I__2110\ : Odrv4
    port map (
            O => \N__11186\,
            I => \rUartTxDataZ0Z_0\
        );

    \I__2109\ : CEMux
    port map (
            O => \N__11183\,
            I => \N__11180\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__11180\,
            I => \N__11176\
        );

    \I__2107\ : CEMux
    port map (
            O => \N__11179\,
            I => \N__11173\
        );

    \I__2106\ : Odrv12
    port map (
            O => \N__11176\,
            I => \rUartTxEn_4_0\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__11173\,
            I => \rUartTxEn_4_0\
        );

    \I__2104\ : CEMux
    port map (
            O => \N__11168\,
            I => \N__11164\
        );

    \I__2103\ : CEMux
    port map (
            O => \N__11167\,
            I => \N__11161\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__11164\,
            I => \rUartRxState_0_0\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__11161\,
            I => \rUartRxState_0_0\
        );

    \I__2100\ : InMux
    port map (
            O => \N__11156\,
            I => \N__11152\
        );

    \I__2099\ : InMux
    port map (
            O => \N__11155\,
            I => \N__11148\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__11152\,
            I => \N__11145\
        );

    \I__2097\ : InMux
    port map (
            O => \N__11151\,
            I => \N__11142\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__11148\,
            I => \N__11139\
        );

    \I__2095\ : Span4Mux_v
    port map (
            O => \N__11145\,
            I => \N__11136\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__11142\,
            I => \N__11131\
        );

    \I__2093\ : Span4Mux_h
    port map (
            O => \N__11139\,
            I => \N__11131\
        );

    \I__2092\ : Span4Mux_v
    port map (
            O => \N__11136\,
            I => \N__11123\
        );

    \I__2091\ : Span4Mux_h
    port map (
            O => \N__11131\,
            I => \N__11123\
        );

    \I__2090\ : InMux
    port map (
            O => \N__11130\,
            I => \N__11118\
        );

    \I__2089\ : InMux
    port map (
            O => \N__11129\,
            I => \N__11118\
        );

    \I__2088\ : InMux
    port map (
            O => \N__11128\,
            I => \N__11115\
        );

    \I__2087\ : Odrv4
    port map (
            O => \N__11123\,
            I => \uart_inst0.uart_inst0.rx_stateZ0Z_0\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__11118\,
            I => \uart_inst0.uart_inst0.rx_stateZ0Z_0\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__11115\,
            I => \uart_inst0.uart_inst0.rx_stateZ0Z_0\
        );

    \I__2084\ : CascadeMux
    port map (
            O => \N__11108\,
            I => \N__11105\
        );

    \I__2083\ : InMux
    port map (
            O => \N__11105\,
            I => \N__11096\
        );

    \I__2082\ : InMux
    port map (
            O => \N__11104\,
            I => \N__11096\
        );

    \I__2081\ : InMux
    port map (
            O => \N__11103\,
            I => \N__11096\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__11096\,
            I => \uart_inst0.wRxWrEn_0\
        );

    \I__2079\ : CascadeMux
    port map (
            O => \N__11093\,
            I => \N__11090\
        );

    \I__2078\ : InMux
    port map (
            O => \N__11090\,
            I => \N__11087\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__11087\,
            I => \N__11084\
        );

    \I__2076\ : Span4Mux_h
    port map (
            O => \N__11084\,
            I => \N__11081\
        );

    \I__2075\ : Odrv4
    port map (
            O => \N__11081\,
            I => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_0_0\
        );

    \I__2074\ : InMux
    port map (
            O => \N__11078\,
            I => \N__11074\
        );

    \I__2073\ : InMux
    port map (
            O => \N__11077\,
            I => \N__11071\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__11074\,
            I => \N__11068\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__11071\,
            I => \fifo_inst_rx_fifo_inst_rRamRdAddr_5\
        );

    \I__2070\ : Odrv4
    port map (
            O => \N__11068\,
            I => \fifo_inst_rx_fifo_inst_rRamRdAddr_5\
        );

    \I__2069\ : InMux
    port map (
            O => \N__11063\,
            I => \N__11059\
        );

    \I__2068\ : InMux
    port map (
            O => \N__11062\,
            I => \N__11056\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__11059\,
            I => \fifo_inst_rx_fifo_inst_rRamRdAddr_4\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__11056\,
            I => \fifo_inst_rx_fifo_inst_rRamRdAddr_4\
        );

    \I__2065\ : InMux
    port map (
            O => \N__11051\,
            I => \N__11048\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__11048\,
            I => \N__11045\
        );

    \I__2063\ : Span4Mux_h
    port map (
            O => \N__11045\,
            I => \N__11041\
        );

    \I__2062\ : InMux
    port map (
            O => \N__11044\,
            I => \N__11038\
        );

    \I__2061\ : Odrv4
    port map (
            O => \N__11041\,
            I => \fifo_inst_rx_fifo_inst_rRamRdAddr_2\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__11038\,
            I => \fifo_inst_rx_fifo_inst_rRamRdAddr_2\
        );

    \I__2059\ : InMux
    port map (
            O => \N__11033\,
            I => \N__11029\
        );

    \I__2058\ : InMux
    port map (
            O => \N__11032\,
            I => \N__11026\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__11029\,
            I => \N__11023\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__11026\,
            I => \fifo_inst_rx_fifo_inst_rRamRdAddr_7\
        );

    \I__2055\ : Odrv4
    port map (
            O => \N__11023\,
            I => \fifo_inst_rx_fifo_inst_rRamRdAddr_7\
        );

    \I__2054\ : InMux
    port map (
            O => \N__11018\,
            I => \N__11014\
        );

    \I__2053\ : InMux
    port map (
            O => \N__11017\,
            I => \N__11011\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__11014\,
            I => \N__11008\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__11011\,
            I => \fifo_inst_rx_fifo_inst_rRamRdAddr_6\
        );

    \I__2050\ : Odrv4
    port map (
            O => \N__11008\,
            I => \fifo_inst_rx_fifo_inst_rRamRdAddr_6\
        );

    \I__2049\ : CascadeMux
    port map (
            O => \N__11003\,
            I => \uart_inst0.tx_uart_fifo_inst.m58_eZ0Z_5_cascade_\
        );

    \I__2048\ : InMux
    port map (
            O => \N__11000\,
            I => \N__10997\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__10997\,
            I => \uart_inst0.tx_uart_fifo_inst.m58_eZ0Z_6\
        );

    \I__2046\ : InMux
    port map (
            O => \N__10994\,
            I => \N__10989\
        );

    \I__2045\ : InMux
    port map (
            O => \N__10993\,
            I => \N__10986\
        );

    \I__2044\ : InMux
    port map (
            O => \N__10992\,
            I => \N__10983\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__10989\,
            I => \uart_inst0.tx_uart_fifo_inst.N_99\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__10986\,
            I => \uart_inst0.tx_uart_fifo_inst.N_99\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__10983\,
            I => \uart_inst0.tx_uart_fifo_inst.N_99\
        );

    \I__2040\ : InMux
    port map (
            O => \N__10976\,
            I => \N__10970\
        );

    \I__2039\ : InMux
    port map (
            O => \N__10975\,
            I => \N__10970\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__10970\,
            I => \rRamRdAddr_RNI0S8U_0\
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__10967\,
            I => \N__10963\
        );

    \I__2036\ : InMux
    port map (
            O => \N__10966\,
            I => \N__10958\
        );

    \I__2035\ : InMux
    port map (
            O => \N__10963\,
            I => \N__10955\
        );

    \I__2034\ : InMux
    port map (
            O => \N__10962\,
            I => \N__10951\
        );

    \I__2033\ : InMux
    port map (
            O => \N__10961\,
            I => \N__10948\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__10958\,
            I => \N__10943\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__10955\,
            I => \N__10943\
        );

    \I__2030\ : CascadeMux
    port map (
            O => \N__10954\,
            I => \N__10939\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__10951\,
            I => \N__10934\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__10948\,
            I => \N__10934\
        );

    \I__2027\ : Span4Mux_h
    port map (
            O => \N__10943\,
            I => \N__10931\
        );

    \I__2026\ : InMux
    port map (
            O => \N__10942\,
            I => \N__10928\
        );

    \I__2025\ : InMux
    port map (
            O => \N__10939\,
            I => \N__10925\
        );

    \I__2024\ : Odrv4
    port map (
            O => \N__10934\,
            I => \fifo_inst_rx_fifo_inst_wRamRdEn\
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__10931\,
            I => \fifo_inst_rx_fifo_inst_wRamRdEn\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__10928\,
            I => \fifo_inst_rx_fifo_inst_wRamRdEn\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__10925\,
            I => \fifo_inst_rx_fifo_inst_wRamRdEn\
        );

    \I__2020\ : CascadeMux
    port map (
            O => \N__10916\,
            I => \uart_inst0.tx_uart_fifo_inst.N_99_cascade_\
        );

    \I__2019\ : InMux
    port map (
            O => \N__10913\,
            I => \N__10909\
        );

    \I__2018\ : InMux
    port map (
            O => \N__10912\,
            I => \N__10906\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__10909\,
            I => \fifo_inst_rx_fifo_inst_rRamRdAddr_0\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__10906\,
            I => \fifo_inst_rx_fifo_inst_rRamRdAddr_0\
        );

    \I__2015\ : InMux
    port map (
            O => \N__10901\,
            I => \N__10898\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__10898\,
            I => \N__10895\
        );

    \I__2013\ : Odrv4
    port map (
            O => \N__10895\,
            I => \rUartRxDataZ0Z_3\
        );

    \I__2012\ : InMux
    port map (
            O => \N__10892\,
            I => \N__10889\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__10889\,
            I => \N__10886\
        );

    \I__2010\ : Span4Mux_v
    port map (
            O => \N__10886\,
            I => \N__10883\
        );

    \I__2009\ : Span4Mux_h
    port map (
            O => \N__10883\,
            I => \N__10880\
        );

    \I__2008\ : Odrv4
    port map (
            O => \N__10880\,
            I => \rUartTxDataZ0Z_3\
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__10877\,
            I => \N__10874\
        );

    \I__2006\ : InMux
    port map (
            O => \N__10874\,
            I => \N__10871\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__10871\,
            I => \N__10868\
        );

    \I__2004\ : Odrv4
    port map (
            O => \N__10868\,
            I => \rUartRxDataZ0Z_4\
        );

    \I__2003\ : InMux
    port map (
            O => \N__10865\,
            I => \N__10862\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__10862\,
            I => \rRxDataZ0Z_4\
        );

    \I__2001\ : InMux
    port map (
            O => \N__10859\,
            I => \N__10856\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__10856\,
            I => \N__10853\
        );

    \I__1999\ : Span4Mux_v
    port map (
            O => \N__10853\,
            I => \N__10850\
        );

    \I__1998\ : Odrv4
    port map (
            O => \N__10850\,
            I => \rUartTxDataZ0Z_4\
        );

    \I__1997\ : CascadeMux
    port map (
            O => \N__10847\,
            I => \N__10844\
        );

    \I__1996\ : InMux
    port map (
            O => \N__10844\,
            I => \N__10841\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__10841\,
            I => \rUartRxDataZ0Z_7\
        );

    \I__1994\ : InMux
    port map (
            O => \N__10838\,
            I => \N__10835\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__10835\,
            I => \N__10832\
        );

    \I__1992\ : Span4Mux_v
    port map (
            O => \N__10832\,
            I => \N__10829\
        );

    \I__1991\ : Odrv4
    port map (
            O => \N__10829\,
            I => \rUartTxDataZ0Z_7\
        );

    \I__1990\ : InMux
    port map (
            O => \N__10826\,
            I => \N__10823\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__10823\,
            I => \N__10820\
        );

    \I__1988\ : Odrv4
    port map (
            O => \N__10820\,
            I => \rUartRxDataZ0Z_2\
        );

    \I__1987\ : InMux
    port map (
            O => \N__10817\,
            I => \N__10814\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__10814\,
            I => \N__10811\
        );

    \I__1985\ : Span4Mux_v
    port map (
            O => \N__10811\,
            I => \N__10808\
        );

    \I__1984\ : Span4Mux_h
    port map (
            O => \N__10808\,
            I => \N__10805\
        );

    \I__1983\ : Odrv4
    port map (
            O => \N__10805\,
            I => \rUartTxDataZ0Z_2\
        );

    \I__1982\ : CascadeMux
    port map (
            O => \N__10802\,
            I => \N__10799\
        );

    \I__1981\ : InMux
    port map (
            O => \N__10799\,
            I => \N__10796\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__10796\,
            I => \N__10793\
        );

    \I__1979\ : Span4Mux_h
    port map (
            O => \N__10793\,
            I => \N__10789\
        );

    \I__1978\ : InMux
    port map (
            O => \N__10792\,
            I => \N__10786\
        );

    \I__1977\ : Odrv4
    port map (
            O => \N__10789\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIM36CZ0\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__10786\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIM36CZ0\
        );

    \I__1975\ : CascadeMux
    port map (
            O => \N__10781\,
            I => \N__10778\
        );

    \I__1974\ : InMux
    port map (
            O => \N__10778\,
            I => \N__10775\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__10775\,
            I => \N__10772\
        );

    \I__1972\ : Span4Mux_s2_v
    port map (
            O => \N__10772\,
            I => \N__10769\
        );

    \I__1971\ : Span4Mux_h
    port map (
            O => \N__10769\,
            I => \N__10765\
        );

    \I__1970\ : InMux
    port map (
            O => \N__10768\,
            I => \N__10762\
        );

    \I__1969\ : Odrv4
    port map (
            O => \N__10765\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIAHVBZ0\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__10762\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIAHVBZ0\
        );

    \I__1967\ : InMux
    port map (
            O => \N__10757\,
            I => \N__10751\
        );

    \I__1966\ : InMux
    port map (
            O => \N__10756\,
            I => \N__10751\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__10751\,
            I => \un1_rRamRdAddr_cry_2_c_RNII9N9\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__10748\,
            I => \N__10745\
        );

    \I__1963\ : InMux
    port map (
            O => \N__10745\,
            I => \N__10742\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__10742\,
            I => \N__10739\
        );

    \I__1961\ : Span4Mux_h
    port map (
            O => \N__10739\,
            I => \N__10736\
        );

    \I__1960\ : Odrv4
    port map (
            O => \N__10736\,
            I => m60
        );

    \I__1959\ : CascadeMux
    port map (
            O => \N__10733\,
            I => \N__10730\
        );

    \I__1958\ : InMux
    port map (
            O => \N__10730\,
            I => \N__10727\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__10727\,
            I => \N__10724\
        );

    \I__1956\ : Span4Mux_h
    port map (
            O => \N__10724\,
            I => \N__10720\
        );

    \I__1955\ : InMux
    port map (
            O => \N__10723\,
            I => \N__10717\
        );

    \I__1954\ : Odrv4
    port map (
            O => \N__10720\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIGQ2CZ0\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__10717\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIGQ2CZ0\
        );

    \I__1952\ : InMux
    port map (
            O => \N__10712\,
            I => \N__10708\
        );

    \I__1951\ : InMux
    port map (
            O => \N__10711\,
            I => \N__10705\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__10708\,
            I => \fifo_inst_rx_fifo_inst_rRamRdAddr_3\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__10705\,
            I => \fifo_inst_rx_fifo_inst_rRamRdAddr_3\
        );

    \I__1948\ : InMux
    port map (
            O => \N__10700\,
            I => \N__10696\
        );

    \I__1947\ : InMux
    port map (
            O => \N__10699\,
            I => \N__10693\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__10696\,
            I => \fifo_inst_rx_fifo_inst_rRamRdAddr_1\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__10693\,
            I => \fifo_inst_rx_fifo_inst_rRamRdAddr_1\
        );

    \I__1944\ : CascadeMux
    port map (
            O => \N__10688\,
            I => \N__10684\
        );

    \I__1943\ : InMux
    port map (
            O => \N__10687\,
            I => \N__10681\
        );

    \I__1942\ : InMux
    port map (
            O => \N__10684\,
            I => \N__10678\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__10681\,
            I => \fifo_inst_rx_fifo_inst_rRamRdAddr_8\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__10678\,
            I => \fifo_inst_rx_fifo_inst_rRamRdAddr_8\
        );

    \I__1939\ : InMux
    port map (
            O => \N__10673\,
            I => \N__10669\
        );

    \I__1938\ : InMux
    port map (
            O => \N__10672\,
            I => \N__10666\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__10669\,
            I => \N__10663\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__10666\,
            I => \N_101\
        );

    \I__1935\ : Odrv4
    port map (
            O => \N__10663\,
            I => \N_101\
        );

    \I__1934\ : InMux
    port map (
            O => \N__10658\,
            I => \N__10653\
        );

    \I__1933\ : InMux
    port map (
            O => \N__10657\,
            I => \N__10649\
        );

    \I__1932\ : InMux
    port map (
            O => \N__10656\,
            I => \N__10646\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__10653\,
            I => \N__10643\
        );

    \I__1930\ : InMux
    port map (
            O => \N__10652\,
            I => \N__10640\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__10649\,
            I => \N__10637\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__10646\,
            I => \N__10633\
        );

    \I__1927\ : Span4Mux_v
    port map (
            O => \N__10643\,
            I => \N__10628\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__10640\,
            I => \N__10628\
        );

    \I__1925\ : Span4Mux_v
    port map (
            O => \N__10637\,
            I => \N__10625\
        );

    \I__1924\ : InMux
    port map (
            O => \N__10636\,
            I => \N__10622\
        );

    \I__1923\ : Odrv4
    port map (
            O => \N__10633\,
            I => \N_97\
        );

    \I__1922\ : Odrv4
    port map (
            O => \N__10628\,
            I => \N_97\
        );

    \I__1921\ : Odrv4
    port map (
            O => \N__10625\,
            I => \N_97\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__10622\,
            I => \N_97\
        );

    \I__1919\ : CascadeMux
    port map (
            O => \N__10613\,
            I => \N__10610\
        );

    \I__1918\ : InMux
    port map (
            O => \N__10610\,
            I => \N__10604\
        );

    \I__1917\ : InMux
    port map (
            O => \N__10609\,
            I => \N__10601\
        );

    \I__1916\ : InMux
    port map (
            O => \N__10608\,
            I => \N__10597\
        );

    \I__1915\ : InMux
    port map (
            O => \N__10607\,
            I => \N__10594\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__10604\,
            I => \N__10588\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__10601\,
            I => \N__10588\
        );

    \I__1912\ : InMux
    port map (
            O => \N__10600\,
            I => \N__10585\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__10597\,
            I => \N__10582\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__10594\,
            I => \N__10579\
        );

    \I__1909\ : CascadeMux
    port map (
            O => \N__10593\,
            I => \N__10576\
        );

    \I__1908\ : Span4Mux_v
    port map (
            O => \N__10588\,
            I => \N__10571\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__10585\,
            I => \N__10571\
        );

    \I__1906\ : Span4Mux_v
    port map (
            O => \N__10582\,
            I => \N__10566\
        );

    \I__1905\ : Span4Mux_v
    port map (
            O => \N__10579\,
            I => \N__10566\
        );

    \I__1904\ : InMux
    port map (
            O => \N__10576\,
            I => \N__10563\
        );

    \I__1903\ : Span4Mux_v
    port map (
            O => \N__10571\,
            I => \N__10560\
        );

    \I__1902\ : Sp12to4
    port map (
            O => \N__10566\,
            I => \N__10555\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__10563\,
            I => \N__10555\
        );

    \I__1900\ : Span4Mux_h
    port map (
            O => \N__10560\,
            I => \N__10552\
        );

    \I__1899\ : Span12Mux_h
    port map (
            O => \N__10555\,
            I => \N__10549\
        );

    \I__1898\ : Sp12to4
    port map (
            O => \N__10552\,
            I => \N__10546\
        );

    \I__1897\ : Span12Mux_v
    port map (
            O => \N__10549\,
            I => \N__10543\
        );

    \I__1896\ : Span12Mux_v
    port map (
            O => \N__10546\,
            I => \N__10540\
        );

    \I__1895\ : Span12Mux_v
    port map (
            O => \N__10543\,
            I => \N__10537\
        );

    \I__1894\ : Odrv12
    port map (
            O => \N__10540\,
            I => \iTxE_n_c\
        );

    \I__1893\ : Odrv12
    port map (
            O => \N__10537\,
            I => \iTxE_n_c\
        );

    \I__1892\ : InMux
    port map (
            O => \N__10532\,
            I => \N__10527\
        );

    \I__1891\ : InMux
    port map (
            O => \N__10531\,
            I => \N__10520\
        );

    \I__1890\ : InMux
    port map (
            O => \N__10530\,
            I => \N__10517\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__10527\,
            I => \N__10514\
        );

    \I__1888\ : InMux
    port map (
            O => \N__10526\,
            I => \N__10511\
        );

    \I__1887\ : InMux
    port map (
            O => \N__10525\,
            I => \N__10508\
        );

    \I__1886\ : InMux
    port map (
            O => \N__10524\,
            I => \N__10503\
        );

    \I__1885\ : InMux
    port map (
            O => \N__10523\,
            I => \N__10503\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__10520\,
            I => \N__10500\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__10517\,
            I => \N__10496\
        );

    \I__1882\ : Span4Mux_h
    port map (
            O => \N__10514\,
            I => \N__10491\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__10511\,
            I => \N__10491\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__10508\,
            I => \N__10484\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__10503\,
            I => \N__10484\
        );

    \I__1878\ : Span4Mux_h
    port map (
            O => \N__10500\,
            I => \N__10484\
        );

    \I__1877\ : InMux
    port map (
            O => \N__10499\,
            I => \N__10481\
        );

    \I__1876\ : Odrv4
    port map (
            O => \N__10496\,
            I => \N_8_0\
        );

    \I__1875\ : Odrv4
    port map (
            O => \N__10491\,
            I => \N_8_0\
        );

    \I__1874\ : Odrv4
    port map (
            O => \N__10484\,
            I => \N_8_0\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__10481\,
            I => \N_8_0\
        );

    \I__1872\ : CascadeMux
    port map (
            O => \N__10472\,
            I => \fifo_inst_ft2232h_inst_un1_rFifoState_1_sqmuxa_0_i_cascade_\
        );

    \I__1871\ : CEMux
    port map (
            O => \N__10469\,
            I => \N__10466\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__10466\,
            I => \N__10463\
        );

    \I__1869\ : Odrv4
    port map (
            O => \N__10463\,
            I => \fifo_inst.ft2232h_inst.un1_rFifoState_1_sqmuxa_0_i_0\
        );

    \I__1868\ : CascadeMux
    port map (
            O => \N__10460\,
            I => \N__10457\
        );

    \I__1867\ : InMux
    port map (
            O => \N__10457\,
            I => \N__10454\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__10454\,
            I => \N__10451\
        );

    \I__1865\ : Span4Mux_h
    port map (
            O => \N__10451\,
            I => \N__10448\
        );

    \I__1864\ : Odrv4
    port map (
            O => \N__10448\,
            I => m59
        );

    \I__1863\ : CascadeMux
    port map (
            O => \N__10445\,
            I => \N__10442\
        );

    \I__1862\ : InMux
    port map (
            O => \N__10442\,
            I => \N__10436\
        );

    \I__1861\ : InMux
    port map (
            O => \N__10441\,
            I => \N__10436\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__10436\,
            I => \un1_rRamRdAddr_cry_2_c_RNIMVKN\
        );

    \I__1859\ : CascadeMux
    port map (
            O => \N__10433\,
            I => \N__10430\
        );

    \I__1858\ : InMux
    port map (
            O => \N__10430\,
            I => \N__10427\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__10427\,
            I => \N__10424\
        );

    \I__1856\ : Span4Mux_s2_v
    port map (
            O => \N__10424\,
            I => \N__10421\
        );

    \I__1855\ : Odrv4
    port map (
            O => \N__10421\,
            I => m74
        );

    \I__1854\ : InMux
    port map (
            O => \N__10418\,
            I => \N__10414\
        );

    \I__1853\ : InMux
    port map (
            O => \N__10417\,
            I => \N__10411\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__10414\,
            I => \fifo_inst_tx_fifo_inst_rRamRdAddr_5\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__10411\,
            I => \fifo_inst_tx_fifo_inst_rRamRdAddr_5\
        );

    \I__1850\ : InMux
    port map (
            O => \N__10406\,
            I => \N__10402\
        );

    \I__1849\ : InMux
    port map (
            O => \N__10405\,
            I => \N__10399\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__10402\,
            I => \fifo_inst_tx_fifo_inst_rRamRdAddr_7\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__10399\,
            I => \fifo_inst_tx_fifo_inst_rRamRdAddr_7\
        );

    \I__1846\ : InMux
    port map (
            O => \N__10394\,
            I => \N__10390\
        );

    \I__1845\ : InMux
    port map (
            O => \N__10393\,
            I => \N__10387\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__10390\,
            I => \fifo_inst_tx_fifo_inst_rRamRdAddr_6\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__10387\,
            I => \fifo_inst_tx_fifo_inst_rRamRdAddr_6\
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__10382\,
            I => \uart_inst0.tx_uart_fifo_inst.m72_eZ0Z_5_cascade_\
        );

    \I__1841\ : CascadeMux
    port map (
            O => \N__10379\,
            I => \uart_inst0.tx_uart_fifo_inst.N_100_cascade_\
        );

    \I__1840\ : CascadeMux
    port map (
            O => \N__10376\,
            I => \N__10373\
        );

    \I__1839\ : InMux
    port map (
            O => \N__10373\,
            I => \N__10370\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__10370\,
            I => \N__10367\
        );

    \I__1837\ : Span4Mux_s2_v
    port map (
            O => \N__10367\,
            I => \N__10364\
        );

    \I__1836\ : Odrv4
    port map (
            O => \N__10364\,
            I => m73
        );

    \I__1835\ : InMux
    port map (
            O => \N__10361\,
            I => \N__10357\
        );

    \I__1834\ : InMux
    port map (
            O => \N__10360\,
            I => \N__10354\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__10357\,
            I => \fifo_inst_tx_fifo_inst_rRamRdAddr_3\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__10354\,
            I => \fifo_inst_tx_fifo_inst_rRamRdAddr_3\
        );

    \I__1831\ : InMux
    port map (
            O => \N__10349\,
            I => \N__10345\
        );

    \I__1830\ : InMux
    port map (
            O => \N__10348\,
            I => \N__10342\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__10345\,
            I => \fifo_inst_tx_fifo_inst_rRamRdAddr_1\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__10342\,
            I => \fifo_inst_tx_fifo_inst_rRamRdAddr_1\
        );

    \I__1827\ : CascadeMux
    port map (
            O => \N__10337\,
            I => \N__10334\
        );

    \I__1826\ : InMux
    port map (
            O => \N__10334\,
            I => \N__10330\
        );

    \I__1825\ : InMux
    port map (
            O => \N__10333\,
            I => \N__10327\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__10330\,
            I => \N__10324\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__10327\,
            I => \fifo_inst_tx_fifo_inst_rRamRdAddr_8\
        );

    \I__1822\ : Odrv4
    port map (
            O => \N__10324\,
            I => \fifo_inst_tx_fifo_inst_rRamRdAddr_8\
        );

    \I__1821\ : InMux
    port map (
            O => \N__10319\,
            I => \N__10316\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__10316\,
            I => \uart_inst0.tx_uart_fifo_inst.m72_eZ0Z_6\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__10313\,
            I => \N__10310\
        );

    \I__1818\ : InMux
    port map (
            O => \N__10310\,
            I => \N__10307\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__10307\,
            I => \N__10304\
        );

    \I__1816\ : Span4Mux_s2_v
    port map (
            O => \N__10304\,
            I => \N__10300\
        );

    \I__1815\ : InMux
    port map (
            O => \N__10303\,
            I => \N__10297\
        );

    \I__1814\ : Odrv4
    port map (
            O => \N__10300\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIKG0QZ0\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__10297\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIKG0QZ0\
        );

    \I__1812\ : InMux
    port map (
            O => \N__10292\,
            I => \N__10288\
        );

    \I__1811\ : InMux
    port map (
            O => \N__10291\,
            I => \N__10285\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__10288\,
            I => \fifo_inst_tx_fifo_inst_rRamRdAddr_4\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__10285\,
            I => \fifo_inst_tx_fifo_inst_rRamRdAddr_4\
        );

    \I__1808\ : InMux
    port map (
            O => \N__10280\,
            I => \N__10266\
        );

    \I__1807\ : InMux
    port map (
            O => \N__10279\,
            I => \N__10266\
        );

    \I__1806\ : InMux
    port map (
            O => \N__10278\,
            I => \N__10266\
        );

    \I__1805\ : InMux
    port map (
            O => \N__10277\,
            I => \N__10266\
        );

    \I__1804\ : CEMux
    port map (
            O => \N__10276\,
            I => \N__10262\
        );

    \I__1803\ : CascadeMux
    port map (
            O => \N__10275\,
            I => \N__10259\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__10266\,
            I => \N__10256\
        );

    \I__1801\ : InMux
    port map (
            O => \N__10265\,
            I => \N__10253\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__10262\,
            I => \N__10250\
        );

    \I__1799\ : InMux
    port map (
            O => \N__10259\,
            I => \N__10247\
        );

    \I__1798\ : Odrv4
    port map (
            O => \N__10256\,
            I => \fifo_inst_tx_fifo_inst_wRamRdEn\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__10253\,
            I => \fifo_inst_tx_fifo_inst_wRamRdEn\
        );

    \I__1796\ : Odrv4
    port map (
            O => \N__10250\,
            I => \fifo_inst_tx_fifo_inst_wRamRdEn\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__10247\,
            I => \fifo_inst_tx_fifo_inst_wRamRdEn\
        );

    \I__1794\ : CascadeMux
    port map (
            O => \N__10238\,
            I => \N__10235\
        );

    \I__1793\ : InMux
    port map (
            O => \N__10235\,
            I => \N__10229\
        );

    \I__1792\ : InMux
    port map (
            O => \N__10234\,
            I => \N__10229\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__10229\,
            I => \rRamRdAddr_RNI9KL42_0\
        );

    \I__1790\ : InMux
    port map (
            O => \N__10226\,
            I => \N__10217\
        );

    \I__1789\ : InMux
    port map (
            O => \N__10225\,
            I => \N__10217\
        );

    \I__1788\ : InMux
    port map (
            O => \N__10224\,
            I => \N__10217\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__10217\,
            I => \uart_inst0.tx_uart_fifo_inst.N_100\
        );

    \I__1786\ : InMux
    port map (
            O => \N__10214\,
            I => \N__10210\
        );

    \I__1785\ : InMux
    port map (
            O => \N__10213\,
            I => \N__10207\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__10210\,
            I => \fifo_inst_tx_fifo_inst_rRamRdAddr_0\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__10207\,
            I => \fifo_inst_tx_fifo_inst_rRamRdAddr_0\
        );

    \I__1782\ : CascadeMux
    port map (
            O => \N__10202\,
            I => \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_11_3_cascade_\
        );

    \I__1781\ : InMux
    port map (
            O => \N__10199\,
            I => \N__10191\
        );

    \I__1780\ : InMux
    port map (
            O => \N__10198\,
            I => \N__10191\
        );

    \I__1779\ : InMux
    port map (
            O => \N__10197\,
            I => \N__10188\
        );

    \I__1778\ : InMux
    port map (
            O => \N__10196\,
            I => \N__10185\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__10191\,
            I => \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__10188\,
            I => \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__10185\,
            I => \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__10178\,
            I => \N__10175\
        );

    \I__1773\ : InMux
    port map (
            O => \N__10175\,
            I => \N__10170\
        );

    \I__1772\ : InMux
    port map (
            O => \N__10174\,
            I => \N__10167\
        );

    \I__1771\ : InMux
    port map (
            O => \N__10173\,
            I => \N__10164\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__10170\,
            I => \N__10157\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__10167\,
            I => \N__10154\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__10164\,
            I => \N__10151\
        );

    \I__1767\ : InMux
    port map (
            O => \N__10163\,
            I => \N__10148\
        );

    \I__1766\ : CascadeMux
    port map (
            O => \N__10162\,
            I => \N__10144\
        );

    \I__1765\ : InMux
    port map (
            O => \N__10161\,
            I => \N__10138\
        );

    \I__1764\ : InMux
    port map (
            O => \N__10160\,
            I => \N__10138\
        );

    \I__1763\ : Span4Mux_h
    port map (
            O => \N__10157\,
            I => \N__10135\
        );

    \I__1762\ : Span12Mux_h
    port map (
            O => \N__10154\,
            I => \N__10132\
        );

    \I__1761\ : Span4Mux_h
    port map (
            O => \N__10151\,
            I => \N__10127\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__10148\,
            I => \N__10127\
        );

    \I__1759\ : InMux
    port map (
            O => \N__10147\,
            I => \N__10122\
        );

    \I__1758\ : InMux
    port map (
            O => \N__10144\,
            I => \N__10122\
        );

    \I__1757\ : InMux
    port map (
            O => \N__10143\,
            I => \N__10119\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__10138\,
            I => \wTxFull\
        );

    \I__1755\ : Odrv4
    port map (
            O => \N__10135\,
            I => \wTxFull\
        );

    \I__1754\ : Odrv12
    port map (
            O => \N__10132\,
            I => \wTxFull\
        );

    \I__1753\ : Odrv4
    port map (
            O => \N__10127\,
            I => \wTxFull\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__10122\,
            I => \wTxFull\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__10119\,
            I => \wTxFull\
        );

    \I__1750\ : InMux
    port map (
            O => \N__10106\,
            I => \N__10103\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__10103\,
            I => \N__10099\
        );

    \I__1748\ : InMux
    port map (
            O => \N__10102\,
            I => \N__10096\
        );

    \I__1747\ : Span12Mux_v
    port map (
            O => \N__10099\,
            I => \N__10093\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__10096\,
            I => \rTxDataZ0Z_0\
        );

    \I__1745\ : Odrv12
    port map (
            O => \N__10093\,
            I => \rTxDataZ0Z_0\
        );

    \I__1744\ : IoInMux
    port map (
            O => \N__10088\,
            I => \N__10084\
        );

    \I__1743\ : IoInMux
    port map (
            O => \N__10087\,
            I => \N__10081\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__10084\,
            I => \N__10076\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__10081\,
            I => \N__10076\
        );

    \I__1740\ : IoSpan4Mux
    port map (
            O => \N__10076\,
            I => \N__10072\
        );

    \I__1739\ : IoInMux
    port map (
            O => \N__10075\,
            I => \N__10069\
        );

    \I__1738\ : Span4Mux_s3_v
    port map (
            O => \N__10072\,
            I => \N__10065\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__10069\,
            I => \N__10061\
        );

    \I__1736\ : IoInMux
    port map (
            O => \N__10068\,
            I => \N__10058\
        );

    \I__1735\ : Sp12to4
    port map (
            O => \N__10065\,
            I => \N__10052\
        );

    \I__1734\ : IoInMux
    port map (
            O => \N__10064\,
            I => \N__10049\
        );

    \I__1733\ : IoSpan4Mux
    port map (
            O => \N__10061\,
            I => \N__10044\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__10058\,
            I => \N__10044\
        );

    \I__1731\ : IoInMux
    port map (
            O => \N__10057\,
            I => \N__10041\
        );

    \I__1730\ : IoInMux
    port map (
            O => \N__10056\,
            I => \N__10038\
        );

    \I__1729\ : IoInMux
    port map (
            O => \N__10055\,
            I => \N__10035\
        );

    \I__1728\ : Span12Mux_v
    port map (
            O => \N__10052\,
            I => \N__10032\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__10049\,
            I => \N__10029\
        );

    \I__1726\ : IoSpan4Mux
    port map (
            O => \N__10044\,
            I => \N__10024\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__10041\,
            I => \N__10024\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__10038\,
            I => \N__10021\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__10035\,
            I => \N__10018\
        );

    \I__1722\ : Span12Mux_v
    port map (
            O => \N__10032\,
            I => \N__10015\
        );

    \I__1721\ : Span4Mux_s1_v
    port map (
            O => \N__10029\,
            I => \N__10012\
        );

    \I__1720\ : Span4Mux_s1_v
    port map (
            O => \N__10024\,
            I => \N__10009\
        );

    \I__1719\ : Span4Mux_s1_v
    port map (
            O => \N__10021\,
            I => \N__10004\
        );

    \I__1718\ : Span4Mux_s1_v
    port map (
            O => \N__10018\,
            I => \N__10004\
        );

    \I__1717\ : Odrv12
    port map (
            O => \N__10015\,
            I => \rTxBusReady\
        );

    \I__1716\ : Odrv4
    port map (
            O => \N__10012\,
            I => \rTxBusReady\
        );

    \I__1715\ : Odrv4
    port map (
            O => \N__10009\,
            I => \rTxBusReady\
        );

    \I__1714\ : Odrv4
    port map (
            O => \N__10004\,
            I => \rTxBusReady\
        );

    \I__1713\ : CascadeMux
    port map (
            O => \N__9995\,
            I => \uart_inst0.uart_inst0.tx_state_ns_0_0_0_cascade_\
        );

    \I__1712\ : InMux
    port map (
            O => \N__9992\,
            I => \N__9989\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__9989\,
            I => \N__9985\
        );

    \I__1710\ : InMux
    port map (
            O => \N__9988\,
            I => \N__9982\
        );

    \I__1709\ : Odrv4
    port map (
            O => \N__9985\,
            I => \uart_inst0.uart_inst0.tx_state_1_sqmuxa_1_0_a3_0\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__9982\,
            I => \uart_inst0.uart_inst0.tx_state_1_sqmuxa_1_0_a3_0\
        );

    \I__1707\ : SRMux
    port map (
            O => \N__9977\,
            I => \N__9974\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__9974\,
            I => \N__9971\
        );

    \I__1705\ : Span4Mux_h
    port map (
            O => \N__9971\,
            I => \N__9967\
        );

    \I__1704\ : InMux
    port map (
            O => \N__9970\,
            I => \N__9964\
        );

    \I__1703\ : Odrv4
    port map (
            O => \N__9967\,
            I => \uart_inst0.uart_inst0.tx_state_RNI1319Z0Z_0\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__9964\,
            I => \uart_inst0.uart_inst0.tx_state_RNI1319Z0Z_0\
        );

    \I__1701\ : InMux
    port map (
            O => \N__9959\,
            I => \N__9952\
        );

    \I__1700\ : InMux
    port map (
            O => \N__9958\,
            I => \N__9947\
        );

    \I__1699\ : InMux
    port map (
            O => \N__9957\,
            I => \N__9947\
        );

    \I__1698\ : InMux
    port map (
            O => \N__9956\,
            I => \N__9944\
        );

    \I__1697\ : InMux
    port map (
            O => \N__9955\,
            I => \N__9941\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__9952\,
            I => \N__9938\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__9947\,
            I => \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_1\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__9944\,
            I => \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_1\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__9941\,
            I => \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_1\
        );

    \I__1692\ : Odrv4
    port map (
            O => \N__9938\,
            I => \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_1\
        );

    \I__1691\ : InMux
    port map (
            O => \N__9929\,
            I => \N__9918\
        );

    \I__1690\ : InMux
    port map (
            O => \N__9928\,
            I => \N__9918\
        );

    \I__1689\ : InMux
    port map (
            O => \N__9927\,
            I => \N__9918\
        );

    \I__1688\ : InMux
    port map (
            O => \N__9926\,
            I => \N__9915\
        );

    \I__1687\ : InMux
    port map (
            O => \N__9925\,
            I => \N__9912\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__9918\,
            I => \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_0\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__9915\,
            I => \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_0\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__9912\,
            I => \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_0\
        );

    \I__1683\ : CascadeMux
    port map (
            O => \N__9905\,
            I => \uart_inst0.uart_inst0.un1_tx_bits_remaining_ac0_1_a0_0_cascade_\
        );

    \I__1682\ : InMux
    port map (
            O => \N__9902\,
            I => \N__9899\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__9899\,
            I => \uart_inst0.uart_inst0.un1_tx_bits_remaining_ac0_1\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__9896\,
            I => \uart_inst0.uart_inst0.un1_rx_state49_i_cascade_\
        );

    \I__1679\ : CascadeMux
    port map (
            O => \N__9893\,
            I => \uart_inst0.uart_inst0.tx_countdown_RNO_0Z0Z_3_cascade_\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__9890\,
            I => \uart_inst0.uart_inst0.N_147_0_cascade_\
        );

    \I__1677\ : CascadeMux
    port map (
            O => \N__9887\,
            I => \uart_inst0.uart_inst0.N_277_cascade_\
        );

    \I__1676\ : InMux
    port map (
            O => \N__9884\,
            I => \N__9881\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__9881\,
            I => \uart_inst0.uart_inst0.rx_state_srsts_0_a5_1_0\
        );

    \I__1674\ : CascadeMux
    port map (
            O => \N__9878\,
            I => \uart_inst0.uart_inst0.N_280_cascade_\
        );

    \I__1673\ : InMux
    port map (
            O => \N__9875\,
            I => \N__9870\
        );

    \I__1672\ : InMux
    port map (
            O => \N__9874\,
            I => \N__9865\
        );

    \I__1671\ : InMux
    port map (
            O => \N__9873\,
            I => \N__9865\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__9870\,
            I => \uart_inst0.uart_inst0.rx_stateZ0Z_4\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__9865\,
            I => \uart_inst0.uart_inst0.rx_stateZ0Z_4\
        );

    \I__1668\ : InMux
    port map (
            O => \N__9860\,
            I => \N__9857\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__9857\,
            I => \uart_inst0.uart_inst0.N_261_0\
        );

    \I__1666\ : InMux
    port map (
            O => \N__9854\,
            I => \N__9851\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__9851\,
            I => \N__9845\
        );

    \I__1664\ : CascadeMux
    port map (
            O => \N__9850\,
            I => \N__9842\
        );

    \I__1663\ : InMux
    port map (
            O => \N__9849\,
            I => \N__9839\
        );

    \I__1662\ : CascadeMux
    port map (
            O => \N__9848\,
            I => \N__9836\
        );

    \I__1661\ : Span4Mux_h
    port map (
            O => \N__9845\,
            I => \N__9833\
        );

    \I__1660\ : InMux
    port map (
            O => \N__9842\,
            I => \N__9829\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__9839\,
            I => \N__9826\
        );

    \I__1658\ : InMux
    port map (
            O => \N__9836\,
            I => \N__9823\
        );

    \I__1657\ : Span4Mux_v
    port map (
            O => \N__9833\,
            I => \N__9820\
        );

    \I__1656\ : InMux
    port map (
            O => \N__9832\,
            I => \N__9817\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__9829\,
            I => \N__9814\
        );

    \I__1654\ : Odrv4
    port map (
            O => \N__9826\,
            I => \uart_inst0.wTxRdEmpty\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__9823\,
            I => \uart_inst0.wTxRdEmpty\
        );

    \I__1652\ : Odrv4
    port map (
            O => \N__9820\,
            I => \uart_inst0.wTxRdEmpty\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__9817\,
            I => \uart_inst0.wTxRdEmpty\
        );

    \I__1650\ : Odrv12
    port map (
            O => \N__9814\,
            I => \uart_inst0.wTxRdEmpty\
        );

    \I__1649\ : CascadeMux
    port map (
            O => \N__9803\,
            I => \uart_inst0.uart_inst0.rx_state_srsts_0_o2_3_3_cascade_\
        );

    \I__1648\ : CascadeMux
    port map (
            O => \N__9800\,
            I => \uart_inst0.uart_inst0.N_257_0_cascade_\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__9797\,
            I => \N__9793\
        );

    \I__1646\ : InMux
    port map (
            O => \N__9796\,
            I => \N__9789\
        );

    \I__1645\ : InMux
    port map (
            O => \N__9793\,
            I => \N__9786\
        );

    \I__1644\ : InMux
    port map (
            O => \N__9792\,
            I => \N__9783\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__9789\,
            I => \N__9780\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__9786\,
            I => \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_2\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__9783\,
            I => \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_2\
        );

    \I__1640\ : Odrv4
    port map (
            O => \N__9780\,
            I => \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_2\
        );

    \I__1639\ : CascadeMux
    port map (
            O => \N__9773\,
            I => \N__9770\
        );

    \I__1638\ : InMux
    port map (
            O => \N__9770\,
            I => \N__9767\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__9767\,
            I => \N__9763\
        );

    \I__1636\ : InMux
    port map (
            O => \N__9766\,
            I => \N__9760\
        );

    \I__1635\ : Span4Mux_h
    port map (
            O => \N__9763\,
            I => \N__9757\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__9760\,
            I => \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_3\
        );

    \I__1633\ : Odrv4
    port map (
            O => \N__9757\,
            I => \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_3\
        );

    \I__1632\ : CascadeMux
    port map (
            O => \N__9752\,
            I => \N__9749\
        );

    \I__1631\ : InMux
    port map (
            O => \N__9749\,
            I => \N__9743\
        );

    \I__1630\ : InMux
    port map (
            O => \N__9748\,
            I => \N__9743\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__9743\,
            I => \uart_inst0.uart_inst0.N_157\
        );

    \I__1628\ : CascadeMux
    port map (
            O => \N__9740\,
            I => \uart_inst0.uart_inst0.N_157_cascade_\
        );

    \I__1627\ : CascadeMux
    port map (
            O => \N__9737\,
            I => \N__9734\
        );

    \I__1626\ : InMux
    port map (
            O => \N__9734\,
            I => \N__9731\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__9731\,
            I => \N__9728\
        );

    \I__1624\ : Odrv12
    port map (
            O => \N__9728\,
            I => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_3\
        );

    \I__1623\ : InMux
    port map (
            O => \N__9725\,
            I => \N__9721\
        );

    \I__1622\ : InMux
    port map (
            O => \N__9724\,
            I => \N__9718\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__9721\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIUJZ0Z84\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__9718\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIUJZ0Z84\
        );

    \I__1619\ : InMux
    port map (
            O => \N__9713\,
            I => \N__9710\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__9710\,
            I => \N__9706\
        );

    \I__1617\ : InMux
    port map (
            O => \N__9709\,
            I => \N__9703\
        );

    \I__1616\ : Odrv4
    port map (
            O => \N__9706\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_4\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__9703\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_4\
        );

    \I__1614\ : InMux
    port map (
            O => \N__9698\,
            I => \N__9695\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__9695\,
            I => \N__9691\
        );

    \I__1612\ : InMux
    port map (
            O => \N__9694\,
            I => \N__9688\
        );

    \I__1611\ : Odrv4
    port map (
            O => \N__9691\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_5\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__9688\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_5\
        );

    \I__1609\ : InMux
    port map (
            O => \N__9683\,
            I => \N__9679\
        );

    \I__1608\ : InMux
    port map (
            O => \N__9682\,
            I => \N__9676\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__9679\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNI2QAZ0Z4\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__9676\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNI2QAZ0Z4\
        );

    \I__1605\ : InMux
    port map (
            O => \N__9671\,
            I => \N__9668\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__9668\,
            I => \N__9664\
        );

    \I__1603\ : InMux
    port map (
            O => \N__9667\,
            I => \N__9661\
        );

    \I__1602\ : Odrv4
    port map (
            O => \N__9664\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_6\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__9661\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_6\
        );

    \I__1600\ : InMux
    port map (
            O => \N__9656\,
            I => \N__9652\
        );

    \I__1599\ : InMux
    port map (
            O => \N__9655\,
            I => \N__9649\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__9652\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI4TBZ0Z4\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__9649\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI4TBZ0Z4\
        );

    \I__1596\ : CascadeMux
    port map (
            O => \N__9644\,
            I => \N__9641\
        );

    \I__1595\ : InMux
    port map (
            O => \N__9641\,
            I => \N__9638\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__9638\,
            I => \N__9635\
        );

    \I__1593\ : Span4Mux_v
    port map (
            O => \N__9635\,
            I => \N__9631\
        );

    \I__1592\ : InMux
    port map (
            O => \N__9634\,
            I => \N__9628\
        );

    \I__1591\ : Odrv4
    port map (
            O => \N__9631\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_7\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__9628\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_7\
        );

    \I__1589\ : InMux
    port map (
            O => \N__9623\,
            I => \N__9619\
        );

    \I__1588\ : InMux
    port map (
            O => \N__9622\,
            I => \N__9616\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__9619\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI60DZ0Z4\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__9616\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI60DZ0Z4\
        );

    \I__1585\ : InMux
    port map (
            O => \N__9611\,
            I => \N__9607\
        );

    \I__1584\ : InMux
    port map (
            O => \N__9610\,
            I => \N__9604\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__9607\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_8\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__9604\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_8\
        );

    \I__1581\ : CascadeMux
    port map (
            O => \N__9599\,
            I => \uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_5_cascade_\
        );

    \I__1580\ : CascadeMux
    port map (
            O => \N__9596\,
            I => \uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7_cascade_\
        );

    \I__1579\ : CEMux
    port map (
            O => \N__9593\,
            I => \N__9584\
        );

    \I__1578\ : CascadeMux
    port map (
            O => \N__9592\,
            I => \N__9581\
        );

    \I__1577\ : InMux
    port map (
            O => \N__9591\,
            I => \N__9578\
        );

    \I__1576\ : InMux
    port map (
            O => \N__9590\,
            I => \N__9571\
        );

    \I__1575\ : InMux
    port map (
            O => \N__9589\,
            I => \N__9571\
        );

    \I__1574\ : InMux
    port map (
            O => \N__9588\,
            I => \N__9571\
        );

    \I__1573\ : InMux
    port map (
            O => \N__9587\,
            I => \N__9568\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__9584\,
            I => \N__9565\
        );

    \I__1571\ : InMux
    port map (
            O => \N__9581\,
            I => \N__9562\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__9578\,
            I => \uart_inst0.tx_uart_fifo_inst.wRamRdEn_1\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__9571\,
            I => \uart_inst0.tx_uart_fifo_inst.wRamRdEn_1\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__9568\,
            I => \uart_inst0.tx_uart_fifo_inst.wRamRdEn_1\
        );

    \I__1567\ : Odrv4
    port map (
            O => \N__9565\,
            I => \uart_inst0.tx_uart_fifo_inst.wRamRdEn_1\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__9562\,
            I => \uart_inst0.tx_uart_fifo_inst.wRamRdEn_1\
        );

    \I__1565\ : CascadeMux
    port map (
            O => \N__9551\,
            I => \N__9548\
        );

    \I__1564\ : InMux
    port map (
            O => \N__9548\,
            I => \N__9545\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__9545\,
            I => \N__9542\
        );

    \I__1562\ : Span4Mux_v
    port map (
            O => \N__9542\,
            I => \N__9539\
        );

    \I__1561\ : Odrv4
    port map (
            O => \N__9539\,
            I => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0\
        );

    \I__1560\ : InMux
    port map (
            O => \N__9536\,
            I => \N__9530\
        );

    \I__1559\ : InMux
    port map (
            O => \N__9535\,
            I => \N__9530\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__9530\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIBDOK2Z0Z_0\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__9527\,
            I => \N__9523\
        );

    \I__1556\ : InMux
    port map (
            O => \N__9526\,
            I => \N__9519\
        );

    \I__1555\ : InMux
    port map (
            O => \N__9523\,
            I => \N__9514\
        );

    \I__1554\ : InMux
    port map (
            O => \N__9522\,
            I => \N__9514\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__9519\,
            I => \uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__9514\,
            I => \uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7\
        );

    \I__1551\ : InMux
    port map (
            O => \N__9509\,
            I => \N__9501\
        );

    \I__1550\ : InMux
    port map (
            O => \N__9508\,
            I => \N__9501\
        );

    \I__1549\ : InMux
    port map (
            O => \N__9507\,
            I => \N__9496\
        );

    \I__1548\ : CascadeMux
    port map (
            O => \N__9506\,
            I => \N__9493\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__9501\,
            I => \N__9490\
        );

    \I__1546\ : InMux
    port map (
            O => \N__9500\,
            I => \N__9484\
        );

    \I__1545\ : InMux
    port map (
            O => \N__9499\,
            I => \N__9481\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__9496\,
            I => \N__9478\
        );

    \I__1543\ : InMux
    port map (
            O => \N__9493\,
            I => \N__9475\
        );

    \I__1542\ : Span4Mux_v
    port map (
            O => \N__9490\,
            I => \N__9472\
        );

    \I__1541\ : InMux
    port map (
            O => \N__9489\,
            I => \N__9465\
        );

    \I__1540\ : InMux
    port map (
            O => \N__9488\,
            I => \N__9465\
        );

    \I__1539\ : InMux
    port map (
            O => \N__9487\,
            I => \N__9465\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__9484\,
            I => \uart_inst0.wTxRdEn_0\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__9481\,
            I => \uart_inst0.wTxRdEn_0\
        );

    \I__1536\ : Odrv4
    port map (
            O => \N__9478\,
            I => \uart_inst0.wTxRdEn_0\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__9475\,
            I => \uart_inst0.wTxRdEn_0\
        );

    \I__1534\ : Odrv4
    port map (
            O => \N__9472\,
            I => \uart_inst0.wTxRdEn_0\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__9465\,
            I => \uart_inst0.wTxRdEn_0\
        );

    \I__1532\ : CascadeMux
    port map (
            O => \N__9452\,
            I => \N__9449\
        );

    \I__1531\ : InMux
    port map (
            O => \N__9449\,
            I => \N__9446\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__9446\,
            I => \N__9443\
        );

    \I__1529\ : Odrv12
    port map (
            O => \N__9443\,
            I => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_5\
        );

    \I__1528\ : CascadeMux
    port map (
            O => \N__9440\,
            I => \N__9437\
        );

    \I__1527\ : InMux
    port map (
            O => \N__9437\,
            I => \N__9434\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__9434\,
            I => \N__9431\
        );

    \I__1525\ : Odrv12
    port map (
            O => \N__9431\,
            I => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_6\
        );

    \I__1524\ : CascadeMux
    port map (
            O => \N__9428\,
            I => \N__9425\
        );

    \I__1523\ : InMux
    port map (
            O => \N__9425\,
            I => \N__9422\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__9422\,
            I => \N__9419\
        );

    \I__1521\ : Odrv12
    port map (
            O => \N__9419\,
            I => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_7\
        );

    \I__1520\ : InMux
    port map (
            O => \N__9416\,
            I => \N__9412\
        );

    \I__1519\ : InMux
    port map (
            O => \N__9415\,
            I => \N__9409\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__9412\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_0\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__9409\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_0\
        );

    \I__1516\ : InMux
    port map (
            O => \N__9404\,
            I => \N__9400\
        );

    \I__1515\ : InMux
    port map (
            O => \N__9403\,
            I => \N__9397\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__9400\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_3\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__9397\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_3\
        );

    \I__1512\ : InMux
    port map (
            O => \N__9392\,
            I => \N__9389\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__9389\,
            I => \uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_4\
        );

    \I__1510\ : InMux
    port map (
            O => \N__9386\,
            I => \N__9383\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__9383\,
            I => \rUartRxDataZ0Z_5\
        );

    \I__1508\ : InMux
    port map (
            O => \N__9380\,
            I => \N__9377\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__9377\,
            I => \rUartRxDataZ0Z_6\
        );

    \I__1506\ : InMux
    port map (
            O => \N__9374\,
            I => \N__9371\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__9371\,
            I => \N__9368\
        );

    \I__1504\ : Odrv4
    port map (
            O => \N__9368\,
            I => \rUartRxDataZ0Z_1\
        );

    \I__1503\ : CascadeMux
    port map (
            O => \N__9365\,
            I => \N__9362\
        );

    \I__1502\ : InMux
    port map (
            O => \N__9362\,
            I => \N__9359\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__9359\,
            I => \N__9356\
        );

    \I__1500\ : Span4Mux_h
    port map (
            O => \N__9356\,
            I => \N__9353\
        );

    \I__1499\ : Odrv4
    port map (
            O => \N__9353\,
            I => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_2\
        );

    \I__1498\ : CascadeMux
    port map (
            O => \N__9350\,
            I => \N__9346\
        );

    \I__1497\ : InMux
    port map (
            O => \N__9349\,
            I => \N__9341\
        );

    \I__1496\ : InMux
    port map (
            O => \N__9346\,
            I => \N__9341\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__9341\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNISGZ0Z74\
        );

    \I__1494\ : InMux
    port map (
            O => \N__9338\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_6\
        );

    \I__1493\ : InMux
    port map (
            O => \N__9335\,
            I => \bfn_15_6_0_\
        );

    \I__1492\ : CascadeMux
    port map (
            O => \N__9332\,
            I => \N__9329\
        );

    \I__1491\ : InMux
    port map (
            O => \N__9329\,
            I => \N__9326\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__9326\,
            I => \N__9323\
        );

    \I__1489\ : Span4Mux_h
    port map (
            O => \N__9323\,
            I => \N__9319\
        );

    \I__1488\ : InMux
    port map (
            O => \N__9322\,
            I => \N__9316\
        );

    \I__1487\ : Odrv4
    port map (
            O => \N__9319\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIIT3CZ0\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__9316\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIIT3CZ0\
        );

    \I__1485\ : InMux
    port map (
            O => \N__9311\,
            I => \N__9307\
        );

    \I__1484\ : InMux
    port map (
            O => \N__9310\,
            I => \N__9304\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__9307\,
            I => \N__9299\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__9304\,
            I => \N__9296\
        );

    \I__1481\ : InMux
    port map (
            O => \N__9303\,
            I => \N__9292\
        );

    \I__1480\ : InMux
    port map (
            O => \N__9302\,
            I => \N__9289\
        );

    \I__1479\ : Span4Mux_v
    port map (
            O => \N__9299\,
            I => \N__9283\
        );

    \I__1478\ : Span4Mux_v
    port map (
            O => \N__9296\,
            I => \N__9283\
        );

    \I__1477\ : InMux
    port map (
            O => \N__9295\,
            I => \N__9280\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__9292\,
            I => \N__9275\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__9289\,
            I => \N__9275\
        );

    \I__1474\ : InMux
    port map (
            O => \N__9288\,
            I => \N__9272\
        );

    \I__1473\ : Odrv4
    port map (
            O => \N__9283\,
            I => \rTxEnZ0\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__9280\,
            I => \rTxEnZ0\
        );

    \I__1471\ : Odrv4
    port map (
            O => \N__9275\,
            I => \rTxEnZ0\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__9272\,
            I => \rTxEnZ0\
        );

    \I__1469\ : CascadeMux
    port map (
            O => \N__9263\,
            I => \N__9260\
        );

    \I__1468\ : InMux
    port map (
            O => \N__9260\,
            I => \N__9254\
        );

    \I__1467\ : CascadeMux
    port map (
            O => \N__9259\,
            I => \N__9248\
        );

    \I__1466\ : InMux
    port map (
            O => \N__9258\,
            I => \N__9243\
        );

    \I__1465\ : InMux
    port map (
            O => \N__9257\,
            I => \N__9243\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__9254\,
            I => \N__9240\
        );

    \I__1463\ : InMux
    port map (
            O => \N__9253\,
            I => \N__9232\
        );

    \I__1462\ : InMux
    port map (
            O => \N__9252\,
            I => \N__9232\
        );

    \I__1461\ : InMux
    port map (
            O => \N__9251\,
            I => \N__9227\
        );

    \I__1460\ : InMux
    port map (
            O => \N__9248\,
            I => \N__9227\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__9243\,
            I => \N__9222\
        );

    \I__1458\ : Span4Mux_v
    port map (
            O => \N__9240\,
            I => \N__9222\
        );

    \I__1457\ : InMux
    port map (
            O => \N__9239\,
            I => \N__9219\
        );

    \I__1456\ : InMux
    port map (
            O => \N__9238\,
            I => \N__9214\
        );

    \I__1455\ : InMux
    port map (
            O => \N__9237\,
            I => \N__9214\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__9232\,
            I => \fifo_inst_wTxRdEn\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__9227\,
            I => \fifo_inst_wTxRdEn\
        );

    \I__1452\ : Odrv4
    port map (
            O => \N__9222\,
            I => \fifo_inst_wTxRdEn\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__9219\,
            I => \fifo_inst_wTxRdEn\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__9214\,
            I => \fifo_inst_wTxRdEn\
        );

    \I__1449\ : InMux
    port map (
            O => \N__9203\,
            I => \N__9197\
        );

    \I__1448\ : InMux
    port map (
            O => \N__9202\,
            I => \N__9197\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__9197\,
            I => \N__9194\
        );

    \I__1446\ : Span4Mux_v
    port map (
            O => \N__9194\,
            I => \N__9191\
        );

    \I__1445\ : Odrv4
    port map (
            O => \N__9191\,
            I => \fifo_inst_tx_fifo_inst_rDataCount_0_sqmuxa\
        );

    \I__1444\ : CascadeMux
    port map (
            O => \N__9188\,
            I => \N__9184\
        );

    \I__1443\ : InMux
    port map (
            O => \N__9187\,
            I => \N__9180\
        );

    \I__1442\ : InMux
    port map (
            O => \N__9184\,
            I => \N__9174\
        );

    \I__1441\ : InMux
    port map (
            O => \N__9183\,
            I => \N__9174\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__9180\,
            I => \N__9171\
        );

    \I__1439\ : InMux
    port map (
            O => \N__9179\,
            I => \N__9168\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__9174\,
            I => \fifo_inst_ft2232h_inst_rWrDelay\
        );

    \I__1437\ : Odrv4
    port map (
            O => \N__9171\,
            I => \fifo_inst_ft2232h_inst_rWrDelay\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__9168\,
            I => \fifo_inst_ft2232h_inst_rWrDelay\
        );

    \I__1435\ : InMux
    port map (
            O => \N__9161\,
            I => \N__9156\
        );

    \I__1434\ : InMux
    port map (
            O => \N__9160\,
            I => \N__9150\
        );

    \I__1433\ : InMux
    port map (
            O => \N__9159\,
            I => \N__9150\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__9156\,
            I => \N__9147\
        );

    \I__1431\ : InMux
    port map (
            O => \N__9155\,
            I => \N__9144\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__9150\,
            I => \fifo_inst_ft2232h_inst_rFifoState_4\
        );

    \I__1429\ : Odrv4
    port map (
            O => \N__9147\,
            I => \fifo_inst_ft2232h_inst_rFifoState_4\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__9144\,
            I => \fifo_inst_ft2232h_inst_rFifoState_4\
        );

    \I__1427\ : CascadeMux
    port map (
            O => \N__9137\,
            I => \N__9134\
        );

    \I__1426\ : InMux
    port map (
            O => \N__9134\,
            I => \N__9131\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__9131\,
            I => \N__9128\
        );

    \I__1424\ : Span4Mux_h
    port map (
            O => \N__9128\,
            I => \N__9124\
        );

    \I__1423\ : InMux
    port map (
            O => \N__9127\,
            I => \N__9121\
        );

    \I__1422\ : Odrv4
    port map (
            O => \N__9124\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNIO67CZ0\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__9121\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNIO67CZ0\
        );

    \I__1420\ : InMux
    port map (
            O => \N__9116\,
            I => \N__9113\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__9113\,
            I => \N__9110\
        );

    \I__1418\ : Span4Mux_v
    port map (
            O => \N__9110\,
            I => \N__9107\
        );

    \I__1417\ : Odrv4
    port map (
            O => \N__9107\,
            I => \rUartTxDataZ0Z_6\
        );

    \I__1416\ : InMux
    port map (
            O => \N__9104\,
            I => \N__9101\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__9101\,
            I => \N__9098\
        );

    \I__1414\ : Span4Mux_v
    port map (
            O => \N__9098\,
            I => \N__9095\
        );

    \I__1413\ : Odrv4
    port map (
            O => \N__9095\,
            I => \rUartTxDataZ0Z_5\
        );

    \I__1412\ : InMux
    port map (
            O => \N__9092\,
            I => \N__9089\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__9089\,
            I => \N__9086\
        );

    \I__1410\ : Span4Mux_v
    port map (
            O => \N__9086\,
            I => \N__9083\
        );

    \I__1409\ : Span4Mux_h
    port map (
            O => \N__9083\,
            I => \N__9080\
        );

    \I__1408\ : Odrv4
    port map (
            O => \N__9080\,
            I => \rUartTxDataZ0Z_1\
        );

    \I__1407\ : InMux
    port map (
            O => \N__9077\,
            I => \N__9066\
        );

    \I__1406\ : InMux
    port map (
            O => \N__9076\,
            I => \N__9066\
        );

    \I__1405\ : InMux
    port map (
            O => \N__9075\,
            I => \N__9061\
        );

    \I__1404\ : InMux
    port map (
            O => \N__9074\,
            I => \N__9061\
        );

    \I__1403\ : InMux
    port map (
            O => \N__9073\,
            I => \N__9056\
        );

    \I__1402\ : InMux
    port map (
            O => \N__9072\,
            I => \N__9056\
        );

    \I__1401\ : InMux
    port map (
            O => \N__9071\,
            I => \N__9053\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__9066\,
            I => \fifo_inst_wRxWrEn\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__9061\,
            I => \fifo_inst_wRxWrEn\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__9056\,
            I => \fifo_inst_wRxWrEn\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__9053\,
            I => \fifo_inst_wRxWrEn\
        );

    \I__1396\ : InMux
    port map (
            O => \N__9044\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_0\
        );

    \I__1395\ : CascadeMux
    port map (
            O => \N__9041\,
            I => \N__9038\
        );

    \I__1394\ : InMux
    port map (
            O => \N__9038\,
            I => \N__9035\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__9035\,
            I => \N__9032\
        );

    \I__1392\ : Span4Mux_v
    port map (
            O => \N__9032\,
            I => \N__9028\
        );

    \I__1391\ : InMux
    port map (
            O => \N__9031\,
            I => \N__9025\
        );

    \I__1390\ : Odrv4
    port map (
            O => \N__9028\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNICK0CZ0\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__9025\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNICK0CZ0\
        );

    \I__1388\ : InMux
    port map (
            O => \N__9020\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_1\
        );

    \I__1387\ : InMux
    port map (
            O => \N__9017\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_2\
        );

    \I__1386\ : InMux
    port map (
            O => \N__9014\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_3\
        );

    \I__1385\ : InMux
    port map (
            O => \N__9011\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_4\
        );

    \I__1384\ : CascadeMux
    port map (
            O => \N__9008\,
            I => \N__9005\
        );

    \I__1383\ : InMux
    port map (
            O => \N__9005\,
            I => \N__9002\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__9002\,
            I => \N__8999\
        );

    \I__1381\ : Span4Mux_s2_v
    port map (
            O => \N__8999\,
            I => \N__8996\
        );

    \I__1380\ : Span4Mux_h
    port map (
            O => \N__8996\,
            I => \N__8992\
        );

    \I__1379\ : InMux
    port map (
            O => \N__8995\,
            I => \N__8989\
        );

    \I__1378\ : Odrv4
    port map (
            O => \N__8992\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIK05CZ0\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__8989\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIK05CZ0\
        );

    \I__1376\ : InMux
    port map (
            O => \N__8984\,
            I => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_5\
        );

    \I__1375\ : InMux
    port map (
            O => \N__8981\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_2\
        );

    \I__1374\ : InMux
    port map (
            O => \N__8978\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_3\
        );

    \I__1373\ : CascadeMux
    port map (
            O => \N__8975\,
            I => \N__8972\
        );

    \I__1372\ : InMux
    port map (
            O => \N__8972\,
            I => \N__8969\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__8969\,
            I => \N__8966\
        );

    \I__1370\ : Span4Mux_s2_v
    port map (
            O => \N__8966\,
            I => \N__8962\
        );

    \I__1369\ : InMux
    port map (
            O => \N__8965\,
            I => \N__8959\
        );

    \I__1368\ : Odrv4
    port map (
            O => \N__8962\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIMJ1QZ0\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__8959\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIMJ1QZ0\
        );

    \I__1366\ : InMux
    port map (
            O => \N__8954\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_4\
        );

    \I__1365\ : CascadeMux
    port map (
            O => \N__8951\,
            I => \N__8948\
        );

    \I__1364\ : InMux
    port map (
            O => \N__8948\,
            I => \N__8945\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__8945\,
            I => \N__8942\
        );

    \I__1362\ : Span4Mux_h
    port map (
            O => \N__8942\,
            I => \N__8938\
        );

    \I__1361\ : InMux
    port map (
            O => \N__8941\,
            I => \N__8935\
        );

    \I__1360\ : Odrv4
    port map (
            O => \N__8938\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIOM2QZ0\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__8935\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIOM2QZ0\
        );

    \I__1358\ : InMux
    port map (
            O => \N__8930\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_5\
        );

    \I__1357\ : CascadeMux
    port map (
            O => \N__8927\,
            I => \N__8924\
        );

    \I__1356\ : InMux
    port map (
            O => \N__8924\,
            I => \N__8921\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__8921\,
            I => \N__8918\
        );

    \I__1354\ : Span4Mux_h
    port map (
            O => \N__8918\,
            I => \N__8914\
        );

    \I__1353\ : InMux
    port map (
            O => \N__8917\,
            I => \N__8911\
        );

    \I__1352\ : Odrv4
    port map (
            O => \N__8914\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIQP3QZ0\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__8911\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIQP3QZ0\
        );

    \I__1350\ : InMux
    port map (
            O => \N__8906\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_6\
        );

    \I__1349\ : InMux
    port map (
            O => \N__8903\,
            I => \bfn_15_4_0_\
        );

    \I__1348\ : CascadeMux
    port map (
            O => \N__8900\,
            I => \N__8897\
        );

    \I__1347\ : InMux
    port map (
            O => \N__8897\,
            I => \N__8894\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__8894\,
            I => \N__8891\
        );

    \I__1345\ : Span4Mux_h
    port map (
            O => \N__8891\,
            I => \N__8887\
        );

    \I__1344\ : InMux
    port map (
            O => \N__8890\,
            I => \N__8884\
        );

    \I__1343\ : Odrv4
    port map (
            O => \N__8887\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIE7TPZ0\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__8884\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIE7TPZ0\
        );

    \I__1341\ : CascadeMux
    port map (
            O => \N__8879\,
            I => \N__8876\
        );

    \I__1340\ : InMux
    port map (
            O => \N__8876\,
            I => \N__8873\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__8873\,
            I => \N__8870\
        );

    \I__1338\ : Span4Mux_h
    port map (
            O => \N__8870\,
            I => \N__8866\
        );

    \I__1337\ : InMux
    port map (
            O => \N__8869\,
            I => \N__8863\
        );

    \I__1336\ : Odrv4
    port map (
            O => \N__8866\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNISS4QZ0\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__8863\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNISS4QZ0\
        );

    \I__1334\ : InMux
    port map (
            O => \N__8858\,
            I => \N__8855\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__8855\,
            I => \N__8852\
        );

    \I__1332\ : Span4Mux_s1_v
    port map (
            O => \N__8852\,
            I => \N__8849\
        );

    \I__1331\ : Odrv4
    port map (
            O => \N__8849\,
            I => \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_0\
        );

    \I__1330\ : IoInMux
    port map (
            O => \N__8846\,
            I => \N__8843\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__8843\,
            I => \N__8840\
        );

    \I__1328\ : Span4Mux_s0_v
    port map (
            O => \N__8840\,
            I => \N__8837\
        );

    \I__1327\ : Odrv4
    port map (
            O => \N__8837\,
            I => \wTxRdData_0\
        );

    \I__1326\ : InMux
    port map (
            O => \N__8834\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_0\
        );

    \I__1325\ : InMux
    port map (
            O => \N__8831\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_1\
        );

    \I__1324\ : InMux
    port map (
            O => \N__8828\,
            I => \N__8825\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__8825\,
            I => \uart_inst0.uart_inst0.N_141_0\
        );

    \I__1322\ : InMux
    port map (
            O => \N__8822\,
            I => \N__8819\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__8819\,
            I => \uart_inst0.uart_inst0.N_143_0\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__8816\,
            I => \uart_inst0.uart_inst0.N_143_0_cascade_\
        );

    \I__1319\ : CEMux
    port map (
            O => \N__8813\,
            I => \N__8810\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__8810\,
            I => \N__8807\
        );

    \I__1317\ : Span4Mux_v
    port map (
            O => \N__8807\,
            I => \N__8803\
        );

    \I__1316\ : CEMux
    port map (
            O => \N__8806\,
            I => \N__8800\
        );

    \I__1315\ : Odrv4
    port map (
            O => \N__8803\,
            I => \uart_inst0.uart_inst0.N_143_0_0\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__8800\,
            I => \uart_inst0.uart_inst0.N_143_0_0\
        );

    \I__1313\ : CascadeMux
    port map (
            O => \N__8795\,
            I => \N__8792\
        );

    \I__1312\ : InMux
    port map (
            O => \N__8792\,
            I => \N__8789\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__8789\,
            I => \uart_inst0.uart_inst0.un1_m3_0_a2_2_1\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__8786\,
            I => \uart_inst0.uart_inst0.N_136_0_cascade_\
        );

    \I__1309\ : InMux
    port map (
            O => \N__8783\,
            I => \N__8780\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__8780\,
            I => \uart_inst0.uart_inst0.un1_tx_bits_remaining_c1\
        );

    \I__1307\ : InMux
    port map (
            O => \N__8777\,
            I => \N__8772\
        );

    \I__1306\ : InMux
    port map (
            O => \N__8776\,
            I => \N__8767\
        );

    \I__1305\ : InMux
    port map (
            O => \N__8775\,
            I => \N__8767\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__8772\,
            I => \uart_inst0.uart_inst0.N_136_0\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__8767\,
            I => \uart_inst0.uart_inst0.N_136_0\
        );

    \I__1302\ : InMux
    port map (
            O => \N__8762\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_3\
        );

    \I__1301\ : InMux
    port map (
            O => \N__8759\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_4\
        );

    \I__1300\ : InMux
    port map (
            O => \N__8756\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_5\
        );

    \I__1299\ : InMux
    port map (
            O => \N__8753\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_6\
        );

    \I__1298\ : InMux
    port map (
            O => \N__8750\,
            I => \bfn_14_12_0_\
        );

    \I__1297\ : CascadeMux
    port map (
            O => \N__8747\,
            I => \N__8744\
        );

    \I__1296\ : InMux
    port map (
            O => \N__8744\,
            I => \N__8739\
        );

    \I__1295\ : InMux
    port map (
            O => \N__8743\,
            I => \N__8736\
        );

    \I__1294\ : InMux
    port map (
            O => \N__8742\,
            I => \N__8733\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__8739\,
            I => \N__8730\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__8736\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_7\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__8733\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_7\
        );

    \I__1290\ : Odrv12
    port map (
            O => \N__8730\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_7\
        );

    \I__1289\ : CascadeMux
    port map (
            O => \N__8723\,
            I => \N__8720\
        );

    \I__1288\ : InMux
    port map (
            O => \N__8720\,
            I => \N__8717\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__8717\,
            I => \N__8714\
        );

    \I__1286\ : Span4Mux_h
    port map (
            O => \N__8714\,
            I => \N__8709\
        );

    \I__1285\ : InMux
    port map (
            O => \N__8713\,
            I => \N__8706\
        );

    \I__1284\ : InMux
    port map (
            O => \N__8712\,
            I => \N__8703\
        );

    \I__1283\ : Odrv4
    port map (
            O => \N__8709\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_5\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__8706\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_5\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__8703\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_5\
        );

    \I__1280\ : CascadeMux
    port map (
            O => \N__8696\,
            I => \N__8693\
        );

    \I__1279\ : InMux
    port map (
            O => \N__8693\,
            I => \N__8689\
        );

    \I__1278\ : CascadeMux
    port map (
            O => \N__8692\,
            I => \N__8686\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__8689\,
            I => \N__8682\
        );

    \I__1276\ : InMux
    port map (
            O => \N__8686\,
            I => \N__8679\
        );

    \I__1275\ : InMux
    port map (
            O => \N__8685\,
            I => \N__8676\
        );

    \I__1274\ : Odrv12
    port map (
            O => \N__8682\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_6\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__8679\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_6\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__8676\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_6\
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__8669\,
            I => \N__8666\
        );

    \I__1270\ : InMux
    port map (
            O => \N__8666\,
            I => \N__8663\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__8663\,
            I => \N__8658\
        );

    \I__1268\ : InMux
    port map (
            O => \N__8662\,
            I => \N__8655\
        );

    \I__1267\ : InMux
    port map (
            O => \N__8661\,
            I => \N__8652\
        );

    \I__1266\ : Odrv12
    port map (
            O => \N__8658\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_4\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__8655\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_4\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__8652\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_4\
        );

    \I__1263\ : CascadeMux
    port map (
            O => \N__8645\,
            I => \N__8641\
        );

    \I__1262\ : CascadeMux
    port map (
            O => \N__8644\,
            I => \N__8638\
        );

    \I__1261\ : InMux
    port map (
            O => \N__8641\,
            I => \N__8635\
        );

    \I__1260\ : InMux
    port map (
            O => \N__8638\,
            I => \N__8632\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__8635\,
            I => \N__8629\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__8632\,
            I => \N__8626\
        );

    \I__1257\ : Span4Mux_h
    port map (
            O => \N__8629\,
            I => \N__8623\
        );

    \I__1256\ : Span4Mux_h
    port map (
            O => \N__8626\,
            I => \N__8620\
        );

    \I__1255\ : Odrv4
    port map (
            O => \N__8623\,
            I => \uart_inst0.tx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_5\
        );

    \I__1254\ : Odrv4
    port map (
            O => \N__8620\,
            I => \uart_inst0.tx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_5\
        );

    \I__1253\ : IoInMux
    port map (
            O => \N__8615\,
            I => \N__8612\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__8612\,
            I => \N__8609\
        );

    \I__1251\ : IoSpan4Mux
    port map (
            O => \N__8609\,
            I => \N__8606\
        );

    \I__1250\ : Span4Mux_s0_v
    port map (
            O => \N__8606\,
            I => \N__8603\
        );

    \I__1249\ : Sp12to4
    port map (
            O => \N__8603\,
            I => \N__8599\
        );

    \I__1248\ : CascadeMux
    port map (
            O => \N__8602\,
            I => \N__8596\
        );

    \I__1247\ : Span12Mux_v
    port map (
            O => \N__8599\,
            I => \N__8593\
        );

    \I__1246\ : InMux
    port map (
            O => \N__8596\,
            I => \N__8590\
        );

    \I__1245\ : Odrv12
    port map (
            O => \N__8593\,
            I => \P1A7_c\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__8590\,
            I => \P1A7_c\
        );

    \I__1243\ : InMux
    port map (
            O => \N__8585\,
            I => \N__8576\
        );

    \I__1242\ : InMux
    port map (
            O => \N__8584\,
            I => \N__8563\
        );

    \I__1241\ : InMux
    port map (
            O => \N__8583\,
            I => \N__8563\
        );

    \I__1240\ : InMux
    port map (
            O => \N__8582\,
            I => \N__8563\
        );

    \I__1239\ : InMux
    port map (
            O => \N__8581\,
            I => \N__8563\
        );

    \I__1238\ : InMux
    port map (
            O => \N__8580\,
            I => \N__8563\
        );

    \I__1237\ : InMux
    port map (
            O => \N__8579\,
            I => \N__8559\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__8576\,
            I => \N__8556\
        );

    \I__1235\ : InMux
    port map (
            O => \N__8575\,
            I => \N__8551\
        );

    \I__1234\ : InMux
    port map (
            O => \N__8574\,
            I => \N__8551\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__8563\,
            I => \N__8548\
        );

    \I__1232\ : InMux
    port map (
            O => \N__8562\,
            I => \N__8545\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__8559\,
            I => \uart_inst0.uart_inst0.tx_state_81_d\
        );

    \I__1230\ : Odrv4
    port map (
            O => \N__8556\,
            I => \uart_inst0.uart_inst0.tx_state_81_d\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__8551\,
            I => \uart_inst0.uart_inst0.tx_state_81_d\
        );

    \I__1228\ : Odrv4
    port map (
            O => \N__8548\,
            I => \uart_inst0.uart_inst0.tx_state_81_d\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__8545\,
            I => \uart_inst0.uart_inst0.tx_state_81_d\
        );

    \I__1226\ : InMux
    port map (
            O => \N__8534\,
            I => \N__8531\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__8531\,
            I => \uart_inst0.uart_inst0.rTxDataZ0Z_0\
        );

    \I__1224\ : InMux
    port map (
            O => \N__8528\,
            I => \N__8525\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__8525\,
            I => \uart_inst0.uart_inst0.rTx_6_f1_0\
        );

    \I__1222\ : InMux
    port map (
            O => \N__8522\,
            I => \N__8519\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__8519\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c2\
        );

    \I__1220\ : CascadeMux
    port map (
            O => \N__8516\,
            I => \N__8511\
        );

    \I__1219\ : InMux
    port map (
            O => \N__8515\,
            I => \N__8506\
        );

    \I__1218\ : InMux
    port map (
            O => \N__8514\,
            I => \N__8502\
        );

    \I__1217\ : InMux
    port map (
            O => \N__8511\,
            I => \N__8499\
        );

    \I__1216\ : CEMux
    port map (
            O => \N__8510\,
            I => \N__8496\
        );

    \I__1215\ : CascadeMux
    port map (
            O => \N__8509\,
            I => \N__8493\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__8506\,
            I => \N__8488\
        );

    \I__1213\ : InMux
    port map (
            O => \N__8505\,
            I => \N__8485\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__8502\,
            I => \N__8480\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__8499\,
            I => \N__8480\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__8496\,
            I => \N__8477\
        );

    \I__1209\ : InMux
    port map (
            O => \N__8493\,
            I => \N__8470\
        );

    \I__1208\ : InMux
    port map (
            O => \N__8492\,
            I => \N__8470\
        );

    \I__1207\ : InMux
    port map (
            O => \N__8491\,
            I => \N__8467\
        );

    \I__1206\ : Span4Mux_v
    port map (
            O => \N__8488\,
            I => \N__8462\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__8485\,
            I => \N__8462\
        );

    \I__1204\ : Span4Mux_h
    port map (
            O => \N__8480\,
            I => \N__8457\
        );

    \I__1203\ : Span4Mux_h
    port map (
            O => \N__8477\,
            I => \N__8457\
        );

    \I__1202\ : InMux
    port map (
            O => \N__8476\,
            I => \N__8454\
        );

    \I__1201\ : InMux
    port map (
            O => \N__8475\,
            I => \N__8451\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__8470\,
            I => \N__8448\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__8467\,
            I => \N__8445\
        );

    \I__1198\ : Span4Mux_v
    port map (
            O => \N__8462\,
            I => \N__8440\
        );

    \I__1197\ : Span4Mux_v
    port map (
            O => \N__8457\,
            I => \N__8440\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__8454\,
            I => \uart_inst0.tx_uart_fifo_inst.wRamWrEn_1\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__8451\,
            I => \uart_inst0.tx_uart_fifo_inst.wRamWrEn_1\
        );

    \I__1194\ : Odrv4
    port map (
            O => \N__8448\,
            I => \uart_inst0.tx_uart_fifo_inst.wRamWrEn_1\
        );

    \I__1193\ : Odrv12
    port map (
            O => \N__8445\,
            I => \uart_inst0.tx_uart_fifo_inst.wRamWrEn_1\
        );

    \I__1192\ : Odrv4
    port map (
            O => \N__8440\,
            I => \uart_inst0.tx_uart_fifo_inst.wRamWrEn_1\
        );

    \I__1191\ : CascadeMux
    port map (
            O => \N__8429\,
            I => \N__8426\
        );

    \I__1190\ : InMux
    port map (
            O => \N__8426\,
            I => \N__8423\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__8423\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rDataCount_axbxc1_0\
        );

    \I__1188\ : InMux
    port map (
            O => \N__8420\,
            I => \N__8414\
        );

    \I__1187\ : InMux
    port map (
            O => \N__8419\,
            I => \N__8414\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__8414\,
            I => \N__8411\
        );

    \I__1185\ : Span4Mux_v
    port map (
            O => \N__8411\,
            I => \N__8404\
        );

    \I__1184\ : InMux
    port map (
            O => \N__8410\,
            I => \N__8401\
        );

    \I__1183\ : InMux
    port map (
            O => \N__8409\,
            I => \N__8394\
        );

    \I__1182\ : InMux
    port map (
            O => \N__8408\,
            I => \N__8394\
        );

    \I__1181\ : InMux
    port map (
            O => \N__8407\,
            I => \N__8394\
        );

    \I__1180\ : Odrv4
    port map (
            O => \N__8404\,
            I => \uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_1\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__8401\,
            I => \uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_1\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__8394\,
            I => \uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_1\
        );

    \I__1177\ : InMux
    port map (
            O => \N__8387\,
            I => \N__8383\
        );

    \I__1176\ : CascadeMux
    port map (
            O => \N__8386\,
            I => \N__8378\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__8383\,
            I => \N__8375\
        );

    \I__1174\ : InMux
    port map (
            O => \N__8382\,
            I => \N__8370\
        );

    \I__1173\ : InMux
    port map (
            O => \N__8381\,
            I => \N__8370\
        );

    \I__1172\ : InMux
    port map (
            O => \N__8378\,
            I => \N__8367\
        );

    \I__1171\ : Odrv12
    port map (
            O => \N__8375\,
            I => \uart_inst0.tx_uart_fifo_inst.rDataCountZ0Z_2\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__8370\,
            I => \uart_inst0.tx_uart_fifo_inst.rDataCountZ0Z_2\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__8367\,
            I => \uart_inst0.tx_uart_fifo_inst.rDataCountZ0Z_2\
        );

    \I__1168\ : CascadeMux
    port map (
            O => \N__8360\,
            I => \N__8357\
        );

    \I__1167\ : InMux
    port map (
            O => \N__8357\,
            I => \N__8352\
        );

    \I__1166\ : InMux
    port map (
            O => \N__8356\,
            I => \N__8346\
        );

    \I__1165\ : InMux
    port map (
            O => \N__8355\,
            I => \N__8343\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__8352\,
            I => \N__8340\
        );

    \I__1163\ : InMux
    port map (
            O => \N__8351\,
            I => \N__8337\
        );

    \I__1162\ : InMux
    port map (
            O => \N__8350\,
            I => \N__8332\
        );

    \I__1161\ : InMux
    port map (
            O => \N__8349\,
            I => \N__8332\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__8346\,
            I => \uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_0\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__8343\,
            I => \uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_0\
        );

    \I__1158\ : Odrv12
    port map (
            O => \N__8340\,
            I => \uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_0\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__8337\,
            I => \uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_0\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__8332\,
            I => \uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_0\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__8321\,
            I => \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIJHQM1Z0Z_2_cascade_\
        );

    \I__1154\ : InMux
    port map (
            O => \N__8318\,
            I => \N__8311\
        );

    \I__1153\ : InMux
    port map (
            O => \N__8317\,
            I => \N__8308\
        );

    \I__1152\ : InMux
    port map (
            O => \N__8316\,
            I => \N__8305\
        );

    \I__1151\ : CascadeMux
    port map (
            O => \N__8315\,
            I => \N__8302\
        );

    \I__1150\ : InMux
    port map (
            O => \N__8314\,
            I => \N__8297\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__8311\,
            I => \N__8292\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__8308\,
            I => \N__8292\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__8305\,
            I => \N__8289\
        );

    \I__1146\ : InMux
    port map (
            O => \N__8302\,
            I => \N__8286\
        );

    \I__1145\ : InMux
    port map (
            O => \N__8301\,
            I => \N__8283\
        );

    \I__1144\ : InMux
    port map (
            O => \N__8300\,
            I => \N__8280\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__8297\,
            I => \uart_inst0.tx_uart_fifo_inst.wUartTxFull\
        );

    \I__1142\ : Odrv4
    port map (
            O => \N__8292\,
            I => \uart_inst0.tx_uart_fifo_inst.wUartTxFull\
        );

    \I__1141\ : Odrv12
    port map (
            O => \N__8289\,
            I => \uart_inst0.tx_uart_fifo_inst.wUartTxFull\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__8286\,
            I => \uart_inst0.tx_uart_fifo_inst.wUartTxFull\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__8283\,
            I => \uart_inst0.tx_uart_fifo_inst.wUartTxFull\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__8280\,
            I => \uart_inst0.tx_uart_fifo_inst.wUartTxFull\
        );

    \I__1137\ : InMux
    port map (
            O => \N__8267\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_0\
        );

    \I__1136\ : InMux
    port map (
            O => \N__8264\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_1\
        );

    \I__1135\ : InMux
    port map (
            O => \N__8261\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_2\
        );

    \I__1134\ : InMux
    port map (
            O => \N__8258\,
            I => \N__8253\
        );

    \I__1133\ : InMux
    port map (
            O => \N__8257\,
            I => \N__8248\
        );

    \I__1132\ : InMux
    port map (
            O => \N__8256\,
            I => \N__8248\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__8253\,
            I => \N__8245\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__8248\,
            I => \N__8240\
        );

    \I__1129\ : Span4Mux_s2_v
    port map (
            O => \N__8245\,
            I => \N__8240\
        );

    \I__1128\ : Odrv4
    port map (
            O => \N__8240\,
            I => \fifo_inst_ft2232h_inst_rFifoState_3\
        );

    \I__1127\ : InMux
    port map (
            O => \N__8237\,
            I => \N__8232\
        );

    \I__1126\ : InMux
    port map (
            O => \N__8236\,
            I => \N__8227\
        );

    \I__1125\ : InMux
    port map (
            O => \N__8235\,
            I => \N__8227\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__8232\,
            I => \fifo_inst_rx_fifo_inst_un1_rDataCount15_2_0_0\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__8227\,
            I => \fifo_inst_rx_fifo_inst_un1_rDataCount15_2_0_0\
        );

    \I__1122\ : InMux
    port map (
            O => \N__8222\,
            I => \N__8217\
        );

    \I__1121\ : InMux
    port map (
            O => \N__8221\,
            I => \N__8214\
        );

    \I__1120\ : InMux
    port map (
            O => \N__8220\,
            I => \N__8211\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__8217\,
            I => \fifo_inst_rx_fifo_inst_rDataCount_fast_0\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__8214\,
            I => \fifo_inst_rx_fifo_inst_rDataCount_fast_0\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__8211\,
            I => \fifo_inst_rx_fifo_inst_rDataCount_fast_0\
        );

    \I__1116\ : InMux
    port map (
            O => \N__8204\,
            I => \N__8201\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__8201\,
            I => \N__8196\
        );

    \I__1114\ : InMux
    port map (
            O => \N__8200\,
            I => \N__8193\
        );

    \I__1113\ : InMux
    port map (
            O => \N__8199\,
            I => \N__8190\
        );

    \I__1112\ : Odrv4
    port map (
            O => \N__8196\,
            I => \N_84_mux\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__8193\,
            I => \N_84_mux\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__8190\,
            I => \N_84_mux\
        );

    \I__1109\ : CascadeMux
    port map (
            O => \N__8183\,
            I => \rUartTxEn_4_cascade_\
        );

    \I__1108\ : CascadeMux
    port map (
            O => \N__8180\,
            I => \N__8176\
        );

    \I__1107\ : InMux
    port map (
            O => \N__8179\,
            I => \N__8172\
        );

    \I__1106\ : InMux
    port map (
            O => \N__8176\,
            I => \N__8167\
        );

    \I__1105\ : InMux
    port map (
            O => \N__8175\,
            I => \N__8167\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__8172\,
            I => \rFtdiRxStateZ0Z_0\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__8167\,
            I => \rFtdiRxStateZ0Z_0\
        );

    \I__1102\ : InMux
    port map (
            O => \N__8162\,
            I => \N__8159\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__8159\,
            I => \N__8156\
        );

    \I__1100\ : Span4Mux_s3_v
    port map (
            O => \N__8156\,
            I => \N__8153\
        );

    \I__1099\ : Odrv4
    port map (
            O => \N__8153\,
            I => \fifo_inst.ft2232h_inst.rFifoStatesr_0\
        );

    \I__1098\ : InMux
    port map (
            O => \N__8150\,
            I => \N__8147\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__8147\,
            I => \N__8143\
        );

    \I__1096\ : InMux
    port map (
            O => \N__8146\,
            I => \N__8140\
        );

    \I__1095\ : Span4Mux_h
    port map (
            O => \N__8143\,
            I => \N__8137\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__8140\,
            I => \N__8134\
        );

    \I__1093\ : Span4Mux_v
    port map (
            O => \N__8137\,
            I => \N__8130\
        );

    \I__1092\ : Span4Mux_h
    port map (
            O => \N__8134\,
            I => \N__8127\
        );

    \I__1091\ : InMux
    port map (
            O => \N__8133\,
            I => \N__8124\
        );

    \I__1090\ : Odrv4
    port map (
            O => \N__8130\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_2\
        );

    \I__1089\ : Odrv4
    port map (
            O => \N__8127\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_2\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__8124\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_2\
        );

    \I__1087\ : InMux
    port map (
            O => \N__8117\,
            I => \N__8113\
        );

    \I__1086\ : InMux
    port map (
            O => \N__8116\,
            I => \N__8110\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__8113\,
            I => \N__8107\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__8110\,
            I => \N__8104\
        );

    \I__1083\ : Span4Mux_v
    port map (
            O => \N__8107\,
            I => \N__8098\
        );

    \I__1082\ : Span4Mux_h
    port map (
            O => \N__8104\,
            I => \N__8098\
        );

    \I__1081\ : InMux
    port map (
            O => \N__8103\,
            I => \N__8095\
        );

    \I__1080\ : Span4Mux_v
    port map (
            O => \N__8098\,
            I => \N__8090\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__8095\,
            I => \N__8090\
        );

    \I__1078\ : Span4Mux_h
    port map (
            O => \N__8090\,
            I => \N__8087\
        );

    \I__1077\ : Sp12to4
    port map (
            O => \N__8087\,
            I => \N__8084\
        );

    \I__1076\ : Span12Mux_v
    port map (
            O => \N__8084\,
            I => \N__8081\
        );

    \I__1075\ : Odrv12
    port map (
            O => \N__8081\,
            I => \iRxF_n_c\
        );

    \I__1074\ : InMux
    port map (
            O => \N__8078\,
            I => \N__8074\
        );

    \I__1073\ : InMux
    port map (
            O => \N__8077\,
            I => \N__8071\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__8074\,
            I => \N__8068\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__8071\,
            I => \N__8064\
        );

    \I__1070\ : Span4Mux_h
    port map (
            O => \N__8068\,
            I => \N__8061\
        );

    \I__1069\ : InMux
    port map (
            O => \N__8067\,
            I => \N__8058\
        );

    \I__1068\ : Odrv12
    port map (
            O => \N__8064\,
            I => \fifo_inst_ft2232h_inst_rFifoState_0\
        );

    \I__1067\ : Odrv4
    port map (
            O => \N__8061\,
            I => \fifo_inst_ft2232h_inst_rFifoState_0\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__8058\,
            I => \fifo_inst_ft2232h_inst_rFifoState_0\
        );

    \I__1065\ : CascadeMux
    port map (
            O => \N__8051\,
            I => \fifo_inst.rx_fifo_inst.un1_rDataCount_axbxc3_1_1_cascade_\
        );

    \I__1064\ : CascadeMux
    port map (
            O => \N__8048\,
            I => \uart_inst0.tx_uart_fifo_inst.m15_xZ0Z0_cascade_\
        );

    \I__1063\ : InMux
    port map (
            O => \N__8045\,
            I => \N__8042\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__8042\,
            I => \fifo_inst.rx_fifo_inst.un1_rDataCount_axbxc3_1_1\
        );

    \I__1061\ : CascadeMux
    port map (
            O => \N__8039\,
            I => \N__8036\
        );

    \I__1060\ : InMux
    port map (
            O => \N__8036\,
            I => \N__8031\
        );

    \I__1059\ : InMux
    port map (
            O => \N__8035\,
            I => \N__8026\
        );

    \I__1058\ : InMux
    port map (
            O => \N__8034\,
            I => \N__8026\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__8031\,
            I => \fifo_inst_rx_fifo_inst_rDataCount_fast_3\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__8026\,
            I => \fifo_inst_rx_fifo_inst_rDataCount_fast_3\
        );

    \I__1055\ : IoInMux
    port map (
            O => \N__8021\,
            I => \N__8018\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__8018\,
            I => \N__8015\
        );

    \I__1053\ : IoSpan4Mux
    port map (
            O => \N__8015\,
            I => \N__8011\
        );

    \I__1052\ : IoInMux
    port map (
            O => \N__8014\,
            I => \N__8008\
        );

    \I__1051\ : Span4Mux_s0_v
    port map (
            O => \N__8011\,
            I => \N__8005\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__8008\,
            I => \N__8002\
        );

    \I__1049\ : Sp12to4
    port map (
            O => \N__8005\,
            I => \N__7999\
        );

    \I__1048\ : IoSpan4Mux
    port map (
            O => \N__8002\,
            I => \N__7996\
        );

    \I__1047\ : Span12Mux_v
    port map (
            O => \N__7999\,
            I => \N__7993\
        );

    \I__1046\ : Span4Mux_s3_v
    port map (
            O => \N__7996\,
            I => \N__7990\
        );

    \I__1045\ : Span12Mux_v
    port map (
            O => \N__7993\,
            I => \N__7986\
        );

    \I__1044\ : Span4Mux_h
    port map (
            O => \N__7990\,
            I => \N__7983\
        );

    \I__1043\ : InMux
    port map (
            O => \N__7989\,
            I => \N__7980\
        );

    \I__1042\ : Odrv12
    port map (
            O => \N__7986\,
            I => \P1A4_c\
        );

    \I__1041\ : Odrv4
    port map (
            O => \N__7983\,
            I => \P1A4_c\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__7980\,
            I => \P1A4_c\
        );

    \I__1039\ : CascadeMux
    port map (
            O => \N__7973\,
            I => \uart_inst0.tx_uart_fifo_inst.m8_xZ0Z0_cascade_\
        );

    \I__1038\ : InMux
    port map (
            O => \N__7970\,
            I => \N__7967\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__7967\,
            I => \N__7963\
        );

    \I__1036\ : InMux
    port map (
            O => \N__7966\,
            I => \N__7960\
        );

    \I__1035\ : Odrv4
    port map (
            O => \N__7963\,
            I => \fifo_inst.tx_fifo_inst.un1_rDataCount_axbxc3_2_tz\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__7960\,
            I => \fifo_inst.tx_fifo_inst.un1_rDataCount_axbxc3_2_tz\
        );

    \I__1033\ : CascadeMux
    port map (
            O => \N__7955\,
            I => \N__7952\
        );

    \I__1032\ : InMux
    port map (
            O => \N__7952\,
            I => \N__7948\
        );

    \I__1031\ : CascadeMux
    port map (
            O => \N__7951\,
            I => \N__7945\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__7948\,
            I => \N__7942\
        );

    \I__1029\ : InMux
    port map (
            O => \N__7945\,
            I => \N__7939\
        );

    \I__1028\ : Odrv4
    port map (
            O => \N__7942\,
            I => \fifo_inst.tx_fifo_inst.un1_rDataCount_axbxc3_a0_2\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__7939\,
            I => \fifo_inst.tx_fifo_inst.un1_rDataCount_axbxc3_a0_2\
        );

    \I__1026\ : InMux
    port map (
            O => \N__7934\,
            I => \N__7931\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__7931\,
            I => \fifo_inst.tx_fifo_inst.un1_rDataCount_c2_0\
        );

    \I__1024\ : CEMux
    port map (
            O => \N__7928\,
            I => \N__7924\
        );

    \I__1023\ : InMux
    port map (
            O => \N__7927\,
            I => \N__7920\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__7924\,
            I => \N__7915\
        );

    \I__1021\ : CascadeMux
    port map (
            O => \N__7923\,
            I => \N__7912\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__7920\,
            I => \N__7909\
        );

    \I__1019\ : CascadeMux
    port map (
            O => \N__7919\,
            I => \N__7906\
        );

    \I__1018\ : InMux
    port map (
            O => \N__7918\,
            I => \N__7903\
        );

    \I__1017\ : Span4Mux_h
    port map (
            O => \N__7915\,
            I => \N__7900\
        );

    \I__1016\ : InMux
    port map (
            O => \N__7912\,
            I => \N__7897\
        );

    \I__1015\ : Span4Mux_v
    port map (
            O => \N__7909\,
            I => \N__7894\
        );

    \I__1014\ : InMux
    port map (
            O => \N__7906\,
            I => \N__7891\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__7903\,
            I => \N__7886\
        );

    \I__1012\ : Span4Mux_h
    port map (
            O => \N__7900\,
            I => \N__7886\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__7897\,
            I => \fifo_inst_tx_fifo_inst_wRamWrEn\
        );

    \I__1010\ : Odrv4
    port map (
            O => \N__7894\,
            I => \fifo_inst_tx_fifo_inst_wRamWrEn\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__7891\,
            I => \fifo_inst_tx_fifo_inst_wRamWrEn\
        );

    \I__1008\ : Odrv4
    port map (
            O => \N__7886\,
            I => \fifo_inst_tx_fifo_inst_wRamWrEn\
        );

    \I__1007\ : CascadeMux
    port map (
            O => \N__7877\,
            I => \N__7874\
        );

    \I__1006\ : InMux
    port map (
            O => \N__7874\,
            I => \N__7870\
        );

    \I__1005\ : InMux
    port map (
            O => \N__7873\,
            I => \N__7867\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__7870\,
            I => \N__7863\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__7867\,
            I => \N__7860\
        );

    \I__1002\ : InMux
    port map (
            O => \N__7866\,
            I => \N__7857\
        );

    \I__1001\ : Span4Mux_h
    port map (
            O => \N__7863\,
            I => \N__7854\
        );

    \I__1000\ : Odrv4
    port map (
            O => \N__7860\,
            I => \fifo_inst.tx_fifo_inst.un1_rDataCount_ac0_1_a0_0\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__7857\,
            I => \fifo_inst.tx_fifo_inst.un1_rDataCount_ac0_1_a0_0\
        );

    \I__998\ : Odrv4
    port map (
            O => \N__7854\,
            I => \fifo_inst.tx_fifo_inst.un1_rDataCount_ac0_1_a0_0\
        );

    \I__997\ : CascadeMux
    port map (
            O => \N__7847\,
            I => \fifo_inst.tx_fifo_inst.un1_rDataCount_c2_1_cascade_\
        );

    \I__996\ : InMux
    port map (
            O => \N__7844\,
            I => \N__7841\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__7841\,
            I => \fifo_inst.tx_fifo_inst.un1_rDataCount_ac0_2\
        );

    \I__994\ : InMux
    port map (
            O => \N__7838\,
            I => \N__7834\
        );

    \I__993\ : InMux
    port map (
            O => \N__7837\,
            I => \N__7831\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__7834\,
            I => \fifo_inst_tx_fifo_inst_un1_rDataCount15_2_0_0\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__7831\,
            I => \fifo_inst_tx_fifo_inst_un1_rDataCount15_2_0_0\
        );

    \I__990\ : InMux
    port map (
            O => \N__7826\,
            I => \N__7820\
        );

    \I__989\ : InMux
    port map (
            O => \N__7825\,
            I => \N__7820\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__7820\,
            I => \N__7816\
        );

    \I__987\ : CascadeMux
    port map (
            O => \N__7819\,
            I => \N__7810\
        );

    \I__986\ : Span4Mux_s3_v
    port map (
            O => \N__7816\,
            I => \N__7807\
        );

    \I__985\ : InMux
    port map (
            O => \N__7815\,
            I => \N__7804\
        );

    \I__984\ : InMux
    port map (
            O => \N__7814\,
            I => \N__7799\
        );

    \I__983\ : InMux
    port map (
            O => \N__7813\,
            I => \N__7799\
        );

    \I__982\ : InMux
    port map (
            O => \N__7810\,
            I => \N__7796\
        );

    \I__981\ : Odrv4
    port map (
            O => \N__7807\,
            I => \fifo_inst_tx_fifo_inst_rDataCount_2\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__7804\,
            I => \fifo_inst_tx_fifo_inst_rDataCount_2\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__7799\,
            I => \fifo_inst_tx_fifo_inst_rDataCount_2\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__7796\,
            I => \fifo_inst_tx_fifo_inst_rDataCount_2\
        );

    \I__977\ : InMux
    port map (
            O => \N__7787\,
            I => \N__7780\
        );

    \I__976\ : InMux
    port map (
            O => \N__7786\,
            I => \N__7780\
        );

    \I__975\ : CascadeMux
    port map (
            O => \N__7785\,
            I => \N__7777\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__7780\,
            I => \N__7774\
        );

    \I__973\ : InMux
    port map (
            O => \N__7777\,
            I => \N__7766\
        );

    \I__972\ : Span4Mux_h
    port map (
            O => \N__7774\,
            I => \N__7763\
        );

    \I__971\ : InMux
    port map (
            O => \N__7773\,
            I => \N__7758\
        );

    \I__970\ : InMux
    port map (
            O => \N__7772\,
            I => \N__7758\
        );

    \I__969\ : InMux
    port map (
            O => \N__7771\,
            I => \N__7753\
        );

    \I__968\ : InMux
    port map (
            O => \N__7770\,
            I => \N__7753\
        );

    \I__967\ : InMux
    port map (
            O => \N__7769\,
            I => \N__7750\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__7766\,
            I => \fifo_inst_tx_fifo_inst_rDataCount_1\
        );

    \I__965\ : Odrv4
    port map (
            O => \N__7763\,
            I => \fifo_inst_tx_fifo_inst_rDataCount_1\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__7758\,
            I => \fifo_inst_tx_fifo_inst_rDataCount_1\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__7753\,
            I => \fifo_inst_tx_fifo_inst_rDataCount_1\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__7750\,
            I => \fifo_inst_tx_fifo_inst_rDataCount_1\
        );

    \I__961\ : CascadeMux
    port map (
            O => \N__7739\,
            I => \N__7736\
        );

    \I__960\ : InMux
    port map (
            O => \N__7736\,
            I => \N__7731\
        );

    \I__959\ : InMux
    port map (
            O => \N__7735\,
            I => \N__7726\
        );

    \I__958\ : InMux
    port map (
            O => \N__7734\,
            I => \N__7726\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__7731\,
            I => \fifo_inst_tx_fifo_inst_rDataCount_fast_3\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__7726\,
            I => \fifo_inst_tx_fifo_inst_rDataCount_fast_3\
        );

    \I__955\ : InMux
    port map (
            O => \N__7721\,
            I => \N__7712\
        );

    \I__954\ : InMux
    port map (
            O => \N__7720\,
            I => \N__7712\
        );

    \I__953\ : InMux
    port map (
            O => \N__7719\,
            I => \N__7706\
        );

    \I__952\ : InMux
    port map (
            O => \N__7718\,
            I => \N__7701\
        );

    \I__951\ : InMux
    port map (
            O => \N__7717\,
            I => \N__7701\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__7712\,
            I => \N__7698\
        );

    \I__949\ : InMux
    port map (
            O => \N__7711\,
            I => \N__7695\
        );

    \I__948\ : InMux
    port map (
            O => \N__7710\,
            I => \N__7690\
        );

    \I__947\ : InMux
    port map (
            O => \N__7709\,
            I => \N__7690\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__7706\,
            I => \fifo_inst_tx_fifo_inst_rDataCount_0\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__7701\,
            I => \fifo_inst_tx_fifo_inst_rDataCount_0\
        );

    \I__944\ : Odrv4
    port map (
            O => \N__7698\,
            I => \fifo_inst_tx_fifo_inst_rDataCount_0\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__7695\,
            I => \fifo_inst_tx_fifo_inst_rDataCount_0\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__7690\,
            I => \fifo_inst_tx_fifo_inst_rDataCount_0\
        );

    \I__941\ : InMux
    port map (
            O => \N__7679\,
            I => \N__7676\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__7676\,
            I => \N__7673\
        );

    \I__939\ : Span4Mux_v
    port map (
            O => \N__7673\,
            I => \N__7670\
        );

    \I__938\ : Odrv4
    port map (
            O => \N__7670\,
            I => \uart_inst0.wTxRdData_4\
        );

    \I__937\ : InMux
    port map (
            O => \N__7667\,
            I => \N__7664\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__7664\,
            I => \uart_inst0.uart_inst0.rTxDataZ0Z_4\
        );

    \I__935\ : InMux
    port map (
            O => \N__7661\,
            I => \N__7658\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__7658\,
            I => \uart_inst0.uart_inst0.rTxDataZ0Z_3\
        );

    \I__933\ : InMux
    port map (
            O => \N__7655\,
            I => \N__7652\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__7652\,
            I => \N__7649\
        );

    \I__931\ : Odrv12
    port map (
            O => \N__7649\,
            I => \uart_inst0.wTxRdData_2\
        );

    \I__930\ : InMux
    port map (
            O => \N__7646\,
            I => \N__7643\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__7643\,
            I => \uart_inst0.uart_inst0.rTxDataZ0Z_2\
        );

    \I__928\ : InMux
    port map (
            O => \N__7640\,
            I => \N__7637\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__7637\,
            I => \uart_inst0.uart_inst0.rTxDataZ0Z_6\
        );

    \I__926\ : InMux
    port map (
            O => \N__7634\,
            I => \N__7631\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__7631\,
            I => \N__7628\
        );

    \I__924\ : Odrv12
    port map (
            O => \N__7628\,
            I => \uart_inst0.wTxRdData_5\
        );

    \I__923\ : InMux
    port map (
            O => \N__7625\,
            I => \N__7622\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__7622\,
            I => \uart_inst0.uart_inst0.rTxDataZ0Z_5\
        );

    \I__921\ : InMux
    port map (
            O => \N__7619\,
            I => \N__7616\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__7616\,
            I => \N__7613\
        );

    \I__919\ : Odrv12
    port map (
            O => \N__7613\,
            I => \uart_inst0.wTxRdData_7\
        );

    \I__918\ : CascadeMux
    port map (
            O => \N__7610\,
            I => \N__7607\
        );

    \I__917\ : InMux
    port map (
            O => \N__7607\,
            I => \N__7603\
        );

    \I__916\ : InMux
    port map (
            O => \N__7606\,
            I => \N__7600\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__7603\,
            I => \uart_inst0.uart_inst0.rTxDataZ0Z_7\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__7600\,
            I => \uart_inst0.uart_inst0.rTxDataZ0Z_7\
        );

    \I__913\ : CascadeMux
    port map (
            O => \N__7595\,
            I => \N_97_cascade_\
        );

    \I__912\ : InMux
    port map (
            O => \N__7592\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_3\
        );

    \I__911\ : InMux
    port map (
            O => \N__7589\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_4\
        );

    \I__910\ : InMux
    port map (
            O => \N__7586\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_5\
        );

    \I__909\ : InMux
    port map (
            O => \N__7583\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_6\
        );

    \I__908\ : InMux
    port map (
            O => \N__7580\,
            I => \bfn_13_13_0_\
        );

    \I__907\ : CascadeMux
    port map (
            O => \N__7577\,
            I => \N__7574\
        );

    \I__906\ : InMux
    port map (
            O => \N__7574\,
            I => \N__7571\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__7571\,
            I => \N__7568\
        );

    \I__904\ : Span4Mux_v
    port map (
            O => \N__7568\,
            I => \N__7564\
        );

    \I__903\ : InMux
    port map (
            O => \N__7567\,
            I => \N__7560\
        );

    \I__902\ : Span4Mux_h
    port map (
            O => \N__7564\,
            I => \N__7557\
        );

    \I__901\ : InMux
    port map (
            O => \N__7563\,
            I => \N__7554\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__7560\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_8\
        );

    \I__899\ : Odrv4
    port map (
            O => \N__7557\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_8\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__7554\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_8\
        );

    \I__897\ : InMux
    port map (
            O => \N__7547\,
            I => \N__7544\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__7544\,
            I => \N__7541\
        );

    \I__895\ : Odrv12
    port map (
            O => \N__7541\,
            I => \uart_inst0.wTxRdData_0\
        );

    \I__894\ : InMux
    port map (
            O => \N__7538\,
            I => \N__7535\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__7535\,
            I => \N__7532\
        );

    \I__892\ : Odrv12
    port map (
            O => \N__7532\,
            I => \uart_inst0.wTxRdData_1\
        );

    \I__891\ : InMux
    port map (
            O => \N__7529\,
            I => \N__7526\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__7526\,
            I => \uart_inst0.uart_inst0.rTxDataZ0Z_1\
        );

    \I__889\ : InMux
    port map (
            O => \N__7523\,
            I => \N__7520\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__7520\,
            I => \N__7517\
        );

    \I__887\ : Odrv12
    port map (
            O => \N__7517\,
            I => \uart_inst0.wTxRdData_6\
        );

    \I__886\ : InMux
    port map (
            O => \N__7514\,
            I => \N__7511\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__7511\,
            I => \N__7508\
        );

    \I__884\ : Odrv12
    port map (
            O => \N__7508\,
            I => \uart_inst0.wTxRdData_3\
        );

    \I__883\ : InMux
    port map (
            O => \N__7505\,
            I => \N__7502\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__7502\,
            I => \N__7499\
        );

    \I__881\ : Span4Mux_v
    port map (
            O => \N__7499\,
            I => \N__7496\
        );

    \I__880\ : Span4Mux_h
    port map (
            O => \N__7496\,
            I => \N__7493\
        );

    \I__879\ : Odrv4
    port map (
            O => \N__7493\,
            I => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_3\
        );

    \I__878\ : InMux
    port map (
            O => \N__7490\,
            I => \N__7487\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__7487\,
            I => \N__7484\
        );

    \I__876\ : Span4Mux_h
    port map (
            O => \N__7484\,
            I => \N__7481\
        );

    \I__875\ : Odrv4
    port map (
            O => \N__7481\,
            I => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_4\
        );

    \I__874\ : InMux
    port map (
            O => \N__7478\,
            I => \N__7475\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__7475\,
            I => \N__7472\
        );

    \I__872\ : Span4Mux_h
    port map (
            O => \N__7472\,
            I => \N__7469\
        );

    \I__871\ : Odrv4
    port map (
            O => \N__7469\,
            I => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_5\
        );

    \I__870\ : InMux
    port map (
            O => \N__7466\,
            I => \N__7463\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__7463\,
            I => \N__7460\
        );

    \I__868\ : Odrv12
    port map (
            O => \N__7460\,
            I => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_6\
        );

    \I__867\ : InMux
    port map (
            O => \N__7457\,
            I => \N__7454\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__7454\,
            I => \N__7451\
        );

    \I__865\ : Span4Mux_h
    port map (
            O => \N__7451\,
            I => \N__7448\
        );

    \I__864\ : Odrv4
    port map (
            O => \N__7448\,
            I => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_7\
        );

    \I__863\ : CascadeMux
    port map (
            O => \N__7445\,
            I => \N__7442\
        );

    \I__862\ : InMux
    port map (
            O => \N__7442\,
            I => \N__7439\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__7439\,
            I => \N__7436\
        );

    \I__860\ : Span4Mux_h
    port map (
            O => \N__7436\,
            I => \N__7432\
        );

    \I__859\ : InMux
    port map (
            O => \N__7435\,
            I => \N__7428\
        );

    \I__858\ : Span4Mux_h
    port map (
            O => \N__7432\,
            I => \N__7425\
        );

    \I__857\ : InMux
    port map (
            O => \N__7431\,
            I => \N__7422\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__7428\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ1Z_0\
        );

    \I__855\ : Odrv4
    port map (
            O => \N__7425\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ1Z_0\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__7422\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ1Z_0\
        );

    \I__853\ : InMux
    port map (
            O => \N__7415\,
            I => \N__7412\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__7412\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNO_0Z0Z_0\
        );

    \I__851\ : CascadeMux
    port map (
            O => \N__7409\,
            I => \N__7406\
        );

    \I__850\ : InMux
    port map (
            O => \N__7406\,
            I => \N__7402\
        );

    \I__849\ : InMux
    port map (
            O => \N__7405\,
            I => \N__7398\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__7402\,
            I => \N__7395\
        );

    \I__847\ : InMux
    port map (
            O => \N__7401\,
            I => \N__7392\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__7398\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ1Z_1\
        );

    \I__845\ : Odrv12
    port map (
            O => \N__7395\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ1Z_1\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__7392\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ1Z_1\
        );

    \I__843\ : InMux
    port map (
            O => \N__7385\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_0\
        );

    \I__842\ : CascadeMux
    port map (
            O => \N__7382\,
            I => \N__7379\
        );

    \I__841\ : InMux
    port map (
            O => \N__7379\,
            I => \N__7376\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__7376\,
            I => \N__7372\
        );

    \I__839\ : InMux
    port map (
            O => \N__7375\,
            I => \N__7368\
        );

    \I__838\ : Span4Mux_h
    port map (
            O => \N__7372\,
            I => \N__7365\
        );

    \I__837\ : InMux
    port map (
            O => \N__7371\,
            I => \N__7362\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__7368\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ0Z_2\
        );

    \I__835\ : Odrv4
    port map (
            O => \N__7365\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ0Z_2\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__7362\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ0Z_2\
        );

    \I__833\ : InMux
    port map (
            O => \N__7355\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_1\
        );

    \I__832\ : CascadeMux
    port map (
            O => \N__7352\,
            I => \N__7349\
        );

    \I__831\ : InMux
    port map (
            O => \N__7349\,
            I => \N__7346\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__7346\,
            I => \N__7343\
        );

    \I__829\ : Span4Mux_h
    port map (
            O => \N__7343\,
            I => \N__7340\
        );

    \I__828\ : Span4Mux_h
    port map (
            O => \N__7340\,
            I => \N__7335\
        );

    \I__827\ : InMux
    port map (
            O => \N__7339\,
            I => \N__7332\
        );

    \I__826\ : InMux
    port map (
            O => \N__7338\,
            I => \N__7329\
        );

    \I__825\ : Odrv4
    port map (
            O => \N__7335\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_3\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__7332\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_3\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__7329\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_3\
        );

    \I__822\ : InMux
    port map (
            O => \N__7322\,
            I => \N__7319\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__7319\,
            I => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNO_0Z0Z_3\
        );

    \I__820\ : InMux
    port map (
            O => \N__7316\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_2\
        );

    \I__819\ : InMux
    port map (
            O => \N__7313\,
            I => \N__7310\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__7310\,
            I => \N__7306\
        );

    \I__817\ : InMux
    port map (
            O => \N__7309\,
            I => \N__7303\
        );

    \I__816\ : Odrv4
    port map (
            O => \N__7306\,
            I => \rUartTxEnZ0\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__7303\,
            I => \rUartTxEnZ0\
        );

    \I__814\ : InMux
    port map (
            O => \N__7298\,
            I => \N__7295\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__7295\,
            I => \N__7292\
        );

    \I__812\ : Span4Mux_v
    port map (
            O => \N__7292\,
            I => \N__7289\
        );

    \I__811\ : Odrv4
    port map (
            O => \N__7289\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c3_0_0\
        );

    \I__810\ : CascadeMux
    port map (
            O => \N__7286\,
            I => \N__7283\
        );

    \I__809\ : InMux
    port map (
            O => \N__7283\,
            I => \N__7280\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__7280\,
            I => \N__7277\
        );

    \I__807\ : Span4Mux_v
    port map (
            O => \N__7277\,
            I => \N__7274\
        );

    \I__806\ : Odrv4
    port map (
            O => \N__7274\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c2_d\
        );

    \I__805\ : InMux
    port map (
            O => \N__7271\,
            I => \N__7267\
        );

    \I__804\ : InMux
    port map (
            O => \N__7270\,
            I => \N__7264\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__7267\,
            I => \N__7258\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__7264\,
            I => \N__7258\
        );

    \I__801\ : InMux
    port map (
            O => \N__7263\,
            I => \N__7255\
        );

    \I__800\ : Odrv12
    port map (
            O => \N__7258\,
            I => \uart_inst0.tx_uart_fifo_inst.rDataCount_0_sqmuxa\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__7255\,
            I => \uart_inst0.tx_uart_fifo_inst.rDataCount_0_sqmuxa\
        );

    \I__798\ : CascadeMux
    port map (
            O => \N__7250\,
            I => \uart_inst0.wTxRdEmpty_cascade_\
        );

    \I__797\ : InMux
    port map (
            O => \N__7247\,
            I => \N__7244\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__7244\,
            I => \N__7241\
        );

    \I__795\ : Span4Mux_h
    port map (
            O => \N__7241\,
            I => \N__7238\
        );

    \I__794\ : Span4Mux_h
    port map (
            O => \N__7238\,
            I => \N__7235\
        );

    \I__793\ : Odrv4
    port map (
            O => \N__7235\,
            I => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_0\
        );

    \I__792\ : InMux
    port map (
            O => \N__7232\,
            I => \N__7229\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__7229\,
            I => \N__7226\
        );

    \I__790\ : Span4Mux_h
    port map (
            O => \N__7226\,
            I => \N__7223\
        );

    \I__789\ : Span4Mux_h
    port map (
            O => \N__7223\,
            I => \N__7220\
        );

    \I__788\ : Odrv4
    port map (
            O => \N__7220\,
            I => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_1\
        );

    \I__787\ : InMux
    port map (
            O => \N__7217\,
            I => \N__7214\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__7214\,
            I => \N__7211\
        );

    \I__785\ : Span12Mux_h
    port map (
            O => \N__7211\,
            I => \N__7208\
        );

    \I__784\ : Odrv12
    port map (
            O => \N__7208\,
            I => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_2\
        );

    \I__783\ : CascadeMux
    port map (
            O => \N__7205\,
            I => \uart_inst0.tx_uart_fifo_inst.m65_bmZ0_cascade_\
        );

    \I__782\ : CascadeMux
    port map (
            O => \N__7202\,
            I => \fifo_inst.rx_fifo_inst.un1_rDataCount_c2_1_1_0_cascade_\
        );

    \I__781\ : InMux
    port map (
            O => \N__7199\,
            I => \N__7196\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__7196\,
            I => \uart_inst0.tx_uart_fifo_inst.m65_nsZ0Z_1\
        );

    \I__779\ : InMux
    port map (
            O => \N__7193\,
            I => \N__7190\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__7190\,
            I => \fifo_inst.rx_fifo_inst.un1_rDataCount_c2_1\
        );

    \I__777\ : CascadeMux
    port map (
            O => \N__7187\,
            I => \N__7184\
        );

    \I__776\ : InMux
    port map (
            O => \N__7184\,
            I => \N__7178\
        );

    \I__775\ : InMux
    port map (
            O => \N__7183\,
            I => \N__7178\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__7178\,
            I => \fifo_inst_rx_fifo_inst_rDataCount_0_sqmuxa\
        );

    \I__773\ : CascadeMux
    port map (
            O => \N__7175\,
            I => \N__7172\
        );

    \I__772\ : InMux
    port map (
            O => \N__7172\,
            I => \N__7169\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__7169\,
            I => \fifo_inst.rx_fifo_inst.un1_rDataCount_ac0_2\
        );

    \I__770\ : InMux
    port map (
            O => \N__7166\,
            I => \N__7163\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__7163\,
            I => \uart_inst0.tx_uart_fifo_inst.m78_bmZ0\
        );

    \I__768\ : CascadeMux
    port map (
            O => \N__7160\,
            I => \uart_inst0.tx_uart_fifo_inst.m78_nsZ0Z_1_cascade_\
        );

    \I__767\ : CEMux
    port map (
            O => \N__7157\,
            I => \N__7154\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__7154\,
            I => \N__7151\
        );

    \I__765\ : Odrv4
    port map (
            O => \N__7151\,
            I => \fifo_inst.ft2232h_inst.un1_rFifoState_12_0_i_0\
        );

    \I__764\ : CascadeMux
    port map (
            O => \N__7148\,
            I => \uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c2_d_cascade_\
        );

    \I__763\ : CascadeMux
    port map (
            O => \N__7145\,
            I => \N_84_mux_cascade_\
        );

    \I__762\ : CascadeMux
    port map (
            O => \N__7142\,
            I => \N__7139\
        );

    \I__761\ : InMux
    port map (
            O => \N__7139\,
            I => \N__7136\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__7136\,
            I => \N__7132\
        );

    \I__759\ : InMux
    port map (
            O => \N__7135\,
            I => \N__7128\
        );

    \I__758\ : Span4Mux_h
    port map (
            O => \N__7132\,
            I => \N__7125\
        );

    \I__757\ : InMux
    port map (
            O => \N__7131\,
            I => \N__7122\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__7128\,
            I => \N__7119\
        );

    \I__755\ : Odrv4
    port map (
            O => \N__7125\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_5\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__7122\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_5\
        );

    \I__753\ : Odrv4
    port map (
            O => \N__7119\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_5\
        );

    \I__752\ : InMux
    port map (
            O => \N__7112\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_4\
        );

    \I__751\ : CascadeMux
    port map (
            O => \N__7109\,
            I => \N__7106\
        );

    \I__750\ : InMux
    port map (
            O => \N__7106\,
            I => \N__7103\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__7103\,
            I => \N__7098\
        );

    \I__748\ : InMux
    port map (
            O => \N__7102\,
            I => \N__7095\
        );

    \I__747\ : InMux
    port map (
            O => \N__7101\,
            I => \N__7092\
        );

    \I__746\ : Odrv12
    port map (
            O => \N__7098\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_6\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__7095\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_6\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__7092\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_6\
        );

    \I__743\ : InMux
    port map (
            O => \N__7085\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_5\
        );

    \I__742\ : CascadeMux
    port map (
            O => \N__7082\,
            I => \N__7079\
        );

    \I__741\ : InMux
    port map (
            O => \N__7079\,
            I => \N__7075\
        );

    \I__740\ : InMux
    port map (
            O => \N__7078\,
            I => \N__7071\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__7075\,
            I => \N__7068\
        );

    \I__738\ : InMux
    port map (
            O => \N__7074\,
            I => \N__7065\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__7071\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_7\
        );

    \I__736\ : Odrv12
    port map (
            O => \N__7068\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_7\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__7065\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_7\
        );

    \I__734\ : InMux
    port map (
            O => \N__7058\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_6\
        );

    \I__733\ : InMux
    port map (
            O => \N__7055\,
            I => \bfn_13_3_0_\
        );

    \I__732\ : CascadeMux
    port map (
            O => \N__7052\,
            I => \N__7049\
        );

    \I__731\ : InMux
    port map (
            O => \N__7049\,
            I => \N__7046\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__7046\,
            I => \N__7042\
        );

    \I__729\ : CascadeMux
    port map (
            O => \N__7045\,
            I => \N__7039\
        );

    \I__728\ : Span4Mux_s2_v
    port map (
            O => \N__7042\,
            I => \N__7035\
        );

    \I__727\ : InMux
    port map (
            O => \N__7039\,
            I => \N__7032\
        );

    \I__726\ : InMux
    port map (
            O => \N__7038\,
            I => \N__7029\
        );

    \I__725\ : Span4Mux_h
    port map (
            O => \N__7035\,
            I => \N__7026\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__7032\,
            I => \N__7023\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__7029\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_8\
        );

    \I__722\ : Odrv4
    port map (
            O => \N__7026\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_8\
        );

    \I__721\ : Odrv4
    port map (
            O => \N__7023\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_8\
        );

    \I__720\ : CascadeMux
    port map (
            O => \N__7016\,
            I => \fifo_inst_ft2232h_inst_un1_rFifoState_12_0_i_cascade_\
        );

    \I__719\ : CascadeMux
    port map (
            O => \N__7013\,
            I => \N__7010\
        );

    \I__718\ : InMux
    port map (
            O => \N__7010\,
            I => \N__7007\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__7007\,
            I => \fifo_inst.tx_fifo_inst.un1_rDataCount_ac0_1_a1_1\
        );

    \I__716\ : CascadeMux
    port map (
            O => \N__7004\,
            I => \uart_inst0.tx_uart_fifo_inst.m68_eZ0Z_5_cascade_\
        );

    \I__715\ : InMux
    port map (
            O => \N__7001\,
            I => \N__6998\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__6998\,
            I => \uart_inst0.tx_uart_fifo_inst.m68_eZ0Z_6\
        );

    \I__713\ : InMux
    port map (
            O => \N__6995\,
            I => \N__6991\
        );

    \I__712\ : InMux
    port map (
            O => \N__6994\,
            I => \N__6988\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__6991\,
            I => \uart_inst0.tx_uart_fifo_inst.N_92\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__6988\,
            I => \uart_inst0.tx_uart_fifo_inst.N_92\
        );

    \I__709\ : CascadeMux
    port map (
            O => \N__6983\,
            I => \N__6980\
        );

    \I__708\ : InMux
    port map (
            O => \N__6980\,
            I => \N__6977\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__6977\,
            I => \N__6974\
        );

    \I__706\ : Span4Mux_v
    port map (
            O => \N__6974\,
            I => \N__6971\
        );

    \I__705\ : Span4Mux_h
    port map (
            O => \N__6971\,
            I => \N__6966\
        );

    \I__704\ : InMux
    port map (
            O => \N__6970\,
            I => \N__6963\
        );

    \I__703\ : InMux
    port map (
            O => \N__6969\,
            I => \N__6960\
        );

    \I__702\ : Odrv4
    port map (
            O => \N__6966\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_0\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__6963\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_0\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__6960\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_0\
        );

    \I__699\ : InMux
    port map (
            O => \N__6953\,
            I => \N__6950\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__6950\,
            I => \rRamWrAddr_RNI10581_0\
        );

    \I__697\ : CascadeMux
    port map (
            O => \N__6947\,
            I => \N__6944\
        );

    \I__696\ : InMux
    port map (
            O => \N__6944\,
            I => \N__6941\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__6941\,
            I => \N__6936\
        );

    \I__694\ : InMux
    port map (
            O => \N__6940\,
            I => \N__6933\
        );

    \I__693\ : InMux
    port map (
            O => \N__6939\,
            I => \N__6930\
        );

    \I__692\ : Odrv12
    port map (
            O => \N__6936\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_1\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__6933\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_1\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__6930\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_1\
        );

    \I__689\ : InMux
    port map (
            O => \N__6923\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_0\
        );

    \I__688\ : CascadeMux
    port map (
            O => \N__6920\,
            I => \N__6917\
        );

    \I__687\ : InMux
    port map (
            O => \N__6917\,
            I => \N__6914\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__6914\,
            I => \N__6911\
        );

    \I__685\ : Span4Mux_h
    port map (
            O => \N__6911\,
            I => \N__6906\
        );

    \I__684\ : InMux
    port map (
            O => \N__6910\,
            I => \N__6903\
        );

    \I__683\ : InMux
    port map (
            O => \N__6909\,
            I => \N__6900\
        );

    \I__682\ : Odrv4
    port map (
            O => \N__6906\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_2\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__6903\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_2\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__6900\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_2\
        );

    \I__679\ : InMux
    port map (
            O => \N__6893\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_1\
        );

    \I__678\ : CascadeMux
    port map (
            O => \N__6890\,
            I => \N__6887\
        );

    \I__677\ : InMux
    port map (
            O => \N__6887\,
            I => \N__6884\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__6884\,
            I => \N__6881\
        );

    \I__675\ : Span12Mux_v
    port map (
            O => \N__6881\,
            I => \N__6876\
        );

    \I__674\ : InMux
    port map (
            O => \N__6880\,
            I => \N__6873\
        );

    \I__673\ : InMux
    port map (
            O => \N__6879\,
            I => \N__6870\
        );

    \I__672\ : Odrv12
    port map (
            O => \N__6876\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_3\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__6873\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_3\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__6870\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_3\
        );

    \I__669\ : InMux
    port map (
            O => \N__6863\,
            I => \N__6860\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__6860\,
            I => \un1_rRamWrAddr_cry_2_c_RNISJKU\
        );

    \I__667\ : InMux
    port map (
            O => \N__6857\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_2\
        );

    \I__666\ : CascadeMux
    port map (
            O => \N__6854\,
            I => \N__6851\
        );

    \I__665\ : InMux
    port map (
            O => \N__6851\,
            I => \N__6847\
        );

    \I__664\ : CascadeMux
    port map (
            O => \N__6850\,
            I => \N__6844\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__6847\,
            I => \N__6840\
        );

    \I__662\ : InMux
    port map (
            O => \N__6844\,
            I => \N__6837\
        );

    \I__661\ : InMux
    port map (
            O => \N__6843\,
            I => \N__6834\
        );

    \I__660\ : Span12Mux_s1_v
    port map (
            O => \N__6840\,
            I => \N__6829\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__6837\,
            I => \N__6829\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__6834\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_4\
        );

    \I__657\ : Odrv12
    port map (
            O => \N__6829\,
            I => \fifo_inst_tx_fifo_inst_rRamWrAddr_4\
        );

    \I__656\ : InMux
    port map (
            O => \N__6824\,
            I => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_3\
        );

    \I__655\ : IoInMux
    port map (
            O => \N__6821\,
            I => \N__6817\
        );

    \I__654\ : IoInMux
    port map (
            O => \N__6820\,
            I => \N__6814\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__6817\,
            I => \N__6811\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__6814\,
            I => \N__6808\
        );

    \I__651\ : Span4Mux_s3_v
    port map (
            O => \N__6811\,
            I => \N__6805\
        );

    \I__650\ : Span4Mux_s1_v
    port map (
            O => \N__6808\,
            I => \N__6802\
        );

    \I__649\ : Span4Mux_h
    port map (
            O => \N__6805\,
            I => \N__6798\
        );

    \I__648\ : Span4Mux_h
    port map (
            O => \N__6802\,
            I => \N__6795\
        );

    \I__647\ : InMux
    port map (
            O => \N__6801\,
            I => \N__6792\
        );

    \I__646\ : Odrv4
    port map (
            O => \N__6798\,
            I => \P1A3_c\
        );

    \I__645\ : Odrv4
    port map (
            O => \N__6795\,
            I => \P1A3_c\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__6792\,
            I => \P1A3_c\
        );

    \I__643\ : InMux
    port map (
            O => \N__6785\,
            I => \N__6782\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__6782\,
            I => \N_86_mux\
        );

    \I__641\ : CascadeMux
    port map (
            O => \N__6779\,
            I => \uart_inst0.tx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_0_cascade_\
        );

    \I__640\ : InMux
    port map (
            O => \N__6776\,
            I => \N__6772\
        );

    \I__639\ : InMux
    port map (
            O => \N__6775\,
            I => \N__6769\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__6772\,
            I => \uart_inst0.tx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_6\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__6769\,
            I => \uart_inst0.tx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_6\
        );

    \I__636\ : IoInMux
    port map (
            O => \N__6764\,
            I => \N__6761\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__6761\,
            I => \GB_BUFFER_wPllLocked_i_g_THRU_CO\
        );

    \I__634\ : CascadeMux
    port map (
            O => \N__6758\,
            I => \fifo_inst_tx_fifo_inst_wRamWrEn_cascade_\
        );

    \I__633\ : InMux
    port map (
            O => \N__6755\,
            I => \N__6752\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__6752\,
            I => \uart_inst0.uart_inst0.un1_rx_clk_divider_10\
        );

    \I__631\ : InMux
    port map (
            O => \N__6749\,
            I => \N__6746\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__6746\,
            I => \uart_inst0.uart_inst0.un1_rx_clk_divider_9\
        );

    \I__629\ : CascadeMux
    port map (
            O => \N__6743\,
            I => \uart_inst0.uart_inst0.un1_rx_clk_divider_7_cascade_\
        );

    \I__628\ : CascadeMux
    port map (
            O => \N__6740\,
            I => \uart_inst0.uart_inst0.un1_rx_clk_divider_0_cascade_\
        );

    \I__627\ : InMux
    port map (
            O => \N__6737\,
            I => \N__6733\
        );

    \I__626\ : InMux
    port map (
            O => \N__6736\,
            I => \N__6730\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__6733\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_3\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__6730\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_3\
        );

    \I__623\ : InMux
    port map (
            O => \N__6725\,
            I => \N__6721\
        );

    \I__622\ : InMux
    port map (
            O => \N__6724\,
            I => \N__6718\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__6721\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_1\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__6718\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_1\
        );

    \I__619\ : CascadeMux
    port map (
            O => \N__6713\,
            I => \N__6709\
        );

    \I__618\ : InMux
    port map (
            O => \N__6712\,
            I => \N__6706\
        );

    \I__617\ : InMux
    port map (
            O => \N__6709\,
            I => \N__6703\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__6706\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_4\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__6703\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_4\
        );

    \I__614\ : InMux
    port map (
            O => \N__6698\,
            I => \N__6694\
        );

    \I__613\ : InMux
    port map (
            O => \N__6697\,
            I => \N__6691\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__6694\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_2\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__6691\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_2\
        );

    \I__610\ : InMux
    port map (
            O => \N__6686\,
            I => \N__6683\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__6683\,
            I => \uart_inst0.uart_inst0.un1_rx_clk_divider_8\
        );

    \I__608\ : InMux
    port map (
            O => \N__6680\,
            I => \N__6675\
        );

    \I__607\ : InMux
    port map (
            O => \N__6679\,
            I => \N__6672\
        );

    \I__606\ : InMux
    port map (
            O => \N__6678\,
            I => \N__6669\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__6675\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_0\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__6672\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_0\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__6669\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_0\
        );

    \I__602\ : SRMux
    port map (
            O => \N__6662\,
            I => \N__6657\
        );

    \I__601\ : SRMux
    port map (
            O => \N__6661\,
            I => \N__6654\
        );

    \I__600\ : SRMux
    port map (
            O => \N__6660\,
            I => \N__6651\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__6657\,
            I => \uart_inst0.uart_inst0.rx_clk_divider_1_sqmuxa_i\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__6654\,
            I => \uart_inst0.uart_inst0.rx_clk_divider_1_sqmuxa_i\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__6651\,
            I => \uart_inst0.uart_inst0.rx_clk_divider_1_sqmuxa_i\
        );

    \I__596\ : InMux
    port map (
            O => \N__6644\,
            I => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_8\
        );

    \I__595\ : InMux
    port map (
            O => \N__6641\,
            I => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_9\
        );

    \I__594\ : InMux
    port map (
            O => \N__6638\,
            I => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_10\
        );

    \I__593\ : InMux
    port map (
            O => \N__6635\,
            I => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_11\
        );

    \I__592\ : InMux
    port map (
            O => \N__6632\,
            I => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_12\
        );

    \I__591\ : InMux
    port map (
            O => \N__6629\,
            I => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_13\
        );

    \I__590\ : InMux
    port map (
            O => \N__6626\,
            I => \N__6622\
        );

    \I__589\ : InMux
    port map (
            O => \N__6625\,
            I => \N__6619\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__6622\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_8\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__6619\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_8\
        );

    \I__586\ : InMux
    port map (
            O => \N__6614\,
            I => \N__6610\
        );

    \I__585\ : InMux
    port map (
            O => \N__6613\,
            I => \N__6607\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__6610\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_7\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__6607\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_7\
        );

    \I__582\ : CascadeMux
    port map (
            O => \N__6602\,
            I => \N__6598\
        );

    \I__581\ : InMux
    port map (
            O => \N__6601\,
            I => \N__6595\
        );

    \I__580\ : InMux
    port map (
            O => \N__6598\,
            I => \N__6592\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__6595\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_14\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__6592\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_14\
        );

    \I__577\ : InMux
    port map (
            O => \N__6587\,
            I => \N__6583\
        );

    \I__576\ : InMux
    port map (
            O => \N__6586\,
            I => \N__6580\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__6583\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_10\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__6580\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_10\
        );

    \I__573\ : CascadeMux
    port map (
            O => \N__6575\,
            I => \N__6572\
        );

    \I__572\ : InMux
    port map (
            O => \N__6572\,
            I => \N__6568\
        );

    \I__571\ : InMux
    port map (
            O => \N__6571\,
            I => \N__6565\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__6568\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_11\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__6565\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_11\
        );

    \I__568\ : CascadeMux
    port map (
            O => \N__6560\,
            I => \N__6556\
        );

    \I__567\ : InMux
    port map (
            O => \N__6559\,
            I => \N__6553\
        );

    \I__566\ : InMux
    port map (
            O => \N__6556\,
            I => \N__6550\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__6553\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_12\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__6550\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_12\
        );

    \I__563\ : CascadeMux
    port map (
            O => \N__6545\,
            I => \N__6542\
        );

    \I__562\ : InMux
    port map (
            O => \N__6542\,
            I => \N__6538\
        );

    \I__561\ : InMux
    port map (
            O => \N__6541\,
            I => \N__6535\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__6538\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_9\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__6535\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_9\
        );

    \I__558\ : CascadeMux
    port map (
            O => \N__6530\,
            I => \N__6527\
        );

    \I__557\ : InMux
    port map (
            O => \N__6527\,
            I => \N__6523\
        );

    \I__556\ : InMux
    port map (
            O => \N__6526\,
            I => \N__6520\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__6523\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_13\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__6520\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_13\
        );

    \I__553\ : InMux
    port map (
            O => \N__6515\,
            I => \N__6511\
        );

    \I__552\ : InMux
    port map (
            O => \N__6514\,
            I => \N__6508\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__6511\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_6\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__6508\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_6\
        );

    \I__549\ : InMux
    port map (
            O => \N__6503\,
            I => \N__6499\
        );

    \I__548\ : InMux
    port map (
            O => \N__6502\,
            I => \N__6496\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__6499\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_5\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__6496\,
            I => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_5\
        );

    \I__545\ : InMux
    port map (
            O => \N__6491\,
            I => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_0\
        );

    \I__544\ : InMux
    port map (
            O => \N__6488\,
            I => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_1\
        );

    \I__543\ : InMux
    port map (
            O => \N__6485\,
            I => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_2\
        );

    \I__542\ : InMux
    port map (
            O => \N__6482\,
            I => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_3\
        );

    \I__541\ : InMux
    port map (
            O => \N__6479\,
            I => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_4\
        );

    \I__540\ : InMux
    port map (
            O => \N__6476\,
            I => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_5\
        );

    \I__539\ : InMux
    port map (
            O => \N__6473\,
            I => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_6\
        );

    \I__538\ : InMux
    port map (
            O => \N__6470\,
            I => \bfn_9_15_0_\
        );

    \I__537\ : InMux
    port map (
            O => \N__6467\,
            I => \N__6464\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__6464\,
            I => \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO\
        );

    \I__535\ : IoInMux
    port map (
            O => \N__6461\,
            I => \N__6458\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__6458\,
            I => \N__6455\
        );

    \I__533\ : Span12Mux_s9_v
    port map (
            O => \N__6455\,
            I => \N__6452\
        );

    \I__532\ : Span12Mux_v
    port map (
            O => \N__6452\,
            I => \N__6449\
        );

    \I__531\ : Odrv12
    port map (
            O => \N__6449\,
            I => \BTN_N_c\
        );

    \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_0C\ : INV
    port map (
            O => \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net\,
            I => \N__16957\
        );

    \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_5C\ : INV
    port map (
            O => \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_5C_net\,
            I => \N__16963\
        );

    \INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7C\ : INV
    port map (
            O => \INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7C_net\,
            I => \N__16980\
        );

    \INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_4C\ : INV
    port map (
            O => \INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_4C_net\,
            I => \N__16983\
        );

    \INVfifo_inst.tx_fifo_inst.ram512x8_inst.RDATA_0C\ : INV
    port map (
            O => \INVfifo_inst.tx_fifo_inst.ram512x8_inst.RDATA_0C_net\,
            I => \N__16977\
        );

    \INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0C\ : INV
    port map (
            O => \INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net\,
            I => \N__16924\
        );

    \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN\ : INV
    port map (
            O => \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net\,
            I => \N__16964\
        );

    \INVfifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN\ : INV
    port map (
            O => \INVfifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net\,
            I => \N__16986\
        );

    \INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN\ : INV
    port map (
            O => \INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net\,
            I => \N__16951\
        );

    \INVfifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN\ : INV
    port map (
            O => \INVfifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net\,
            I => \N__16991\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_7\,
            carryinitout => \bfn_9_15_0_\
        );

    \IN_MUX_bfv_16_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_15_0_\
        );

    \IN_MUX_bfv_16_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_18_0_\
        );

    \IN_MUX_bfv_16_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_7_s1\,
            carryinitout => \bfn_16_19_0_\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_12_0_\
        );

    \IN_MUX_bfv_13_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_7\,
            carryinitout => \bfn_13_13_0_\
        );

    \IN_MUX_bfv_14_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_11_0_\
        );

    \IN_MUX_bfv_14_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_7\,
            carryinitout => \bfn_14_12_0_\
        );

    \IN_MUX_bfv_17_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_6_0_\
        );

    \IN_MUX_bfv_17_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_7\,
            carryinitout => \bfn_17_7_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_7\,
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_13_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_2_0_\
        );

    \IN_MUX_bfv_13_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_7\,
            carryinitout => \bfn_13_3_0_\
        );

    \IN_MUX_bfv_15_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_3_0_\
        );

    \IN_MUX_bfv_15_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_7\,
            carryinitout => \bfn_15_4_0_\
        );

    \IN_MUX_bfv_17_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_2_0_\
        );

    \IN_MUX_bfv_17_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_7\,
            carryinitout => \bfn_17_3_0_\
        );

    \IN_MUX_bfv_15_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_5_0_\
        );

    \IN_MUX_bfv_15_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_7\,
            carryinitout => \bfn_15_6_0_\
        );

    \N_292_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__6764\,
            GLOBALBUFFEROUTPUT => \N_292_g\
        );

    \wPllLocked_i_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__14101\,
            GLOBALBUFFEROUTPUT => \wPllLocked_i_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6467\,
            lcout => \wPllLocked\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.wPllLocked_i_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13921\,
            lcout => \wPllLocked_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_0_c_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6679\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_clk_divider_1_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6725\,
            in2 => \N__12338\,
            in3 => \N__6491\,
            lcout => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_1\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_0\,
            carryout => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_1\,
            clk => \N__16923\,
            ce => 'H',
            sr => \N__6661\
        );

    \uart_inst0.uart_inst0.rx_clk_divider_2_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6698\,
            in2 => \N__12342\,
            in3 => \N__6488\,
            lcout => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_2\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_1\,
            carryout => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_2\,
            clk => \N__16923\,
            ce => 'H',
            sr => \N__6661\
        );

    \uart_inst0.uart_inst0.rx_clk_divider_3_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6737\,
            in2 => \N__12339\,
            in3 => \N__6485\,
            lcout => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_3\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_2\,
            carryout => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_3\,
            clk => \N__16923\,
            ce => 'H',
            sr => \N__6661\
        );

    \uart_inst0.uart_inst0.rx_clk_divider_4_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6712\,
            in2 => \N__12343\,
            in3 => \N__6482\,
            lcout => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_4\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_3\,
            carryout => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_4\,
            clk => \N__16923\,
            ce => 'H',
            sr => \N__6661\
        );

    \uart_inst0.uart_inst0.rx_clk_divider_5_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6503\,
            in2 => \N__12340\,
            in3 => \N__6479\,
            lcout => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_5\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_4\,
            carryout => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_5\,
            clk => \N__16923\,
            ce => 'H',
            sr => \N__6661\
        );

    \uart_inst0.uart_inst0.rx_clk_divider_6_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6515\,
            in2 => \N__12344\,
            in3 => \N__6476\,
            lcout => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_6\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_5\,
            carryout => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_6\,
            clk => \N__16923\,
            ce => 'H',
            sr => \N__6661\
        );

    \uart_inst0.uart_inst0.rx_clk_divider_7_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6614\,
            in2 => \N__12341\,
            in3 => \N__6473\,
            lcout => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_7\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_6\,
            carryout => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_7\,
            clk => \N__16923\,
            ce => 'H',
            sr => \N__6661\
        );

    \uart_inst0.uart_inst0.rx_clk_divider_8_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6626\,
            in2 => \N__12404\,
            in3 => \N__6470\,
            lcout => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_8\,
            clk => \N__16917\,
            ce => 'H',
            sr => \N__6662\
        );

    \uart_inst0.uart_inst0.rx_clk_divider_9_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12356\,
            in2 => \N__6545\,
            in3 => \N__6644\,
            lcout => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_9\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_8\,
            carryout => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_9\,
            clk => \N__16917\,
            ce => 'H',
            sr => \N__6662\
        );

    \uart_inst0.uart_inst0.rx_clk_divider_10_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6587\,
            in2 => \N__12402\,
            in3 => \N__6641\,
            lcout => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_10\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_9\,
            carryout => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_10\,
            clk => \N__16917\,
            ce => 'H',
            sr => \N__6662\
        );

    \uart_inst0.uart_inst0.rx_clk_divider_11_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12348\,
            in2 => \N__6575\,
            in3 => \N__6638\,
            lcout => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_11\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_10\,
            carryout => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_11\,
            clk => \N__16917\,
            ce => 'H',
            sr => \N__6662\
        );

    \uart_inst0.uart_inst0.rx_clk_divider_12_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6559\,
            in2 => \N__12403\,
            in3 => \N__6635\,
            lcout => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_12\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_11\,
            carryout => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_12\,
            clk => \N__16917\,
            ce => 'H',
            sr => \N__6662\
        );

    \uart_inst0.uart_inst0.rx_clk_divider_13_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12352\,
            in2 => \N__6530\,
            in3 => \N__6632\,
            lcout => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_13\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_12\,
            carryout => \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_13\,
            clk => \N__16917\,
            ce => 'H',
            sr => \N__6662\
        );

    \uart_inst0.uart_inst0.rx_clk_divider_14_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6601\,
            in2 => \_gnd_net_\,
            in3 => \N__6629\,
            lcout => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16917\,
            ce => 'H',
            sr => \N__6662\
        );

    \uart_inst0.uart_inst0.rx_clk_divider_RNI0H8H_14_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6625\,
            in1 => \N__6613\,
            in2 => \N__6602\,
            in3 => \N__6678\,
            lcout => \uart_inst0.uart_inst0.un1_rx_clk_divider_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_clk_divider_RNIRKBC1_9_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6586\,
            in1 => \N__6571\,
            in2 => \N__6560\,
            in3 => \N__6541\,
            lcout => \uart_inst0.uart_inst0.un1_rx_clk_divider_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_clk_divider_RNISPAG_5_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6526\,
            in1 => \N__6514\,
            in2 => \_gnd_net_\,
            in3 => \N__6502\,
            lcout => OPEN,
            ltout => \uart_inst0.uart_inst0.un1_rx_clk_divider_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_clk_divider_RNITHLH2_1_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6755\,
            in1 => \N__6749\,
            in2 => \N__6743\,
            in3 => \N__6686\,
            lcout => \uart_inst0.uart_inst0.un1_rx_clk_divider_0\,
            ltout => \uart_inst0.uart_inst0.un1_rx_clk_divider_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_state_RNIPLGK2_0_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__13894\,
            in1 => \_gnd_net_\,
            in2 => \N__6740\,
            in3 => \N__11155\,
            lcout => \uart_inst0.uart_inst0.rx_clk_divider_1_sqmuxa_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_clk_divider_RNI6IM3_1_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6736\,
            in1 => \N__6724\,
            in2 => \N__6713\,
            in3 => \N__6697\,
            lcout => \uart_inst0.uart_inst0.un1_rx_clk_divider_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_clk_divider_0_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6680\,
            lcout => \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16909\,
            ce => 'H',
            sr => \N__6660\
        );

    \fifo_inst.tx_fifo_inst.rDataCount_3_LC_12_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__7966\,
            in1 => \N__7866\,
            in2 => \N__7951\,
            in3 => \N__10161\,
            lcout => \wTxFull\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16958\,
            ce => 'H',
            sr => \N__16340\
        );

    \rTxEn_LC_12_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10160\,
            lcout => \rTxEnZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16958\,
            ce => 'H',
            sr => \N__16340\
        );

    \fifo_inst.tx_fifo_inst.rDataCount_RNIA7U81_2_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__7825\,
            in1 => \N__7787\,
            in2 => \N__9259\,
            in3 => \N__7721\,
            lcout => \fifo_inst.tx_fifo_inst.un1_rDataCount_axbxc3_2_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rDataCount_RNIEM211_2_LC_12_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__9303\,
            in1 => \N__9251\,
            in2 => \_gnd_net_\,
            in3 => \N__7826\,
            lcout => \fifo_inst.tx_fifo_inst.un1_rDataCount_axbxc3_a0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rDataCount_RNIDPRL_0_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7786\,
            in2 => \_gnd_net_\,
            in3 => \N__7720\,
            lcout => \fifo_inst.tx_fifo_inst.un1_rDataCount_ac0_1_a0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ft2232h_inst.rRx_n_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__6801\,
            in1 => \N__6785\,
            in2 => \_gnd_net_\,
            in3 => \N__8150\,
            lcout => \P1A3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16946\,
            ce => 'H',
            sr => \N__16350\
        );

    \uart_inst0.tx_uart_fifo_inst.m39_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__8116\,
            in1 => \N__8078\,
            in2 => \_gnd_net_\,
            in3 => \N__12764\,
            lcout => \N_86_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_3_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__6776\,
            in1 => \N__7322\,
            in2 => \N__8645\,
            in3 => \N__8505\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16918\,
            ce => 'H',
            sr => \N__13595\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNIVHG3_8_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7563\,
            in2 => \_gnd_net_\,
            in3 => \N__7338\,
            lcout => OPEN,
            ltout => \uart_inst0.tx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNI0VO8_0_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__7375\,
            in1 => \N__7405\,
            in2 => \N__6779\,
            in3 => \N__7435\,
            lcout => \uart_inst0.tx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ0Z_0_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__6775\,
            in1 => \N__7415\,
            in2 => \N__8644\,
            in3 => \N__8515\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16908\,
            ce => 'H',
            sr => \N__13593\
        );

    \GB_BUFFER_wPllLocked_i_g_THRU_LUT4_0_LC_12_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__16696\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_wPllLocked_i_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rDataCount_RNIQ7UO_3_LC_13_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10143\,
            in2 => \_gnd_net_\,
            in3 => \N__9288\,
            lcout => \fifo_inst_tx_fifo_inst_wRamWrEn\,
            ltout => \fifo_inst_tx_fifo_inst_wRamWrEn_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamWrAddr_3_LC_13_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001101100000000"
        )
    port map (
            in0 => \N__6995\,
            in1 => \N__16619\,
            in2 => \N__6758\,
            in3 => \N__6863\,
            lcout => \fifo_inst_tx_fifo_inst_rRamWrAddr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16971\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamWrAddr_0_LC_13_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000101010"
        )
    port map (
            in0 => \N__6953\,
            in1 => \N__6994\,
            in2 => \N__7923\,
            in3 => \N__16618\,
            lcout => \fifo_inst_tx_fifo_inst_rRamWrAddr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16971\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m68_e_6_LC_13_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__6879\,
            in1 => \N__6939\,
            in2 => \N__7045\,
            in3 => \N__6969\,
            lcout => \uart_inst0.tx_uart_fifo_inst.m68_eZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m68_e_5_LC_13_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7135\,
            in1 => \N__16620\,
            in2 => \N__6854\,
            in3 => \N__6909\,
            lcout => OPEN,
            ltout => \uart_inst0.tx_uart_fifo_inst.m68_eZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m68_e_LC_13_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__7074\,
            in1 => \N__7101\,
            in2 => \N__7004\,
            in3 => \N__7001\,
            lcout => \uart_inst0.tx_uart_fifo_inst.N_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamWrAddr_RNI10581_0_LC_13_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6970\,
            in2 => \N__7919\,
            in3 => \N__7918\,
            lcout => \rRamWrAddr_RNI10581_0\,
            ltout => OPEN,
            carryin => \bfn_13_2_0_\,
            carryout => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamWrAddr_1_LC_13_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16621\,
            in1 => \N__6940\,
            in2 => \_gnd_net_\,
            in3 => \N__6923\,
            lcout => \fifo_inst_tx_fifo_inst_rRamWrAddr_1\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_0\,
            carryout => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_1\,
            clk => \N__16966\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamWrAddr_2_LC_13_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16624\,
            in1 => \N__6910\,
            in2 => \_gnd_net_\,
            in3 => \N__6893\,
            lcout => \fifo_inst_tx_fifo_inst_rRamWrAddr_2\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_1\,
            carryout => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_2\,
            clk => \N__16966\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_2_c_RNISJKU_LC_13_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6880\,
            in2 => \_gnd_net_\,
            in3 => \N__6857\,
            lcout => \un1_rRamWrAddr_cry_2_c_RNISJKU\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_2\,
            carryout => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamWrAddr_4_LC_13_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16625\,
            in1 => \N__6843\,
            in2 => \_gnd_net_\,
            in3 => \N__6824\,
            lcout => \fifo_inst_tx_fifo_inst_rRamWrAddr_4\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_3\,
            carryout => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_4\,
            clk => \N__16966\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamWrAddr_5_LC_13_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16622\,
            in1 => \N__7131\,
            in2 => \_gnd_net_\,
            in3 => \N__7112\,
            lcout => \fifo_inst_tx_fifo_inst_rRamWrAddr_5\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_4\,
            carryout => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_5\,
            clk => \N__16966\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamWrAddr_6_LC_13_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16626\,
            in1 => \N__7102\,
            in2 => \_gnd_net_\,
            in3 => \N__7085\,
            lcout => \fifo_inst_tx_fifo_inst_rRamWrAddr_6\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_5\,
            carryout => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_6\,
            clk => \N__16966\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamWrAddr_7_LC_13_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16623\,
            in1 => \N__7078\,
            in2 => \_gnd_net_\,
            in3 => \N__7058\,
            lcout => \fifo_inst_tx_fifo_inst_rRamWrAddr_7\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_6\,
            carryout => \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_7\,
            clk => \N__16966\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamWrAddr_8_LC_13_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16627\,
            in1 => \N__7038\,
            in2 => \_gnd_net_\,
            in3 => \N__7055\,
            lcout => \fifo_inst_tx_fifo_inst_rRamWrAddr_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16959\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rDataCount_RNO_3_2_LC_13_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9239\,
            in2 => \_gnd_net_\,
            in3 => \N__7772\,
            lcout => \fifo_inst.tx_fifo_inst.un1_rDataCount_ac0_1_a1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.un1_rFifoState_12_0_i_LC_13_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001110"
        )
    port map (
            in0 => \N__10636\,
            in1 => \N__8258\,
            in2 => \N__10613\,
            in3 => \N__10499\,
            lcout => OPEN,
            ltout => \fifo_inst_ft2232h_inst_un1_rFifoState_12_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ft2232h_inst.rTxRdEn_esr_RNO_LC_13_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7016\,
            in3 => \N__14102\,
            lcout => \fifo_inst.ft2232h_inst.un1_rFifoState_12_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m78_bm_LC_13_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__7815\,
            in1 => \N__7773\,
            in2 => \N__10162\,
            in3 => \N__7717\,
            lcout => \uart_inst0.tx_uart_fifo_inst.m78_bmZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rDataCount_RNO_2_2_LC_13_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000000000"
        )
    port map (
            in0 => \N__10147\,
            in1 => \N__9295\,
            in2 => \N__7013\,
            in3 => \N__7718\,
            lcout => \fifo_inst.tx_fifo_inst.un1_rDataCount_c2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m78_ns_1_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101000100"
        )
    port map (
            in0 => \N__10163\,
            in1 => \N__9302\,
            in2 => \_gnd_net_\,
            in3 => \N__9257\,
            lcout => OPEN,
            ltout => \uart_inst0.tx_uart_fifo_inst.m78_nsZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m78_ns_LC_13_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__9258\,
            in1 => \N__7166\,
            in2 => \N__7160\,
            in3 => \N__10523\,
            lcout => \fifo_inst_tx_fifo_inst_un1_rDataCount15_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ft2232h_inst.rTxRdEn_esr_LC_13_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__10608\,
            in1 => \N__10656\,
            in2 => \_gnd_net_\,
            in3 => \N__10524\,
            lcout => \fifo_inst_wTxRdEn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16952\,
            ce => \N__7157\,
            sr => \N__16355\
        );

    \uart_inst0.tx_uart_fifo_inst.rDataCount_RNI1JE32_0_LC_13_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010010100000"
        )
    port map (
            in0 => \N__8491\,
            in1 => \N__8419\,
            in2 => \N__8360\,
            in3 => \N__9509\,
            lcout => \uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c2_d\,
            ltout => \uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c2_d_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.rDataCount_RNO_0_3_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__8420\,
            in1 => \N__7263\,
            in2 => \N__7148\,
            in3 => \N__8387\,
            lcout => \uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIO6DU2_3_LC_13_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100000000"
        )
    port map (
            in0 => \N__7313\,
            in1 => \N__8316\,
            in2 => \N__9850\,
            in3 => \N__9508\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rDataCount_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m14_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8221\,
            in1 => \N__12689\,
            in2 => \N__8039\,
            in3 => \N__12587\,
            lcout => \N_84_mux\,
            ltout => \N_84_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m17_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101000000010"
        )
    port map (
            in0 => \N__15364\,
            in1 => \N__9074\,
            in2 => \N__7145\,
            in3 => \N__12757\,
            lcout => \fifo_inst_rx_fifo_inst_rDataCount_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m65_bm_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__12755\,
            in1 => \N__12690\,
            in2 => \N__12650\,
            in3 => \N__12588\,
            lcout => OPEN,
            ltout => \uart_inst0.tx_uart_fifo_inst.m65_bmZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m65_ns_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100100110001"
        )
    port map (
            in0 => \N__15365\,
            in1 => \N__7199\,
            in2 => \N__7205\,
            in3 => \N__8199\,
            lcout => \fifo_inst_rx_fifo_inst_un1_rDataCount15_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rDataCount_RNO_2_2_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__12756\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9073\,
            lcout => OPEN,
            ltout => \fifo_inst.rx_fifo_inst.un1_rDataCount_c2_1_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rDataCount_RNO_1_2_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001000000000"
        )
    port map (
            in0 => \N__15367\,
            in1 => \N__12592\,
            in2 => \N__7202\,
            in3 => \N__12637\,
            lcout => \fifo_inst.rx_fifo_inst.un1_rDataCount_c2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m65_ns_1_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101000100"
        )
    port map (
            in0 => \N__12754\,
            in1 => \N__9072\,
            in2 => \_gnd_net_\,
            in3 => \N__15363\,
            lcout => \uart_inst0.tx_uart_fifo_inst.m65_nsZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rDataCount_RNO_0_2_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010100000"
        )
    port map (
            in0 => \N__15366\,
            in1 => \N__12758\,
            in2 => \N__12598\,
            in3 => \N__9075\,
            lcout => \fifo_inst.rx_fifo_inst.un1_rDataCount_ac0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rDataCount_1_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100101110110100"
        )
    port map (
            in0 => \N__8237\,
            in1 => \N__12646\,
            in2 => \N__7187\,
            in3 => \N__12594\,
            lcout => \fifo_inst_rx_fifo_inst_rDataCount_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16941\,
            ce => 'H',
            sr => \N__16366\
        );

    \fifo_inst.rx_fifo_inst.rDataCount_2_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100100110110"
        )
    port map (
            in0 => \N__7193\,
            in1 => \N__7183\,
            in2 => \N__7175\,
            in3 => \N__12691\,
            lcout => \fifo_inst_rx_fifo_inst_rDataCount_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16941\,
            ce => 'H',
            sr => \N__16366\
        );

    \rUartTxEn_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__11217\,
            in1 => \N__15376\,
            in2 => \_gnd_net_\,
            in3 => \N__8318\,
            lcout => \rUartTxEnZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16938\,
            ce => 'H',
            sr => \N__16384\
        );

    \rUartRxFlag_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13049\,
            lcout => \rUartRxFlagZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16938\,
            ce => 'H',
            sr => \N__16384\
        );

    \CONSTANT_ONE_LUT4_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIPA3Q_3_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7309\,
            in2 => \_gnd_net_\,
            in3 => \N__8301\,
            lcout => \uart_inst0.tx_uart_fifo_inst.wRamWrEn_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.rDataCountZ0Z_0_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101100110100110"
        )
    port map (
            in0 => \N__8475\,
            in1 => \N__9499\,
            in2 => \N__9848\,
            in3 => \N__8356\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16930\,
            ce => 'H',
            sr => \N__16413\
        );

    \uart_inst0.tx_uart_fifo_inst.rDataCount_3_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100101000110"
        )
    port map (
            in0 => \N__7270\,
            in1 => \N__7298\,
            in2 => \N__7286\,
            in3 => \N__8314\,
            lcout => \uart_inst0.tx_uart_fifo_inst.wUartTxFull\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16930\,
            ce => 'H',
            sr => \N__16413\
        );

    \uart_inst0.tx_uart_fifo_inst.rDataCount_2_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__8522\,
            in1 => \N__7271\,
            in2 => \_gnd_net_\,
            in3 => \N__8382\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rDataCountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16926\,
            ce => 'H',
            sr => \N__16415\
        );

    \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIA3TL1_2_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8381\,
            in1 => \N__8351\,
            in2 => \N__8315\,
            in3 => \N__8410\,
            lcout => \uart_inst0.wTxRdEmpty\,
            ltout => \uart_inst0.wTxRdEmpty_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rTxRdEn_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100000001"
        )
    port map (
            in0 => \N__11591\,
            in1 => \N__11669\,
            in2 => \N__7250\,
            in3 => \N__9500\,
            lcout => \uart_inst0.wTxRdEn_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16926\,
            ce => 'H',
            sr => \N__16415\
        );

    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7247\,
            lcout => \uart_inst0.wTxRdData_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net\,
            ce => \N__9593\,
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_1_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7232\,
            lcout => \uart_inst0.wTxRdData_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net\,
            ce => \N__9593\,
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_2_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7217\,
            lcout => \uart_inst0.wTxRdData_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net\,
            ce => \N__9593\,
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_3_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7505\,
            lcout => \uart_inst0.wTxRdData_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net\,
            ce => \N__9593\,
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_4_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7490\,
            lcout => \uart_inst0.wTxRdData_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net\,
            ce => \N__9593\,
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_5_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7478\,
            lcout => \uart_inst0.wTxRdData_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net\,
            ce => \N__9593\,
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_6_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7466\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart_inst0.wTxRdData_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net\,
            ce => \N__9593\,
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_7_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7457\,
            lcout => \uart_inst0.wTxRdData_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net\,
            ce => \N__9593\,
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNO_0_0_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7431\,
            in2 => \N__8516\,
            in3 => \N__8514\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_13_12_0_\,
            carryout => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ0Z_1_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7401\,
            in2 => \_gnd_net_\,
            in3 => \N__7385\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ1Z_1\,
            ltout => OPEN,
            carryin => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_0\,
            carryout => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_1\,
            clk => \N__16919\,
            ce => 'H',
            sr => \N__13596\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_2_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7371\,
            in2 => \_gnd_net_\,
            in3 => \N__7355\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ0Z_2\,
            ltout => OPEN,
            carryin => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_1\,
            carryout => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_2\,
            clk => \N__16919\,
            ce => 'H',
            sr => \N__13596\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNO_0_3_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7339\,
            in2 => \_gnd_net_\,
            in3 => \N__7316\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_2\,
            carryout => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_4_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8661\,
            in2 => \_gnd_net_\,
            in3 => \N__7592\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_4\,
            ltout => OPEN,
            carryin => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_3\,
            carryout => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_4\,
            clk => \N__16919\,
            ce => 'H',
            sr => \N__13596\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_5_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8712\,
            in2 => \_gnd_net_\,
            in3 => \N__7589\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_5\,
            ltout => OPEN,
            carryin => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_4\,
            carryout => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_5\,
            clk => \N__16919\,
            ce => 'H',
            sr => \N__13596\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_6_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8685\,
            in2 => \_gnd_net_\,
            in3 => \N__7586\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_6\,
            ltout => OPEN,
            carryin => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_5\,
            carryout => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_6\,
            clk => \N__16919\,
            ce => 'H',
            sr => \N__13596\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_7_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8742\,
            in2 => \_gnd_net_\,
            in3 => \N__7583\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_7\,
            ltout => OPEN,
            carryin => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_6\,
            carryout => \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_7\,
            clk => \N__16919\,
            ce => 'H',
            sr => \N__13596\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_8_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7567\,
            in2 => \_gnd_net_\,
            in3 => \N__7580\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16913\,
            ce => 'H',
            sr => \N__13594\
        );

    \uart_inst0.uart_inst0.rTxData_esr_0_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__7529\,
            in1 => \N__8574\,
            in2 => \_gnd_net_\,
            in3 => \N__7547\,
            lcout => \uart_inst0.uart_inst0.rTxDataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16910\,
            ce => \N__8813\,
            sr => \N__16436\
        );

    \uart_inst0.uart_inst0.rTxData_esr_1_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__7646\,
            in1 => \N__8575\,
            in2 => \_gnd_net_\,
            in3 => \N__7538\,
            lcout => \uart_inst0.uart_inst0.rTxDataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16910\,
            ce => \N__8813\,
            sr => \N__16436\
        );

    \uart_inst0.uart_inst0.rTxData_esr_6_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7523\,
            in1 => \N__7606\,
            in2 => \_gnd_net_\,
            in3 => \N__8584\,
            lcout => \uart_inst0.uart_inst0.rTxDataZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16904\,
            ce => \N__8806\,
            sr => \N__16437\
        );

    \uart_inst0.uart_inst0.rTxData_esr_3_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__7667\,
            in1 => \N__8581\,
            in2 => \_gnd_net_\,
            in3 => \N__7514\,
            lcout => \uart_inst0.uart_inst0.rTxDataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16904\,
            ce => \N__8806\,
            sr => \N__16437\
        );

    \uart_inst0.uart_inst0.rTxData_esr_4_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8582\,
            in1 => \N__7625\,
            in2 => \_gnd_net_\,
            in3 => \N__7679\,
            lcout => \uart_inst0.uart_inst0.rTxDataZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16904\,
            ce => \N__8806\,
            sr => \N__16437\
        );

    \uart_inst0.uart_inst0.rTxData_esr_2_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__7661\,
            in1 => \N__8580\,
            in2 => \_gnd_net_\,
            in3 => \N__7655\,
            lcout => \uart_inst0.uart_inst0.rTxDataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16904\,
            ce => \N__8806\,
            sr => \N__16437\
        );

    \uart_inst0.uart_inst0.rTxData_esr_5_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8583\,
            in1 => \N__7640\,
            in2 => \_gnd_net_\,
            in3 => \N__7634\,
            lcout => \uart_inst0.uart_inst0.rTxDataZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16904\,
            ce => \N__8806\,
            sr => \N__16437\
        );

    \uart_inst0.uart_inst0.rTxData_7_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__8562\,
            in1 => \N__7619\,
            in2 => \N__7610\,
            in3 => \N__8822\,
            lcout => \uart_inst0.uart_inst0.rTxDataZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16900\,
            ce => 'H',
            sr => \N__16448\
        );

    \uart_inst0.uart_inst0.tx_bits_remaining_3_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111111101010"
        )
    port map (
            in0 => \N__8585\,
            in1 => \N__8777\,
            in2 => \N__8795\,
            in3 => \N__9766\,
            lcout => \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16897\,
            ce => 'H',
            sr => \N__16453\
        );

    \fifo_inst.ft2232h_inst.rFifoState_RNIM35O_0_LC_14_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__8117\,
            in1 => \N__8067\,
            in2 => \_gnd_net_\,
            in3 => \N__12750\,
            lcout => \N_97\,
            ltout => \N_97_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ft2232h_inst.rFifoState_0_LC_14_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111001110110011"
        )
    port map (
            in0 => \N__10609\,
            in1 => \N__8162\,
            in2 => \N__7595\,
            in3 => \N__10525\,
            lcout => \fifo_inst_ft2232h_inst_rFifoState_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16972\,
            ce => 'H',
            sr => \N__16351\
        );

    \uart_inst0.tx_uart_fifo_inst.m8_x0_LC_14_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__7769\,
            in1 => \N__7709\,
            in2 => \N__7819\,
            in3 => \N__9237\,
            lcout => OPEN,
            ltout => \uart_inst0.tx_uart_fifo_inst.m8_xZ0Z0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m8_ns_LC_14_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__9238\,
            in1 => \_gnd_net_\,
            in2 => \N__7973\,
            in3 => \N__7734\,
            lcout => \fifo_inst_tx_fifo_inst_wRamRdEn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rDataCount_fast_3_LC_14_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__7735\,
            in1 => \N__7970\,
            in2 => \N__7955\,
            in3 => \N__7873\,
            lcout => \fifo_inst_tx_fifo_inst_rDataCount_fast_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16967\,
            ce => 'H',
            sr => \N__16356\
        );

    \fifo_inst.tx_fifo_inst.rDataCount_0_LC_14_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__7710\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7837\,
            lcout => \fifo_inst_tx_fifo_inst_rDataCount_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16967\,
            ce => 'H',
            sr => \N__16356\
        );

    \fifo_inst.tx_fifo_inst.rDataCount_RNO_1_2_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101010"
        )
    port map (
            in0 => \N__7934\,
            in1 => \N__7927\,
            in2 => \N__7877\,
            in3 => \N__9253\,
            lcout => OPEN,
            ltout => \fifo_inst.tx_fifo_inst.un1_rDataCount_c2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rDataCount_2_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100101010110"
        )
    port map (
            in0 => \N__7814\,
            in1 => \N__7844\,
            in2 => \N__7847\,
            in3 => \N__9202\,
            lcout => \fifo_inst_tx_fifo_inst_rDataCount_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16960\,
            ce => 'H',
            sr => \N__16358\
        );

    \fifo_inst.tx_fifo_inst.rDataCount_RNO_0_2_LC_14_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001000000000"
        )
    port map (
            in0 => \N__7771\,
            in1 => \N__9311\,
            in2 => \N__10178\,
            in3 => \N__9252\,
            lcout => \fifo_inst.tx_fifo_inst.un1_rDataCount_ac0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rDataCount_1_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110010010110"
        )
    port map (
            in0 => \N__7719\,
            in1 => \N__9203\,
            in2 => \N__7785\,
            in3 => \N__7838\,
            lcout => \fifo_inst_tx_fifo_inst_rDataCount_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16960\,
            ce => 'H',
            sr => \N__16358\
        );

    \uart_inst0.tx_uart_fifo_inst.m7_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7813\,
            in1 => \N__7770\,
            in2 => \N__7739\,
            in3 => \N__7711\,
            lcout => \N_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rDataCount_RNILHIG_0_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000001010"
        )
    port map (
            in0 => \N__15362\,
            in1 => \N__9076\,
            in2 => \N__12651\,
            in3 => \N__12593\,
            lcout => \fifo_inst.rx_fifo_inst.un1_rDataCount_axbxc3_1_1\,
            ltout => \fifo_inst.rx_fifo_inst.un1_rDataCount_axbxc3_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rDataCount_3_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111110000000"
        )
    port map (
            in0 => \N__12687\,
            in1 => \N__12641\,
            in2 => \N__8051\,
            in3 => \N__12749\,
            lcout => \fifo_inst_wRxWrFull\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16953\,
            ce => 'H',
            sr => \N__16367\
        );

    \fifo_inst.ft2232h_inst.rRxWrEn_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__9077\,
            in1 => \N__17028\,
            in2 => \_gnd_net_\,
            in3 => \N__8146\,
            lcout => \fifo_inst_wRxWrEn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16953\,
            ce => 'H',
            sr => \N__16367\
        );

    \uart_inst0.tx_uart_fifo_inst.m15_x0_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__12586\,
            in1 => \N__12686\,
            in2 => \N__15377\,
            in3 => \N__8220\,
            lcout => OPEN,
            ltout => \uart_inst0.tx_uart_fifo_inst.m15_xZ0Z0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m15_ns_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8034\,
            in2 => \N__8048\,
            in3 => \N__15361\,
            lcout => \fifo_inst_rx_fifo_inst_wRamRdEn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rDataCount_fast_3_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101010100010"
        )
    port map (
            in0 => \N__8035\,
            in1 => \N__8045\,
            in2 => \N__12652\,
            in3 => \N__12688\,
            lcout => \fifo_inst_rx_fifo_inst_rDataCount_fast_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16953\,
            ce => 'H',
            sr => \N__16367\
        );

    \fifo_inst.ft2232h_inst.rFifoState_4_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100001010"
        )
    port map (
            in0 => \N__9160\,
            in1 => \_gnd_net_\,
            in2 => \N__9188\,
            in3 => \N__8256\,
            lcout => \fifo_inst_ft2232h_inst_rFifoState_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16947\,
            ce => 'H',
            sr => \N__16385\
        );

    \rRxEn_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__8200\,
            in1 => \N__8179\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \P1A2_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16947\,
            ce => 'H',
            sr => \N__16385\
        );

    \fifo_inst.ft2232h_inst.rWrDelay_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9183\,
            in2 => \_gnd_net_\,
            in3 => \N__9159\,
            lcout => \fifo_inst_ft2232h_inst_rWrDelay\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16947\,
            ce => 'H',
            sr => \N__16385\
        );

    \fifo_inst.ft2232h_inst.rTx_n_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__7989\,
            in1 => \N__8257\,
            in2 => \_gnd_net_\,
            in3 => \N__10672\,
            lcout => \P1A4_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16947\,
            ce => 'H',
            sr => \N__16385\
        );

    \fifo_inst.rx_fifo_inst.rDataCount_0_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8235\,
            in2 => \_gnd_net_\,
            in3 => \N__12645\,
            lcout => \fifo_inst_rx_fifo_inst_rDataCount_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16947\,
            ce => 'H',
            sr => \N__16385\
        );

    \fifo_inst.ft2232h_inst.rFifoState_3_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__10600\,
            in1 => \N__10658\,
            in2 => \_gnd_net_\,
            in3 => \N__10530\,
            lcout => \fifo_inst_ft2232h_inst_rFifoState_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16947\,
            ce => 'H',
            sr => \N__16385\
        );

    \fifo_inst.rx_fifo_inst.rDataCount_fast_0_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8236\,
            in2 => \_gnd_net_\,
            in3 => \N__8222\,
            lcout => \fifo_inst_rx_fifo_inst_rDataCount_fast_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16947\,
            ce => 'H',
            sr => \N__16385\
        );

    \rFtdiRxState_0_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__8204\,
            in1 => \_gnd_net_\,
            in2 => \N__8180\,
            in3 => \N__14015\,
            lcout => \rFtdiRxStateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16942\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.rDataCount_RNID3RQ_3_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__11216\,
            in1 => \N__15368\,
            in2 => \_gnd_net_\,
            in3 => \N__8317\,
            lcout => OPEN,
            ltout => \rUartTxEn_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.rDataCount_RNI9H5T_3_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8183\,
            in3 => \N__16674\,
            lcout => \rUartTxEn_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m27_e_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__14016\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8175\,
            lcout => \N_27_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ft2232h_inst.rFifoState_RNO_0_0_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__8133\,
            in1 => \N__9187\,
            in2 => \_gnd_net_\,
            in3 => \N__9161\,
            lcout => \fifo_inst.ft2232h_inst.rFifoStatesr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ft2232h_inst.rFifoState_2_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17027\,
            lcout => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16933\,
            ce => 'H',
            sr => \N__16416\
        );

    \fifo_inst.ft2232h_inst.rFifoState_1_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__8103\,
            in1 => \N__8077\,
            in2 => \_gnd_net_\,
            in3 => \N__12762\,
            lcout => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16933\,
            ce => 'H',
            sr => \N__16416\
        );

    \uart_inst0.tx_uart_fifo_inst.rDataCountZ0Z_1_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011010001111000"
        )
    port map (
            in0 => \N__8476\,
            in1 => \N__8355\,
            in2 => \N__8429\,
            in3 => \N__9591\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16933\,
            ce => 'H',
            sr => \N__16416\
        );

    \uart_inst0.tx_uart_fifo_inst.rDataCount_RNO_0_2_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101000001000"
        )
    port map (
            in0 => \N__9489\,
            in1 => \N__8408\,
            in2 => \N__8509\,
            in3 => \N__8350\,
            lcout => \uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.rDataCount_RNO_0_1_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010011010"
        )
    port map (
            in0 => \N__8409\,
            in1 => \N__9832\,
            in2 => \N__9506\,
            in3 => \N__8492\,
            lcout => \uart_inst0.tx_uart_fifo_inst.un1_rDataCount_axbxc1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIJHQM1_2_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__9487\,
            in1 => \N__8407\,
            in2 => \N__8386\,
            in3 => \N__8349\,
            lcout => OPEN,
            ltout => \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIJHQM1Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIKKMI2_3_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9488\,
            in2 => \N__8321\,
            in3 => \N__8300\,
            lcout => \uart_inst0.tx_uart_fifo_inst.wRamRdEn_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIBDOK2_0_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9415\,
            in2 => \N__9592\,
            in3 => \N__9587\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIBDOK2Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_14_11_0_\,
            carryout => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIOA54_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11315\,
            in2 => \_gnd_net_\,
            in3 => \N__8267\,
            lcout => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIOAZ0Z54\,
            ltout => OPEN,
            carryin => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_0\,
            carryout => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIQD64_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11300\,
            in3 => \N__8264\,
            lcout => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIQDZ0Z64\,
            ltout => OPEN,
            carryin => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_1\,
            carryout => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNISG74_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9403\,
            in2 => \_gnd_net_\,
            in3 => \N__8261\,
            lcout => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNISGZ0Z74\,
            ltout => OPEN,
            carryin => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_2\,
            carryout => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIUJ84_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9709\,
            in2 => \_gnd_net_\,
            in3 => \N__8762\,
            lcout => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIUJZ0Z84\,
            ltout => OPEN,
            carryin => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_3\,
            carryout => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNI0N94_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9694\,
            in2 => \_gnd_net_\,
            in3 => \N__8759\,
            lcout => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNI0NZ0Z94\,
            ltout => OPEN,
            carryin => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_4\,
            carryout => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNI2QA4_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9667\,
            in2 => \_gnd_net_\,
            in3 => \N__8756\,
            lcout => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNI2QAZ0Z4\,
            ltout => OPEN,
            carryin => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_5\,
            carryout => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI4TB4_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9634\,
            in2 => \_gnd_net_\,
            in3 => \N__8753\,
            lcout => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI4TBZ0Z4\,
            ltout => OPEN,
            carryin => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_6\,
            carryout => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI60D4_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9611\,
            in2 => \_gnd_net_\,
            in3 => \N__8750\,
            lcout => \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI60DZ0Z4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNIU317_4_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8743\,
            in1 => \N__8713\,
            in2 => \N__8692\,
            in3 => \N__8662\,
            lcout => \uart_inst0.tx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rTx_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011000001110100"
        )
    port map (
            in0 => \N__8579\,
            in1 => \N__8828\,
            in2 => \N__8602\,
            in3 => \N__8528\,
            lcout => \P1A7_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16914\,
            ce => 'H',
            sr => \N__16438\
        );

    \uart_inst0.uart_inst0.tx_state_RNI5LM6_0_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11565\,
            in2 => \_gnd_net_\,
            in3 => \N__11660\,
            lcout => \uart_inst0.uart_inst0.tx_state_81_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rTx_RNO_1_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__11861\,
            in1 => \N__8534\,
            in2 => \_gnd_net_\,
            in3 => \N__9988\,
            lcout => \uart_inst0.uart_inst0.rTx_6_f1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rTx_RNO_0_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101000001010"
        )
    port map (
            in0 => \N__11661\,
            in1 => \_gnd_net_\,
            in2 => \N__11582\,
            in3 => \N__11860\,
            lcout => \uart_inst0.uart_inst0.N_141_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_state_RNI9VFM2_0_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101000001010"
        )
    port map (
            in0 => \N__11648\,
            in1 => \N__9748\,
            in2 => \N__11579\,
            in3 => \N__11853\,
            lcout => \uart_inst0.uart_inst0.N_143_0\,
            ltout => \uart_inst0.uart_inst0.N_143_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_state_RNI5DQO2_0_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__14068\,
            in1 => \_gnd_net_\,
            in2 => \N__8816\,
            in3 => \_gnd_net_\,
            lcout => \uart_inst0.uart_inst0.N_143_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_bits_remaining_RNO_0_3_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__9928\,
            in1 => \N__9792\,
            in2 => \_gnd_net_\,
            in3 => \N__9956\,
            lcout => \uart_inst0.uart_inst0.un1_m3_0_a2_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_bits_remaining_RNO_0_1_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__11650\,
            in1 => \N__11855\,
            in2 => \N__11580\,
            in3 => \N__9927\,
            lcout => \uart_inst0.uart_inst0.un1_tx_bits_remaining_c1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_state_RNI9VFM2_0_0_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__11854\,
            in1 => \N__11556\,
            in2 => \N__9752\,
            in3 => \N__11649\,
            lcout => \uart_inst0.uart_inst0.N_136_0\,
            ltout => \uart_inst0.uart_inst0.N_136_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_bits_remaining_0_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9970\,
            in2 => \N__8786\,
            in3 => \N__9929\,
            lcout => \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16905\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_bits_remaining_1_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__8783\,
            in1 => \N__8775\,
            in2 => \_gnd_net_\,
            in3 => \N__9957\,
            lcout => \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16901\,
            ce => 'H',
            sr => \N__9977\
        );

    \uart_inst0.uart_inst0.tx_bits_remaining_2_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000101011010"
        )
    port map (
            in0 => \N__9902\,
            in1 => \N__9958\,
            in2 => \N__9797\,
            in3 => \N__8776\,
            lcout => \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16901\,
            ce => 'H',
            sr => \N__9977\
        );

    \uart_inst0.uart_inst0.tx_countdown_0_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100110101010"
        )
    port map (
            in0 => \N__14548\,
            in1 => \N__11875\,
            in2 => \_gnd_net_\,
            in3 => \N__10198\,
            lcout => \uart_inst0.uart_inst0.tx_countdownZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16898\,
            ce => 'H',
            sr => \N__13591\
        );

    \uart_inst0.uart_inst0.tx_countdown_1_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011000110"
        )
    port map (
            in0 => \N__10199\,
            in1 => \N__14591\,
            in2 => \N__11879\,
            in3 => \N__14549\,
            lcout => \uart_inst0.uart_inst0.tx_countdownZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16898\,
            ce => 'H',
            sr => \N__13591\
        );

    \fifo_inst.tx_fifo_inst.ram512x8_inst.RDATA_0_LC_15_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8858\,
            lcout => \wTxRdData_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVfifo_inst.tx_fifo_inst.ram512x8_inst.RDATA_0C_net\,
            ce => \N__10276\,
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_6_LC_15_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8941\,
            lcout => \fifo_inst_tx_fifo_inst_rRamRdAddr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16975\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_5_LC_15_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8965\,
            lcout => \fifo_inst_tx_fifo_inst_rRamRdAddr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16975\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_7_LC_15_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8917\,
            lcout => \fifo_inst_tx_fifo_inst_rRamRdAddr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16975\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_RNI9KL42_0_LC_15_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10214\,
            in2 => \N__10275\,
            in3 => \N__10265\,
            lcout => \rRamRdAddr_RNI9KL42_0\,
            ltout => OPEN,
            carryin => \bfn_15_3_0_\,
            carryout => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIE7TP_LC_15_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16628\,
            in1 => \N__10349\,
            in2 => \_gnd_net_\,
            in3 => \N__8834\,
            lcout => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIE7TPZ0\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_0\,
            carryout => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIGAUP_LC_15_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16631\,
            in1 => \N__12779\,
            in2 => \_gnd_net_\,
            in3 => \N__8831\,
            lcout => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIGAUPZ0\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_1\,
            carryout => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_2_c_RNIMVKN_LC_15_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10361\,
            in2 => \_gnd_net_\,
            in3 => \N__8981\,
            lcout => \un1_rRamRdAddr_cry_2_c_RNIMVKN\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_2\,
            carryout => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIKG0Q_LC_15_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16632\,
            in1 => \N__10292\,
            in2 => \_gnd_net_\,
            in3 => \N__8978\,
            lcout => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIKG0QZ0\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_3\,
            carryout => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIMJ1Q_LC_15_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16629\,
            in1 => \N__10418\,
            in2 => \_gnd_net_\,
            in3 => \N__8954\,
            lcout => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIMJ1QZ0\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_4\,
            carryout => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIOM2Q_LC_15_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16633\,
            in1 => \N__10393\,
            in2 => \_gnd_net_\,
            in3 => \N__8930\,
            lcout => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIOM2QZ0\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_5\,
            carryout => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIQP3Q_LC_15_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16630\,
            in1 => \N__10406\,
            in2 => \_gnd_net_\,
            in3 => \N__8906\,
            lcout => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIQP3QZ0\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_6\,
            carryout => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNISS4Q_LC_15_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16649\,
            in1 => \N__10333\,
            in2 => \_gnd_net_\,
            in3 => \N__8903\,
            lcout => \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNISS4QZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_1_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8890\,
            lcout => \fifo_inst_tx_fifo_inst_rRamRdAddr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16968\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rRamRdAddr_2_LC_15_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9031\,
            lcout => \fifo_inst_rx_fifo_inst_rRamRdAddr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16968\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_8_LC_15_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8869\,
            lcout => \fifo_inst_tx_fifo_inst_rRamRdAddr_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16968\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rRamRdAddr_6_LC_15_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8995\,
            lcout => \fifo_inst_rx_fifo_inst_rRamRdAddr_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16968\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m12_LC_15_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12725\,
            in2 => \_gnd_net_\,
            in3 => \N__9071\,
            lcout => \fifo_inst_rx_fifo_inst_wRamWrEn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rRamRdAddr_RNI0S8U_0_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10913\,
            in2 => \N__10954\,
            in3 => \N__10942\,
            lcout => \rRamRdAddr_RNI0S8U_0\,
            ltout => OPEN,
            carryin => \bfn_15_5_0_\,
            carryout => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIAHVB_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16660\,
            in1 => \N__10700\,
            in2 => \_gnd_net_\,
            in3 => \N__9044\,
            lcout => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIAHVBZ0\,
            ltout => OPEN,
            carryin => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_0\,
            carryout => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNICK0C_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16663\,
            in1 => \N__11044\,
            in2 => \_gnd_net_\,
            in3 => \N__9020\,
            lcout => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNICK0CZ0\,
            ltout => OPEN,
            carryin => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_1\,
            carryout => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_2_c_RNII9N9_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10712\,
            in2 => \_gnd_net_\,
            in3 => \N__9017\,
            lcout => \un1_rRamRdAddr_cry_2_c_RNII9N9\,
            ltout => OPEN,
            carryin => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_2\,
            carryout => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIGQ2C_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16664\,
            in1 => \N__11063\,
            in2 => \_gnd_net_\,
            in3 => \N__9014\,
            lcout => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIGQ2CZ0\,
            ltout => OPEN,
            carryin => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_3\,
            carryout => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIIT3C_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16661\,
            in1 => \N__11077\,
            in2 => \_gnd_net_\,
            in3 => \N__9011\,
            lcout => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIIT3CZ0\,
            ltout => OPEN,
            carryin => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_4\,
            carryout => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIK05C_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16665\,
            in1 => \N__11018\,
            in2 => \_gnd_net_\,
            in3 => \N__8984\,
            lcout => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIK05CZ0\,
            ltout => OPEN,
            carryin => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_5\,
            carryout => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIM36C_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16662\,
            in1 => \N__11032\,
            in2 => \_gnd_net_\,
            in3 => \N__9338\,
            lcout => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIM36CZ0\,
            ltout => OPEN,
            carryin => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_6\,
            carryout => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNIO67C_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__10687\,
            in1 => \N__16670\,
            in2 => \_gnd_net_\,
            in3 => \N__9335\,
            lcout => \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNIO67CZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rRamRdAddr_5_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9322\,
            lcout => \fifo_inst_rx_fifo_inst_rRamRdAddr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16954\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m10_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010110000"
        )
    port map (
            in0 => \N__10174\,
            in1 => \N__9310\,
            in2 => \N__9263\,
            in3 => \N__10526\,
            lcout => \fifo_inst_tx_fifo_inst_rDataCount_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m23_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9179\,
            in2 => \_gnd_net_\,
            in3 => \N__9155\,
            lcout => \N_101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rRamRdAddr_8_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9127\,
            lcout => \fifo_inst_rx_fifo_inst_rRamRdAddr_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16954\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rUartTxData_ess_6_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9380\,
            in1 => \N__12548\,
            in2 => \_gnd_net_\,
            in3 => \N__11230\,
            lcout => \rUartTxDataZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16948\,
            ce => \N__11179\,
            sr => \N__16414\
        );

    \rUartTxData_esr_5_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__11229\,
            in1 => \N__9386\,
            in2 => \_gnd_net_\,
            in3 => \N__12872\,
            lcout => \rUartTxDataZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16948\,
            ce => \N__11179\,
            sr => \N__16414\
        );

    \rUartTxData_esr_1_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9374\,
            in1 => \N__12536\,
            in2 => \_gnd_net_\,
            in3 => \N__11228\,
            lcout => \rUartTxDataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16948\,
            ce => \N__11179\,
            sr => \N__16414\
        );

    \rUartRxData_esr_5_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15008\,
            lcout => \rUartRxDataZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16943\,
            ce => \N__11167\,
            sr => \N__16417\
        );

    \rUartRxData_esr_7_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14894\,
            lcout => \rUartRxDataZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16943\,
            ce => \N__11167\,
            sr => \N__16417\
        );

    \rUartRxData_esr_6_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14984\,
            lcout => \rUartRxDataZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16943\,
            ce => \N__11167\,
            sr => \N__16417\
        );

    \rUartRxData_esr_2_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15551\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \rUartRxDataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16939\,
            ce => \N__11168\,
            sr => \N__16420\
        );

    \rUartRxData_esr_0_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14864\,
            lcout => \rUartRxDataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16939\,
            ce => \N__11168\,
            sr => \N__16420\
        );

    \rUartRxData_esr_3_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15536\,
            lcout => \rUartRxDataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16939\,
            ce => \N__11168\,
            sr => \N__16420\
        );

    \rUartRxData_esr_4_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15521\,
            lcout => \rUartRxDataZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16939\,
            ce => \N__11168\,
            sr => \N__16420\
        );

    \rUartRxData_esr_1_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15566\,
            lcout => \rUartRxDataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16939\,
            ce => \N__11168\,
            sr => \N__16420\
        );

    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_2_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__16676\,
            in1 => \N__9522\,
            in2 => \N__9350\,
            in3 => \N__9589\,
            lcout => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_3_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__9590\,
            in1 => \N__9349\,
            in2 => \_gnd_net_\,
            in3 => \N__9526\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16934\,
            ce => 'H',
            sr => \N__13600\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIIP78_4_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9671\,
            in1 => \N__9698\,
            in2 => \N__9644\,
            in3 => \N__9713\,
            lcout => OPEN,
            ltout => \uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIJ3HI_1_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__9392\,
            in1 => \N__11296\,
            in2 => \N__9599\,
            in3 => \N__11314\,
            lcout => \uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7\,
            ltout => \uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000100"
        )
    port map (
            in0 => \N__16677\,
            in1 => \N__9535\,
            in2 => \N__9596\,
            in3 => \N__9588\,
            lcout => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ0Z_0_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010101010"
        )
    port map (
            in0 => \N__9536\,
            in1 => \N__9849\,
            in2 => \N__9527\,
            in3 => \N__9507\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16934\,
            ce => 'H',
            sr => \N__13600\
        );

    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_5_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16680\,
            in2 => \_gnd_net_\,
            in3 => \N__9682\,
            lcout => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_6_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__16681\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9655\,
            lcout => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_7_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16682\,
            in2 => \_gnd_net_\,
            in3 => \N__9622\,
            lcout => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIGL56_8_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__9416\,
            in1 => \N__9610\,
            in2 => \_gnd_net_\,
            in3 => \N__9404\,
            lcout => \uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_3_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__16679\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9724\,
            lcout => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_4_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9725\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16927\,
            ce => 'H',
            sr => \N__13598\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_5_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15595\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16927\,
            ce => 'H',
            sr => \N__13598\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_6_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9683\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16927\,
            ce => 'H',
            sr => \N__13598\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_7_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9656\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16927\,
            ce => 'H',
            sr => \N__13598\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_8_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9623\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16927\,
            ce => 'H',
            sr => \N__13598\
        );

    \uart_inst0.uart_inst0.rx_countdown_4_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__11333\,
            in1 => \N__11752\,
            in2 => \_gnd_net_\,
            in3 => \N__11762\,
            lcout => \uart_inst0.uart_inst0.rx_countdownZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16920\,
            ce => \N__11710\,
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_countdown_2_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__11749\,
            in1 => \N__11363\,
            in2 => \N__14013\,
            in3 => \N__11693\,
            lcout => \uart_inst0.uart_inst0.rx_countdownZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16920\,
            ce => \N__11710\,
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_countdown_3_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__11342\,
            in1 => \N__11275\,
            in2 => \N__14012\,
            in3 => \N__11750\,
            lcout => \uart_inst0.uart_inst0.rx_countdownZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16920\,
            ce => \N__11710\,
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_countdown_1_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__11384\,
            in1 => \N__11151\,
            in2 => \N__14011\,
            in3 => \N__11748\,
            lcout => \uart_inst0.uart_inst0.rx_countdownZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16920\,
            ce => \N__11710\,
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_countdown_0_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__11751\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11432\,
            lcout => \uart_inst0.uart_inst0.rx_countdownZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16920\,
            ce => \N__11710\,
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_state_RNO_2_0_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11274\,
            in1 => \N__13780\,
            in2 => \N__13263\,
            in3 => \N__16034\,
            lcout => \uart_inst0.uart_inst0.rx_state_srsts_0_a5_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_state_RNI1VB3_5_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__14014\,
            in1 => \N__11273\,
            in2 => \_gnd_net_\,
            in3 => \N__11128\,
            lcout => \uart_inst0.uart_inst0.rx_countdown_2_sqmuxa_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_countdown_RNIEE7V1_5_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11331\,
            in1 => \N__11353\,
            in2 => \N__11726\,
            in3 => \N__11374\,
            lcout => \uart_inst0.uart_inst0.rx_state_srsts_0_o2_3_3\,
            ltout => \uart_inst0.uart_inst0.rx_state_srsts_0_o2_3_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_countdown_RNIFVQU2_0_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__11430\,
            in1 => \_gnd_net_\,
            in2 => \N__9803\,
            in3 => \N__11404\,
            lcout => \uart_inst0.uart_inst0.N_257_0\,
            ltout => \uart_inst0.uart_inst0.N_257_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_state_RNIJD833_1_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011111111"
        )
    port map (
            in0 => \N__13250\,
            in1 => \N__16033\,
            in2 => \N__9800\,
            in3 => \N__11455\,
            lcout => \uart_inst0.uart_inst0.N_252_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_bits_remaining_RNIMJMP_3_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9796\,
            in1 => \N__9959\,
            in2 => \N__9773\,
            in3 => \N__9925\,
            lcout => \uart_inst0.uart_inst0.N_157\,
            ltout => \uart_inst0.uart_inst0.N_157_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_state_RNIR8D01_0_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11552\,
            in2 => \N__9740\,
            in3 => \N__11659\,
            lcout => \uart_inst0.uart_inst0.tx_state_1_sqmuxa_1_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_countdown_RNIEM2M1_0_2_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13630\,
            in1 => \N__14592\,
            in2 => \N__13684\,
            in3 => \N__14550\,
            lcout => \uart_inst0.uart_inst0.N_147_0\,
            ltout => \uart_inst0.uart_inst0.N_147_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_state_1_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010001000"
        )
    port map (
            in0 => \N__14004\,
            in1 => \N__11575\,
            in2 => \N__9890\,
            in3 => \N__11658\,
            lcout => \uart_inst0.uart_inst0.tx_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16911\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_state_RNO_0_1_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110011"
        )
    port map (
            in0 => \N__13317\,
            in1 => \N__13254\,
            in2 => \_gnd_net_\,
            in3 => \N__11129\,
            lcout => OPEN,
            ltout => \uart_inst0.uart_inst0.N_277_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_state_1_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001100"
        )
    port map (
            in0 => \N__11130\,
            in1 => \N__14023\,
            in2 => \N__9887\,
            in3 => \N__13823\,
            lcout => \uart_inst0.uart_inst0.rx_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16911\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_state_4_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011000000"
        )
    port map (
            in0 => \N__13824\,
            in1 => \N__14003\,
            in2 => \N__11282\,
            in3 => \N__9875\,
            lcout => \uart_inst0.uart_inst0.rx_stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16911\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_state_RNO_1_0_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__11691\,
            in1 => \N__9874\,
            in2 => \N__13787\,
            in3 => \N__13822\,
            lcout => OPEN,
            ltout => \uart_inst0.uart_inst0.N_280_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_state_0_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111111101"
        )
    port map (
            in0 => \N__14022\,
            in1 => \N__9884\,
            in2 => \N__9878\,
            in3 => \N__9860\,
            lcout => \uart_inst0.uart_inst0.rx_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16911\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_state_RNO_0_0_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__11482\,
            in1 => \N__13316\,
            in2 => \_gnd_net_\,
            in3 => \N__9873\,
            lcout => \uart_inst0.uart_inst0.N_261_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_countdown_RNIEM2M1_2_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13634\,
            in1 => \N__14590\,
            in2 => \N__13679\,
            in3 => \N__14543\,
            lcout => \uart_inst0.uart_inst0.N_147_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_state_RNO_0_0_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111011010"
        )
    port map (
            in0 => \N__11654\,
            in1 => \N__11858\,
            in2 => \N__11581\,
            in3 => \N__9854\,
            lcout => OPEN,
            ltout => \uart_inst0.uart_inst0.tx_state_ns_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_state_0_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110000001100"
        )
    port map (
            in0 => \N__11859\,
            in1 => \N__13999\,
            in2 => \N__9995\,
            in3 => \N__9992\,
            lcout => \uart_inst0.uart_inst0.tx_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16906\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_state_RNI1319_0_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100001111"
        )
    port map (
            in0 => \N__11560\,
            in1 => \_gnd_net_\,
            in2 => \N__14021\,
            in3 => \N__11651\,
            lcout => \uart_inst0.uart_inst0.tx_state_RNI1319Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_bits_remaining_RNO_1_2_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9955\,
            in2 => \_gnd_net_\,
            in3 => \N__9926\,
            lcout => OPEN,
            ltout => \uart_inst0.uart_inst0.un1_tx_bits_remaining_ac0_1_a0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_bits_remaining_RNO_0_2_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__11561\,
            in1 => \N__11857\,
            in2 => \N__9905\,
            in3 => \N__11652\,
            lcout => \uart_inst0.uart_inst0.un1_tx_bits_remaining_ac0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_countdown_RNIEGNA5_2_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100110011"
        )
    port map (
            in0 => \N__11856\,
            in1 => \N__13998\,
            in2 => \_gnd_net_\,
            in3 => \N__10196\,
            lcout => \uart_inst0.uart_inst0.un1_rx_state49_i\,
            ltout => \uart_inst0.uart_inst0.un1_rx_state49_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_clk_divider_esr_RNO_0_14_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9896\,
            in3 => \N__13510\,
            lcout => \uart_inst0.uart_inst0.N_147_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_countdown_RNO_0_3_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__14547\,
            in1 => \N__11501\,
            in2 => \N__13680\,
            in3 => \N__10197\,
            lcout => OPEN,
            ltout => \uart_inst0.uart_inst0.tx_countdown_RNO_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_countdown_3_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001110000"
        )
    port map (
            in0 => \N__11873\,
            in1 => \N__11587\,
            in2 => \N__9893\,
            in3 => \N__11665\,
            lcout => \uart_inst0.uart_inst0.tx_countdownZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16902\,
            ce => 'H',
            sr => \N__13592\
        );

    \uart_inst0.uart_inst0.tx_clk_divider_esr_RNIIIJI_14_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__11955\,
            in1 => \N__11988\,
            in2 => \_gnd_net_\,
            in3 => \N__12115\,
            lcout => \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_11_3\,
            ltout => \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_11_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_clk_divider_esr_RNI4CAI3_14_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14381\,
            in1 => \N__14470\,
            in2 => \N__10202\,
            in3 => \N__14500\,
            lcout => \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_clk_divider_RNIQUQ11_4_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12045\,
            in1 => \N__12018\,
            in2 => \N__12077\,
            in3 => \N__11787\,
            lcout => \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_clk_divider_RNIEC1S_10_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12502\,
            in1 => \N__11901\,
            in2 => \N__12148\,
            in3 => \N__11925\,
            lcout => \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_11_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_clk_divider_10_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001100110"
        )
    port map (
            in0 => \N__11926\,
            in1 => \N__13549\,
            in2 => \_gnd_net_\,
            in3 => \N__11912\,
            lcout => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16899\,
            ce => 'H',
            sr => \N__14636\
        );

    \uart_inst0.uart_inst0.tx_clk_divider_11_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100100010"
        )
    port map (
            in0 => \N__13550\,
            in1 => \N__11888\,
            in2 => \_gnd_net_\,
            in3 => \N__11902\,
            lcout => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16899\,
            ce => 'H',
            sr => \N__14636\
        );

    \uart_inst0.uart_inst0.tx_clk_divider_13_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001011010"
        )
    port map (
            in0 => \N__12144\,
            in1 => \_gnd_net_\,
            in2 => \N__13556\,
            in3 => \N__12128\,
            lcout => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16899\,
            ce => 'H',
            sr => \N__14636\
        );

    \uart_inst0.uart_inst0.tx_clk_divider_5_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101110100100010"
        )
    port map (
            in0 => \N__13554\,
            in1 => \N__12056\,
            in2 => \_gnd_net_\,
            in3 => \N__12076\,
            lcout => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16899\,
            ce => 'H',
            sr => \N__14636\
        );

    \uart_inst0.uart_inst0.tx_clk_divider_6_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101110100100010"
        )
    port map (
            in0 => \N__13555\,
            in1 => \N__12029\,
            in2 => \_gnd_net_\,
            in3 => \N__12047\,
            lcout => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16899\,
            ce => 'H',
            sr => \N__14636\
        );

    \rTxData_0_LC_16_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__14020\,
            in1 => \N__10102\,
            in2 => \_gnd_net_\,
            in3 => \N__10173\,
            lcout => \rTxDataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16981\,
            ce => 'H',
            sr => \N__16357\
        );

    \fifo_inst.ft2232h_inst.rTxBusReady_esr_LC_16_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__10607\,
            in1 => \N__10652\,
            in2 => \_gnd_net_\,
            in3 => \N__10532\,
            lcout => \rTxBusReady\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16978\,
            ce => \N__10469\,
            sr => \N__16359\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_3_LC_16_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000010110000"
        )
    port map (
            in0 => \N__10226\,
            in1 => \N__16645\,
            in2 => \N__10445\,
            in3 => \N__10280\,
            lcout => \fifo_inst_tx_fifo_inst_rRamRdAddr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16976\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m74_LC_16_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011100000000"
        )
    port map (
            in0 => \N__10278\,
            in1 => \N__10224\,
            in2 => \N__16698\,
            in3 => \N__10441\,
            lcout => m74,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m72_e_5_LC_16_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10417\,
            in1 => \N__10291\,
            in2 => \N__16697\,
            in3 => \N__12775\,
            lcout => OPEN,
            ltout => \uart_inst0.tx_uart_fifo_inst.m72_eZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m72_e_LC_16_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__10405\,
            in1 => \N__10394\,
            in2 => \N__10382\,
            in3 => \N__10319\,
            lcout => \uart_inst0.tx_uart_fifo_inst.N_100\,
            ltout => \uart_inst0.tx_uart_fifo_inst.N_100_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m73_LC_16_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011000100"
        )
    port map (
            in0 => \N__16644\,
            in1 => \N__10234\,
            in2 => \N__10379\,
            in3 => \N__10277\,
            lcout => m73,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m72_e_6_LC_16_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__10360\,
            in1 => \N__10348\,
            in2 => \N__10337\,
            in3 => \N__10213\,
            lcout => \uart_inst0.tx_uart_fifo_inst.m72_eZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_4_LC_16_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10303\,
            lcout => \fifo_inst_tx_fifo_inst_rRamRdAddr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16976\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_0_LC_16_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000000110000"
        )
    port map (
            in0 => \N__10279\,
            in1 => \N__16640\,
            in2 => \N__10238\,
            in3 => \N__10225\,
            lcout => \fifo_inst_tx_fifo_inst_rRamRdAddr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16976\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rRamRdAddr_7_LC_16_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10792\,
            lcout => \fifo_inst_rx_fifo_inst_rRamRdAddr_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16973\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rRamRdAddr_3_LC_16_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010010001100"
        )
    port map (
            in0 => \N__10994\,
            in1 => \N__10757\,
            in2 => \N__16699\,
            in3 => \N__10966\,
            lcout => \fifo_inst_rx_fifo_inst_rRamRdAddr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16973\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rRamRdAddr_1_LC_16_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10768\,
            lcout => \fifo_inst_rx_fifo_inst_rRamRdAddr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16973\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m60_LC_16_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100000000"
        )
    port map (
            in0 => \N__16653\,
            in1 => \N__10993\,
            in2 => \N__10967\,
            in3 => \N__10756\,
            lcout => m60,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rRamRdAddr_4_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10723\,
            lcout => \fifo_inst_rx_fifo_inst_rRamRdAddr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16969\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m58_e_6_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__10711\,
            in1 => \N__10699\,
            in2 => \N__10688\,
            in3 => \N__10912\,
            lcout => \uart_inst0.tx_uart_fifo_inst.m58_eZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.un1_rFifoState_1_sqmuxa_0_i_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101110"
        )
    port map (
            in0 => \N__10673\,
            in1 => \N__10657\,
            in2 => \N__10593\,
            in3 => \N__10531\,
            lcout => OPEN,
            ltout => \fifo_inst_ft2232h_inst_un1_rFifoState_1_sqmuxa_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ft2232h_inst.rTxBusReady_esr_RNO_LC_16_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10472\,
            in3 => \N__14100\,
            lcout => \fifo_inst.ft2232h_inst.un1_rFifoState_1_sqmuxa_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m59_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010010001100"
        )
    port map (
            in0 => \N__10992\,
            in1 => \N__10975\,
            in2 => \N__16701\,
            in3 => \N__10961\,
            lcout => m59,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m58_e_5_LC_16_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11078\,
            in1 => \N__11062\,
            in2 => \N__16702\,
            in3 => \N__11051\,
            lcout => OPEN,
            ltout => \uart_inst0.tx_uart_fifo_inst.m58_eZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m58_e_LC_16_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__11033\,
            in1 => \N__11017\,
            in2 => \N__11003\,
            in3 => \N__11000\,
            lcout => \uart_inst0.tx_uart_fifo_inst.N_99\,
            ltout => \uart_inst0.tx_uart_fifo_inst.N_99_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rRamRdAddr_0_LC_16_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000101010"
        )
    port map (
            in0 => \N__10976\,
            in1 => \N__10962\,
            in2 => \N__10916\,
            in3 => \N__16666\,
            lcout => \fifo_inst_rx_fifo_inst_rRamRdAddr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16969\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rRxData_4_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14774\,
            lcout => \rRxDataZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16961\,
            ce => \N__12850\,
            sr => \_gnd_net_\
        );

    \rUartTxData_esr_3_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10901\,
            in1 => \N__12512\,
            in2 => \_gnd_net_\,
            in3 => \N__11244\,
            lcout => \rUartTxDataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16955\,
            ce => \N__11183\,
            sr => \N__16418\
        );

    \rUartTxData_esr_4_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__11245\,
            in1 => \_gnd_net_\,
            in2 => \N__10877\,
            in3 => \N__10865\,
            lcout => \rUartTxDataZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16955\,
            ce => \N__11183\,
            sr => \N__16418\
        );

    \rUartTxData_esr_7_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__12860\,
            in1 => \_gnd_net_\,
            in2 => \N__10847\,
            in3 => \N__11246\,
            lcout => \rUartTxDataZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16955\,
            ce => \N__11183\,
            sr => \N__16418\
        );

    \rUartTxData_esr_2_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__11243\,
            in1 => \_gnd_net_\,
            in2 => \N__12524\,
            in3 => \N__10826\,
            lcout => \rUartTxDataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16955\,
            ce => \N__11183\,
            sr => \N__16418\
        );

    \rUartTxData_esr_0_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__12881\,
            in1 => \N__11255\,
            in2 => \_gnd_net_\,
            in3 => \N__11242\,
            lcout => \rUartTxDataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16955\,
            ce => \N__11183\,
            sr => \N__16418\
        );

    \rUartRxState_RNITBQ5_0_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16675\,
            in2 => \_gnd_net_\,
            in3 => \N__13040\,
            lcout => \rUartRxState_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.rDataCount_RNO_0_1_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__13140\,
            in1 => \N__13093\,
            in2 => \_gnd_net_\,
            in3 => \N__14949\,
            lcout => \uart_inst0.rx_uart_fifo_inst.un1_rDataCount15_2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.rDataCount_RNIG8UP_3_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11103\,
            in2 => \_gnd_net_\,
            in3 => \N__12929\,
            lcout => \uart_inst0.rx_uart_fifo_inst.wRamWrEn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rRxWrEn_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011110100"
        )
    port map (
            in0 => \N__12930\,
            in1 => \N__11483\,
            in2 => \N__11108\,
            in3 => \N__11156\,
            lcout => \uart_inst0.wRxWrEn_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16944\,
            ce => 'H',
            sr => \N__16425\
        );

    \uart_inst0.rx_uart_fifo_inst.rDataCount_RNO_0_3_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011100011111"
        )
    port map (
            in0 => \N__13002\,
            in1 => \N__13094\,
            in2 => \N__14962\,
            in3 => \N__11104\,
            lcout => \uart_inst0.rx_uart_fifo_inst.un1_rDataCount_axbxc3_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_0_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16678\,
            in2 => \_gnd_net_\,
            in3 => \N__13216\,
            lcout => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_1_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13217\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16935\,
            ce => 'H',
            sr => \N__13601\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_2_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15710\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16935\,
            ce => 'H',
            sr => \N__13601\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_4_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15491\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16935\,
            ce => 'H',
            sr => \N__13601\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_5_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15446\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16935\,
            ce => 'H',
            sr => \N__13601\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_6_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15512\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16935\,
            ce => 'H',
            sr => \N__13601\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_7_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15731\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16935\,
            ce => 'H',
            sr => \N__13601\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ0Z_1_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13484\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16935\,
            ce => 'H',
            sr => \N__13601\
        );

    \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_2_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15623\,
            lcout => \uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16935\,
            ce => 'H',
            sr => \N__13601\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_8_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15689\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16931\,
            ce => 'H',
            sr => \N__13599\
        );

    \uart_inst0.uart_inst0.rRxData_7_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13290\,
            in1 => \N__16137\,
            in2 => \_gnd_net_\,
            in3 => \N__14036\,
            lcout => \uart_inst0.wRxWrData_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16928\,
            ce => 'H',
            sr => \N__16449\
        );

    \uart_inst0.uart_inst0.rx_state_5_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000000000"
        )
    port map (
            in0 => \N__13779\,
            in1 => \N__13259\,
            in2 => \N__13319\,
            in3 => \N__15937\,
            lcout => \uart_inst0.uart_inst0.rx_stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16925\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_countdown_RNIBD513_0_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__11402\,
            in1 => \N__11428\,
            in2 => \N__13986\,
            in3 => \N__11464\,
            lcout => \uart_inst0.uart_inst0.N_283\,
            ltout => \uart_inst0.uart_inst0.N_283_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_state_6_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000010000000"
        )
    port map (
            in0 => \N__13315\,
            in1 => \N__13778\,
            in2 => \N__11486\,
            in3 => \_gnd_net_\,
            lcout => \uart_inst0.uart_inst0.rx_stateZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16925\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_countdown_RNIHNBV2_0_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__11403\,
            in1 => \N__11429\,
            in2 => \N__16044\,
            in3 => \N__11465\,
            lcout => \uart_inst0.uart_inst0.rRxData_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_state_RNI3F11_1_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16032\,
            in2 => \_gnd_net_\,
            in3 => \N__13258\,
            lcout => \uart_inst0.uart_inst0.N_258_0\,
            ltout => \uart_inst0.uart_inst0.N_258_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_state_RNIGVTK5_5_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111011101"
        )
    port map (
            in0 => \N__11456\,
            in1 => \N__11444\,
            in2 => \N__11435\,
            in3 => \N__13825\,
            lcout => \uart_inst0.uart_inst0.rx_countdowne_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_countdown_cry_c_0_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11431\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_15_0_\,
            carryout => \uart_inst0.uart_inst0.rx_countdown_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_countdown_RNO_0_1_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11405\,
            in2 => \N__12405\,
            in3 => \N__11378\,
            lcout => \uart_inst0.uart_inst0.rx_countdown_s_1\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.rx_countdown_cry_0\,
            carryout => \uart_inst0.uart_inst0.rx_countdown_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_countdown_RNO_0_2_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11375\,
            in2 => \N__12407\,
            in3 => \N__11357\,
            lcout => \uart_inst0.uart_inst0.rx_countdown_s_2\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.rx_countdown_cry_1\,
            carryout => \uart_inst0.uart_inst0.rx_countdown_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_countdown_RNO_0_3_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11354\,
            in2 => \N__12406\,
            in3 => \N__11336\,
            lcout => \uart_inst0.uart_inst0.rx_countdown_s_3\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.rx_countdown_cry_2\,
            carryout => \uart_inst0.uart_inst0.rx_countdown_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_countdown_cry_3_THRU_LUT4_0_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11332\,
            in2 => \N__12408\,
            in3 => \N__11756\,
            lcout => \uart_inst0.uart_inst0.rx_countdown_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.rx_countdown_cry_3\,
            carryout => \uart_inst0.uart_inst0.rx_countdown_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_countdown_5_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__11753\,
            in1 => \N__11725\,
            in2 => \_gnd_net_\,
            in3 => \N__11729\,
            lcout => \uart_inst0.uart_inst0.rx_countdownZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16921\,
            ce => \N__11711\,
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_state_RNO_1_2_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__13724\,
            in1 => \N__13739\,
            in2 => \N__13264\,
            in3 => \N__13818\,
            lcout => OPEN,
            ltout => \uart_inst0.uart_inst0.N_276_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_state_2_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__14005\,
            in1 => \N__11692\,
            in2 => \N__11672\,
            in3 => \N__11492\,
            lcout => \uart_inst0.uart_inst0.rx_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16915\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_countdown_RNO_0_2_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__14600\,
            in1 => \N__11653\,
            in2 => \N__11583\,
            in3 => \N__14555\,
            lcout => \uart_inst0.uart_inst0.tx_N_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_countdown_RNO_1_3_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__13628\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14599\,
            lcout => \uart_inst0.uart_inst0.un1_m3_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_state_RNO_0_2_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110011"
        )
    port map (
            in0 => \N__13318\,
            in1 => \N__16022\,
            in2 => \_gnd_net_\,
            in3 => \N__13817\,
            lcout => \uart_inst0.uart_inst0.N_275\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_clk_divider_7_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100110101010"
        )
    port map (
            in0 => \N__12020\,
            in1 => \N__12002\,
            in2 => \_gnd_net_\,
            in3 => \N__13545\,
            lcout => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16912\,
            ce => 'H',
            sr => \N__14635\
        );

    \uart_inst0.uart_inst0.tx_clk_divider_8_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100100010"
        )
    port map (
            in0 => \N__13546\,
            in1 => \N__11972\,
            in2 => \_gnd_net_\,
            in3 => \N__11992\,
            lcout => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16912\,
            ce => 'H',
            sr => \N__14635\
        );

    \uart_inst0.uart_inst0.tx_clk_divider_9_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100110101010"
        )
    port map (
            in0 => \N__11959\,
            in1 => \N__11939\,
            in2 => \_gnd_net_\,
            in3 => \N__13547\,
            lcout => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16912\,
            ce => 'H',
            sr => \N__14635\
        );

    \uart_inst0.uart_inst0.tx_clk_divider_12_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100100010"
        )
    port map (
            in0 => \N__13541\,
            in1 => \N__12482\,
            in2 => \_gnd_net_\,
            in3 => \N__12501\,
            lcout => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16912\,
            ce => 'H',
            sr => \N__14635\
        );

    \uart_inst0.uart_inst0.tx_clk_divider_4_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101101000100"
        )
    port map (
            in0 => \N__11771\,
            in1 => \N__13544\,
            in2 => \_gnd_net_\,
            in3 => \N__11789\,
            lcout => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16912\,
            ce => 'H',
            sr => \N__14635\
        );

    \uart_inst0.uart_inst0.tx_clk_divider_1_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010100001010"
        )
    port map (
            in0 => \N__13542\,
            in1 => \_gnd_net_\,
            in2 => \N__11813\,
            in3 => \N__14399\,
            lcout => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16912\,
            ce => 'H',
            sr => \N__14635\
        );

    \uart_inst0.uart_inst0.tx_clk_divider_2_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110100100010"
        )
    port map (
            in0 => \N__13543\,
            in1 => \N__11801\,
            in2 => \_gnd_net_\,
            in3 => \N__14450\,
            lcout => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16912\,
            ce => 'H',
            sr => \N__14635\
        );

    \uart_inst0.uart_inst0.tx_clk_divider_0_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100110011001"
        )
    port map (
            in0 => \N__11874\,
            in1 => \N__14432\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_16_18_0_\,
            carryout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_0_s1\,
            clk => \N__16907\,
            ce => 'H',
            sr => \N__14642\
        );

    \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_0_s1_THRU_LUT4_0_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14398\,
            in2 => \N__12449\,
            in3 => \N__11804\,
            lcout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_0_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_0_s1\,
            carryout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_1_s1_THRU_LUT4_0_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14449\,
            in2 => \N__12453\,
            in3 => \N__11795\,
            lcout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_1_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_1_s1\,
            carryout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_2_s1_THRU_LUT4_0_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14418\,
            in2 => \N__12450\,
            in3 => \N__11792\,
            lcout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_2_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_2_s1\,
            carryout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_3_s1_THRU_LUT4_0_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11788\,
            in2 => \N__12454\,
            in3 => \N__11765\,
            lcout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_3_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_3_s1\,
            carryout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_4_s1_THRU_LUT4_0_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12075\,
            in2 => \N__12451\,
            in3 => \N__12050\,
            lcout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_4_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_4_s1\,
            carryout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_5_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_5_s1_THRU_LUT4_0_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12046\,
            in2 => \N__12455\,
            in3 => \N__12023\,
            lcout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_5_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_5_s1\,
            carryout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_6_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_6_s1_THRU_LUT4_0_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12019\,
            in2 => \N__12452\,
            in3 => \N__11996\,
            lcout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_6_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_6_s1\,
            carryout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_7_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_7_s1_THRU_LUT4_0_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11993\,
            in2 => \N__12459\,
            in3 => \N__11963\,
            lcout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_7_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_16_19_0_\,
            carryout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_8_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_8_s1_THRU_LUT4_0_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11960\,
            in2 => \N__12457\,
            in3 => \N__11930\,
            lcout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_8_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_8_s1\,
            carryout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_9_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_9_s1_THRU_LUT4_0_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11927\,
            in2 => \N__12460\,
            in3 => \N__11906\,
            lcout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_9_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_9_s1\,
            carryout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_10_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_10_s1_THRU_LUT4_0_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11903\,
            in2 => \N__12456\,
            in3 => \N__11882\,
            lcout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_10_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_10_s1\,
            carryout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_11_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_11_s1_THRU_LUT4_0_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12503\,
            in2 => \N__12458\,
            in3 => \N__12473\,
            lcout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_11_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_11_s1\,
            carryout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_12_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_12_s1_THRU_LUT4_0_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12439\,
            in2 => \N__12149\,
            in3 => \N__12122\,
            lcout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_12_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_12_s1\,
            carryout => \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_13_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_clk_divider_esr_14_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12116\,
            in2 => \_gnd_net_\,
            in3 => \N__12119\,
            lcout => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16903\,
            ce => \N__12104\,
            sr => \N__14637\
        );

    \fifo_inst.rx_fifo_inst.rRamWrAddr_RNI9D19_0_LC_17_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14797\,
            in2 => \N__14843\,
            in3 => \N__14840\,
            lcout => \rRamWrAddr_RNI9D19_0\,
            ltout => OPEN,
            carryin => \bfn_17_2_0_\,
            carryout => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rRamWrAddr_1_LC_17_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16634\,
            in1 => \N__14155\,
            in2 => \_gnd_net_\,
            in3 => \N__12092\,
            lcout => \fifo_inst_rx_fifo_inst_rRamWrAddr_1\,
            ltout => OPEN,
            carryin => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_0\,
            carryout => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_1\,
            clk => \N__16982\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rRamWrAddr_2_LC_17_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16637\,
            in1 => \N__14274\,
            in2 => \_gnd_net_\,
            in3 => \N__12089\,
            lcout => \fifo_inst_rx_fifo_inst_rRamWrAddr_2\,
            ltout => OPEN,
            carryin => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_1\,
            carryout => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_2\,
            clk => \N__16982\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_2_c_RNIOTMG_LC_17_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14182\,
            in2 => \_gnd_net_\,
            in3 => \N__12086\,
            lcout => \un1_rRamWrAddr_cry_2_c_RNIOTMG\,
            ltout => OPEN,
            carryin => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_2\,
            carryout => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rRamWrAddr_4_LC_17_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16638\,
            in1 => \N__14308\,
            in2 => \_gnd_net_\,
            in3 => \N__12083\,
            lcout => \fifo_inst_rx_fifo_inst_rRamWrAddr_4\,
            ltout => OPEN,
            carryin => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_3\,
            carryout => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_4\,
            clk => \N__16982\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rRamWrAddr_5_LC_17_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16635\,
            in1 => \N__14332\,
            in2 => \_gnd_net_\,
            in3 => \N__12080\,
            lcout => \fifo_inst_rx_fifo_inst_rRamWrAddr_5\,
            ltout => OPEN,
            carryin => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_4\,
            carryout => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_5\,
            clk => \N__16982\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rRamWrAddr_6_LC_17_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16639\,
            in1 => \N__14218\,
            in2 => \_gnd_net_\,
            in3 => \N__12812\,
            lcout => \fifo_inst_rx_fifo_inst_rRamWrAddr_6\,
            ltout => OPEN,
            carryin => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_5\,
            carryout => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_6\,
            clk => \N__16982\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rRamWrAddr_7_LC_17_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16636\,
            in1 => \N__14248\,
            in2 => \_gnd_net_\,
            in3 => \N__12809\,
            lcout => \fifo_inst_rx_fifo_inst_rRamWrAddr_7\,
            ltout => OPEN,
            carryin => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_6\,
            carryout => \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_7\,
            clk => \N__16982\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rRamWrAddr_8_LC_17_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__16659\,
            in1 => \N__14130\,
            in2 => \_gnd_net_\,
            in3 => \N__12806\,
            lcout => \fifo_inst_rx_fifo_inst_rRamWrAddr_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16979\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_2_LC_17_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12796\,
            lcout => \fifo_inst_tx_fifo_inst_rRamRdAddr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16979\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.N_84_mux_i_LC_17_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12763\,
            in1 => \N__12695\,
            in2 => \N__12656\,
            in3 => \N__12599\,
            lcout => \N_84_mux_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rRxData_6_LC_17_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14653\,
            lcout => \rRxDataZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16974\,
            ce => \N__12851\,
            sr => \_gnd_net_\
        );

    \rRxData_1_LC_17_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14689\,
            lcout => \rRxDataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16974\,
            ce => \N__12851\,
            sr => \_gnd_net_\
        );

    \rRxData_2_LC_17_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14671\,
            lcout => \rRxDataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16974\,
            ce => \N__12851\,
            sr => \_gnd_net_\
        );

    \rRxData_3_LC_17_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14750\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \rRxDataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16974\,
            ce => \N__12851\,
            sr => \_gnd_net_\
        );

    \rRxData_0_LC_17_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15319\,
            lcout => \rRxDataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16974\,
            ce => \N__12851\,
            sr => \_gnd_net_\
        );

    \rRxData_5_LC_17_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14710\,
            lcout => \rRxDataZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16974\,
            ce => \N__12851\,
            sr => \_gnd_net_\
        );

    \rRxData_7_LC_17_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14728\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \rRxDataZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16974\,
            ce => \N__12851\,
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNO_0_0_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15168\,
            in2 => \N__13157\,
            in3 => \N__13154\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNO_0_0_0\,
            ltout => OPEN,
            carryin => \bfn_17_6_0_\,
            carryout => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_1_LC_17_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15198\,
            in2 => \_gnd_net_\,
            in3 => \N__12827\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_1\,
            ltout => OPEN,
            carryin => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_0\,
            carryout => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_1\,
            clk => \N__16970\,
            ce => 'H',
            sr => \N__13604\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_2_LC_17_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15225\,
            in2 => \_gnd_net_\,
            in3 => \N__12824\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_2\,
            ltout => OPEN,
            carryin => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_1\,
            carryout => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_2\,
            clk => \N__16970\,
            ce => 'H',
            sr => \N__13604\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNO_0_3_LC_17_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15253\,
            in2 => \_gnd_net_\,
            in3 => \N__12821\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNO_0_0_3\,
            ltout => OPEN,
            carryin => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_2\,
            carryout => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_4_LC_17_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15042\,
            in2 => \_gnd_net_\,
            in3 => \N__12818\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_4\,
            ltout => OPEN,
            carryin => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_3\,
            carryout => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_4\,
            clk => \N__16970\,
            ce => 'H',
            sr => \N__13604\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_5_LC_17_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15099\,
            in2 => \_gnd_net_\,
            in3 => \N__12815\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_5\,
            ltout => OPEN,
            carryin => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_4\,
            carryout => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_5\,
            clk => \N__16970\,
            ce => 'H',
            sr => \N__13604\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_6_LC_17_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15126\,
            in2 => \_gnd_net_\,
            in3 => \N__12905\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_6\,
            ltout => OPEN,
            carryin => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_5\,
            carryout => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_6\,
            clk => \N__16970\,
            ce => 'H',
            sr => \N__13604\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_7_LC_17_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15072\,
            in2 => \_gnd_net_\,
            in3 => \N__12902\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_7\,
            ltout => OPEN,
            carryin => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_6\,
            carryout => \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_7\,
            clk => \N__16970\,
            ce => 'H',
            sr => \N__13604\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_8_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15286\,
            in2 => \_gnd_net_\,
            in3 => \N__12899\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16962\,
            ce => 'H',
            sr => \N__13603\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_3_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__13146\,
            in1 => \N__15025\,
            in2 => \N__15152\,
            in3 => \N__12896\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16962\,
            ce => 'H',
            sr => \N__13603\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_0_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__15148\,
            in1 => \N__12890\,
            in2 => \N__15026\,
            in3 => \N__13147\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16962\,
            ce => 'H',
            sr => \N__13603\
        );

    \rUartRxState_0_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__14024\,
            in1 => \N__13041\,
            in2 => \_gnd_net_\,
            in3 => \N__13372\,
            lcout => \rUartRxStateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16956\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.rDataCount_RNO_0_2_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100011100000"
        )
    port map (
            in0 => \N__12966\,
            in1 => \N__13092\,
            in2 => \N__14961\,
            in3 => \N__13142\,
            lcout => \uart_inst0.rx_uart_fifo_inst.un1_rDataCount_c2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.rDataCount_RNI2JT81_0_2_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13091\,
            in1 => \N__12934\,
            in2 => \N__12968\,
            in3 => \N__13001\,
            lcout => \wUartRxEmpty\,
            ltout => \wUartRxEmpty_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.rDataCount_RNITL9D2_2_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13141\,
            in2 => \N__12884\,
            in3 => \N__14950\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rDataCount_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.rDataCount_RNI2JT81_2_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13000\,
            in1 => \N__12962\,
            in2 => \N__12935\,
            in3 => \N__13090\,
            lcout => \uart_inst0.rx_uart_fifo_inst.wUartRxEmpty_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.rDataCount_0_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100101110110100"
        )
    port map (
            in0 => \N__13371\,
            in1 => \N__14960\,
            in2 => \N__13156\,
            in3 => \N__13089\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16949\,
            ce => 'H',
            sr => \N__16429\
        );

    \uart_inst0.rx_uart_fifo_inst.rDataCount_RNI3V391_2_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__13088\,
            in1 => \N__14943\,
            in2 => \N__13003\,
            in3 => \N__12957\,
            lcout => OPEN,
            ltout => \uart_inst0.rx_uart_fifo_inst.rDataCount_RNI3V391Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.rDataCount_RNIO7PT1_3_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__14944\,
            in1 => \_gnd_net_\,
            in2 => \N__13061\,
            in3 => \N__12927\,
            lcout => \uart_inst0.rx_uart_fifo_inst.wRamRdEn\,
            ltout => \uart_inst0.rx_uart_fifo_inst.wRamRdEn_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.rDataCount_1_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100101000110"
        )
    port map (
            in0 => \N__13058\,
            in1 => \N__13012\,
            in2 => \N__13052\,
            in3 => \N__12958\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16949\,
            ce => 'H',
            sr => \N__16429\
        );

    \rUartRxEn_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__13370\,
            in1 => \N__13042\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \rUartRxEnZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16949\,
            ce => 'H',
            sr => \N__16429\
        );

    \uart_inst0.rx_uart_fifo_inst.rDataCount_2_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001011010010110"
        )
    port map (
            in0 => \N__13019\,
            in1 => \N__13013\,
            in2 => \N__13004\,
            in3 => \_gnd_net_\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16949\,
            ce => 'H',
            sr => \N__16429\
        );

    \uart_inst0.rx_uart_fifo_inst.rDataCount_3_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100010000"
        )
    port map (
            in0 => \N__14945\,
            in1 => \N__12974\,
            in2 => \N__12967\,
            in3 => \N__12928\,
            lcout => \uart_inst0.wRxWrFull_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16949\,
            ce => 'H',
            sr => \N__16429\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNID4JC2_0_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13352\,
            in2 => \N__15798\,
            in3 => \N__15790\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNID4JC2Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIK0HS_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13180\,
            in2 => \_gnd_net_\,
            in3 => \N__13205\,
            lcout => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIK0HSZ0\,
            ltout => OPEN,
            carryin => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_0\,
            carryout => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIM3IS_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13168\,
            in2 => \_gnd_net_\,
            in3 => \N__13202\,
            lcout => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIM3ISZ0\,
            ltout => OPEN,
            carryin => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_1\,
            carryout => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNIO6JS_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13337\,
            in3 => \N__13199\,
            lcout => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNIO6JSZ0\,
            ltout => OPEN,
            carryin => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_2\,
            carryout => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIQ9KS_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13414\,
            in2 => \_gnd_net_\,
            in3 => \N__13196\,
            lcout => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIQ9KSZ0\,
            ltout => OPEN,
            carryin => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_3\,
            carryout => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNISCLS_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13441\,
            in2 => \_gnd_net_\,
            in3 => \N__13193\,
            lcout => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNISCLSZ0\,
            ltout => OPEN,
            carryin => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_4\,
            carryout => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIUFMS_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13457\,
            in3 => \N__13190\,
            lcout => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIUFMSZ0\,
            ltout => OPEN,
            carryin => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_5\,
            carryout => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI0JNS_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13426\,
            in2 => \_gnd_net_\,
            in3 => \N__13187\,
            lcout => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI0JNSZ0\,
            ltout => OPEN,
            carryin => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_6\,
            carryout => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI2MOS_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13394\,
            in2 => \_gnd_net_\,
            in3 => \N__13184\,
            lcout => \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI2MOSZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNI17A54_1_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__13385\,
            in1 => \N__13181\,
            in2 => \N__13403\,
            in3 => \N__13169\,
            lcout => \uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_0_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16693\,
            in2 => \_gnd_net_\,
            in3 => \N__13483\,
            lcout => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNIA98R1_4_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13456\,
            in1 => \N__13442\,
            in2 => \N__13430\,
            in3 => \N__13415\,
            lcout => \uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNIA1EC1_8_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__13393\,
            in1 => \N__13333\,
            in2 => \_gnd_net_\,
            in3 => \N__13351\,
            lcout => \uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_0_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010011001100"
        )
    port map (
            in0 => \N__15824\,
            in1 => \N__15470\,
            in2 => \N__13379\,
            in3 => \N__14963\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16936\,
            ce => 'H',
            sr => \N__13602\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_3_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__15823\,
            in1 => \N__15755\,
            in2 => \_gnd_net_\,
            in3 => \N__15800\,
            lcout => \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16936\,
            ce => 'H',
            sr => \N__13602\
        );

    \uart_inst0.uart_inst0.rx_bits_remaining_RNINTCJ_2_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__15891\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15637\,
            lcout => \uart_inst0.uart_inst0.N_274_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_bits_remaining_RNO_0_2_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__16035\,
            in1 => \N__15969\,
            in2 => \_gnd_net_\,
            in3 => \N__15922\,
            lcout => \uart_inst0.uart_inst0.un1_rx_bits_remaining_c1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_state_RNID5M13_2_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16036\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15920\,
            lcout => \uart_inst0.uart_inst0.rx_bits_remaining_2_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_state_RNI4UTC3_1_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__15921\,
            in1 => \N__13298\,
            in2 => \_gnd_net_\,
            in3 => \N__13265\,
            lcout => \uart_inst0.uart_inst0.rx_state_2_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_countdown_RNID5M13_0_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__14081\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14035\,
            lcout => \uart_inst0.uart_inst0.rRxData_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_state_RNO_0_3_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__13946\,
            in1 => \N__13771\,
            in2 => \_gnd_net_\,
            in3 => \N__13829\,
            lcout => OPEN,
            ltout => \uart_inst0.uart_inst0.N_273_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_state_3_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__15655\,
            in1 => \N__13720\,
            in2 => \N__13790\,
            in3 => \N__13738\,
            lcout => \uart_inst0.uart_inst0.rx_stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16929\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_bits_remaining_RNINTCJ_3_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13696\,
            in2 => \_gnd_net_\,
            in3 => \N__15965\,
            lcout => \uart_inst0.uart_inst0.rx_state_srsts_0_a5_0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_bits_remaining_RNO_0_3_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010000000000"
        )
    port map (
            in0 => \N__13719\,
            in1 => \N__16037\,
            in2 => \N__15973\,
            in3 => \N__15923\,
            lcout => OPEN,
            ltout => \uart_inst0.uart_inst0.un1_rx_bits_remaining_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_bits_remaining_3_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000100010010"
        )
    port map (
            in0 => \N__13697\,
            in1 => \N__15864\,
            in2 => \N__13700\,
            in3 => \N__15654\,
            lcout => \uart_inst0.uart_inst0.rx_bits_remainingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16929\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_countdown_2_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001011011100"
        )
    port map (
            in0 => \N__13685\,
            in1 => \N__13629\,
            in2 => \N__13643\,
            in3 => \N__14459\,
            lcout => \uart_inst0.uart_inst0.tx_countdownZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16922\,
            ce => 'H',
            sr => \N__13597\
        );

    \uart_inst0.uart_inst0.tx_clk_divider_3_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101110100100010"
        )
    port map (
            in0 => \N__13548\,
            in1 => \N__13490\,
            in2 => \_gnd_net_\,
            in3 => \N__14419\,
            lcout => \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16916\,
            ce => 'H',
            sr => \N__14638\
        );

    \uart_inst0.uart_inst0.tx_countdown_RNO_2_2_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__14593\,
            in1 => \N__14551\,
            in2 => \_gnd_net_\,
            in3 => \N__14504\,
            lcout => OPEN,
            ltout => \uart_inst0.uart_inst0.tx_m5_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_countdown_RNO_1_2_LC_17_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14489\,
            in1 => \N__14380\,
            in2 => \N__14480\,
            in3 => \N__14477\,
            lcout => \uart_inst0.uart_inst0.tx_N_11_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.tx_clk_divider_RNIAEQ11_0_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14448\,
            in1 => \N__14431\,
            in2 => \N__14420\,
            in3 => \N__14397\,
            lcout => \uart_inst0.uart_inst0.tx_m5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ft2232h_inst.rRxData_5_LC_18_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__14366\,
            in1 => \N__17040\,
            in2 => \_gnd_net_\,
            in3 => \N__14356\,
            lcout => \fifo_inst.wRxWrData_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16988\,
            ce => 'H',
            sr => \N__16368\
        );

    \uart_inst0.tx_uart_fifo_inst.m54_e_5_LC_18_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14331\,
            in1 => \N__14307\,
            in2 => \N__14287\,
            in3 => \N__16658\,
            lcout => OPEN,
            ltout => \uart_inst0.tx_uart_fifo_inst.m54_eZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m54_e_LC_18_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__14244\,
            in1 => \N__14217\,
            in2 => \N__14201\,
            in3 => \N__14108\,
            lcout => \uart_inst0.tx_uart_fifo_inst.N_91\,
            ltout => \uart_inst0.tx_uart_fifo_inst.N_91_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rRamWrAddr_3_LC_18_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101001100000000"
        )
    port map (
            in0 => \N__14842\,
            in1 => \N__16657\,
            in2 => \N__14198\,
            in3 => \N__14195\,
            lcout => \fifo_inst_rx_fifo_inst_rRamWrAddr_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16984\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.m54_e_6_LC_18_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__14181\,
            in1 => \N__14154\,
            in2 => \N__14131\,
            in3 => \N__14796\,
            lcout => \uart_inst0.tx_uart_fifo_inst.m54_eZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.rRamWrAddr_0_LC_18_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001010001010"
        )
    port map (
            in0 => \N__14855\,
            in1 => \N__14849\,
            in2 => \N__16700\,
            in3 => \N__14841\,
            lcout => \fifo_inst_rx_fifo_inst_rRamWrAddr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16984\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_4_LC_18_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__15412\,
            in1 => \N__14770\,
            in2 => \_gnd_net_\,
            in3 => \N__14780\,
            lcout => \wRxData_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_4C_net\,
            ce => \N__15308\,
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_3_LC_18_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__15411\,
            in1 => \N__14749\,
            in2 => \_gnd_net_\,
            in3 => \N__14756\,
            lcout => \wRxData_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_4C_net\,
            ce => \N__15308\,
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7_LC_18_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15402\,
            in1 => \N__14735\,
            in2 => \_gnd_net_\,
            in3 => \N__14729\,
            lcout => \wRxData_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7C_net\,
            ce => \N__15304\,
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_5_LC_18_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__15400\,
            in1 => \N__14711\,
            in2 => \_gnd_net_\,
            in3 => \N__14717\,
            lcout => \wRxData_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7C_net\,
            ce => \N__15304\,
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_1_LC_18_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14693\,
            in1 => \N__14699\,
            in2 => \_gnd_net_\,
            in3 => \N__15398\,
            lcout => \wRxData_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7C_net\,
            ce => \N__15304\,
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_2_LC_18_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__15399\,
            in1 => \N__14672\,
            in2 => \_gnd_net_\,
            in3 => \N__14678\,
            lcout => \wRxData_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7C_net\,
            ce => \N__15304\,
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_6_LC_18_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__15401\,
            in1 => \N__14654\,
            in2 => \_gnd_net_\,
            in3 => \N__14660\,
            lcout => \wRxData_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7C_net\,
            ce => \N__15304\,
            sr => \_gnd_net_\
        );

    \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_0_LC_18_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__15320\,
            in1 => \N__15425\,
            in2 => \_gnd_net_\,
            in3 => \N__15397\,
            lcout => \wRxData_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7C_net\,
            ce => \N__15304\,
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNIRP0T_8_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15276\,
            in2 => \_gnd_net_\,
            in3 => \N__15252\,
            lcout => OPEN,
            ltout => \uart_inst0.rx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNIMIH82_0_LC_18_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__15229\,
            in1 => \N__15202\,
            in2 => \N__15182\,
            in3 => \N__15172\,
            lcout => \uart_inst0.rx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNIMJ1Q1_4_LC_18_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15127\,
            in1 => \N__15100\,
            in2 => \N__15079\,
            in3 => \N__15043\,
            lcout => \uart_inst0.rx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_5_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15014\,
            in1 => \N__15007\,
            in2 => \_gnd_net_\,
            in3 => \N__14947\,
            lcout => \wUartRxData_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_5C_net\,
            ce => \N__14879\,
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_6_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__14946\,
            in1 => \_gnd_net_\,
            in2 => \N__14993\,
            in3 => \N__14983\,
            lcout => \wUartRxData_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_5C_net\,
            ce => \N__14879\,
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_7_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__14893\,
            in1 => \N__14969\,
            in2 => \_gnd_net_\,
            in3 => \N__14948\,
            lcout => \wUartRxData_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_5C_net\,
            ce => \N__14879\,
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_0_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14870\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \wUartRxData_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net\,
            ce => \N__15789\,
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_1_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15572\,
            lcout => \wUartRxData_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net\,
            ce => \N__15789\,
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_2_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15557\,
            lcout => \wUartRxData_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net\,
            ce => \N__15789\,
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_3_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15542\,
            lcout => \wUartRxData_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net\,
            ce => \N__15789\,
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_4_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15527\,
            lcout => \wUartRxData_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net\,
            ce => \N__15789\,
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_5_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16684\,
            in2 => \_gnd_net_\,
            in3 => \N__15511\,
            lcout => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_3_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16686\,
            in2 => \_gnd_net_\,
            in3 => \N__15490\,
            lcout => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__15822\,
            in1 => \N__15466\,
            in2 => \N__16703\,
            in3 => \N__15794\,
            lcout => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_4_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16687\,
            in2 => \_gnd_net_\,
            in3 => \N__15445\,
            lcout => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_2_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100000000"
        )
    port map (
            in0 => \N__16685\,
            in1 => \N__15821\,
            in2 => \N__15799\,
            in3 => \N__15751\,
            lcout => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_6_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16688\,
            in2 => \_gnd_net_\,
            in3 => \N__15730\,
            lcout => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_1_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16683\,
            in2 => \_gnd_net_\,
            in3 => \N__15709\,
            lcout => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_7_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16689\,
            in2 => \_gnd_net_\,
            in3 => \N__15688\,
            lcout => \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rx_bits_remaining_2_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110000101111000"
        )
    port map (
            in0 => \N__15896\,
            in1 => \N__15668\,
            in2 => \N__15641\,
            in3 => \N__15659\,
            lcout => \uart_inst0.uart_inst0.rx_bits_remainingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16945\,
            ce => 'H',
            sr => \N__15874\
        );

    \uart_inst0.uart_inst0.rx_bits_remaining_0_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__15938\,
            in1 => \N__15964\,
            in2 => \_gnd_net_\,
            in3 => \N__16049\,
            lcout => \uart_inst0.uart_inst0.rx_bits_remainingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16945\,
            ce => 'H',
            sr => \N__15874\
        );

    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_1_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16694\,
            in2 => \_gnd_net_\,
            in3 => \N__15622\,
            lcout => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_4_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16695\,
            in2 => \_gnd_net_\,
            in3 => \N__15596\,
            lcout => \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uart_inst0.uart_inst0.rRxData_esr_1_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16081\,
            lcout => \uart_inst0.wRxWrData_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16940\,
            ce => \N__16067\,
            sr => \N__16454\
        );

    \uart_inst0.uart_inst0.rRxData_esr_4_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16162\,
            lcout => \uart_inst0.wRxWrData_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16940\,
            ce => \N__16067\,
            sr => \N__16454\
        );

    \uart_inst0.uart_inst0.rRxData_esr_3_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16210\,
            lcout => \uart_inst0.wRxWrData_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16940\,
            ce => \N__16067\,
            sr => \N__16454\
        );

    \uart_inst0.uart_inst0.rRxData_esr_0_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16192\,
            lcout => \uart_inst0.wRxWrData_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16940\,
            ce => \N__16067\,
            sr => \N__16454\
        );

    \uart_inst0.uart_inst0.rRxData_esr_5_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16114\,
            lcout => \uart_inst0.wRxWrData_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16940\,
            ce => \N__16067\,
            sr => \N__16454\
        );

    \uart_inst0.uart_inst0.rRxData_esr_6_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16148\,
            lcout => \uart_inst0.wRxWrData_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16940\,
            ce => \N__16067\,
            sr => \N__16454\
        );

    \uart_inst0.uart_inst0.rRxData_esr_2_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16096\,
            lcout => \uart_inst0.wRxWrData_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16937\,
            ce => \N__16066\,
            sr => \N__16455\
        );

    \uart_inst0.uart_inst0.rx_bits_remaining_1_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010011010101010"
        )
    port map (
            in0 => \N__15895\,
            in1 => \N__16048\,
            in2 => \N__15974\,
            in3 => \N__15933\,
            lcout => \uart_inst0.uart_inst0.rx_bits_remainingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16932\,
            ce => 'H',
            sr => \N__15875\
        );

    \fifo_inst.ft2232h_inst.rRxData_2_LC_20_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__15848\,
            in1 => \N__17060\,
            in2 => \_gnd_net_\,
            in3 => \N__15836\,
            lcout => \fifo_inst.wRxWrData_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16989\,
            ce => 'H',
            sr => \N__16419\
        );

    \fifo_inst.ft2232h_inst.rRxData_1_LC_20_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__17225\,
            in1 => \N__17059\,
            in2 => \_gnd_net_\,
            in3 => \N__17209\,
            lcout => \fifo_inst.wRxWrData_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16989\,
            ce => 'H',
            sr => \N__16419\
        );

    \fifo_inst.ft2232h_inst.rRxData_3_LC_20_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17061\,
            in1 => \N__17195\,
            in2 => \_gnd_net_\,
            in3 => \N__17182\,
            lcout => \fifo_inst.wRxWrData_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16989\,
            ce => 'H',
            sr => \N__16419\
        );

    \fifo_inst.ft2232h_inst.rRxData_4_LC_20_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__17168\,
            in1 => \N__17062\,
            in2 => \_gnd_net_\,
            in3 => \N__17156\,
            lcout => \fifo_inst.wRxWrData_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16989\,
            ce => 'H',
            sr => \N__16419\
        );

    \fifo_inst.ft2232h_inst.rRxData_0_LC_20_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__17144\,
            in1 => \N__17058\,
            in2 => \_gnd_net_\,
            in3 => \N__17129\,
            lcout => \fifo_inst.wRxWrData_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16989\,
            ce => 'H',
            sr => \N__16419\
        );

    \fifo_inst.ft2232h_inst.rRxData_7_LC_20_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__17063\,
            in1 => \N__17117\,
            in2 => \_gnd_net_\,
            in3 => \N__17096\,
            lcout => \fifo_inst.wRxWrData_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16989\,
            ce => 'H',
            sr => \N__16419\
        );

    \fifo_inst.ft2232h_inst.rRxData_6_LC_20_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__17084\,
            in1 => \N__17057\,
            in2 => \_gnd_net_\,
            in3 => \N__17005\,
            lcout => \fifo_inst.wRxWrData_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__16987\,
            ce => 'H',
            sr => \N__16421\
        );
end \INTERFACE\;
