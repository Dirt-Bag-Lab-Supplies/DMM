-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Mar 29 2020 02:25:20

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    ioFifoData : inout std_logic_vector(7 downto 0);
    P1A9 : out std_logic;
    P1A1 : in std_logic;
    P1A8 : out std_logic;
    oRx_n : out std_logic;
    P1A7 : out std_logic;
    P1A3 : out std_logic;
    iTxE_n : in std_logic;
    iRxF_n : in std_logic;
    iClk : in std_logic;
    P1A2 : out std_logic;
    BTN_N : in std_logic;
    BTN1 : in std_logic;
    oTx_n : out std_logic;
    P1A4 : out std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__15651\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15627\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15617\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15608\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15599\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15574\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15572\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15564\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15556\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15545\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15536\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15502\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15493\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15483\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15465\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15447\ : std_logic;
signal \N__15444\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15438\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15423\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15417\ : std_logic;
signal \N__15414\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15410\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15360\ : std_logic;
signal \N__15359\ : std_logic;
signal \N__15358\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15343\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15290\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15286\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15283\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15280\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15278\ : std_logic;
signal \N__15275\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15253\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15241\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15232\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15229\ : std_logic;
signal \N__15226\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15177\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15168\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15154\ : std_logic;
signal \N__15151\ : std_logic;
signal \N__15148\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15107\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15086\ : std_logic;
signal \N__15083\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15081\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15053\ : std_logic;
signal \N__15052\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15049\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15047\ : std_logic;
signal \N__15046\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15043\ : std_logic;
signal \N__15042\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15040\ : std_logic;
signal \N__15039\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15026\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15023\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15021\ : std_logic;
signal \N__15020\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15015\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15013\ : std_logic;
signal \N__15012\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15005\ : std_logic;
signal \N__15004\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__15001\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14859\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14853\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14836\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14826\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14823\ : std_logic;
signal \N__14820\ : std_logic;
signal \N__14819\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14816\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14813\ : std_logic;
signal \N__14812\ : std_logic;
signal \N__14809\ : std_logic;
signal \N__14806\ : std_logic;
signal \N__14789\ : std_logic;
signal \N__14786\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14777\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14773\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14767\ : std_logic;
signal \N__14764\ : std_logic;
signal \N__14761\ : std_logic;
signal \N__14758\ : std_logic;
signal \N__14755\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14737\ : std_logic;
signal \N__14730\ : std_logic;
signal \N__14727\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14707\ : std_logic;
signal \N__14704\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14694\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14679\ : std_logic;
signal \N__14676\ : std_logic;
signal \N__14673\ : std_logic;
signal \N__14670\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14666\ : std_logic;
signal \N__14663\ : std_logic;
signal \N__14658\ : std_logic;
signal \N__14655\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14649\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14633\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14613\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14604\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14589\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14576\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14568\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14562\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14552\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14549\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14537\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14517\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14508\ : std_logic;
signal \N__14505\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14497\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14457\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14452\ : std_logic;
signal \N__14451\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14436\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14428\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14421\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14358\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14343\ : std_logic;
signal \N__14340\ : std_logic;
signal \N__14337\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14330\ : std_logic;
signal \N__14325\ : std_logic;
signal \N__14324\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14322\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14307\ : std_logic;
signal \N__14304\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14289\ : std_logic;
signal \N__14286\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14280\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14274\ : std_logic;
signal \N__14271\ : std_logic;
signal \N__14268\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14235\ : std_logic;
signal \N__14232\ : std_logic;
signal \N__14229\ : std_logic;
signal \N__14226\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14209\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14175\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14172\ : std_logic;
signal \N__14169\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14157\ : std_logic;
signal \N__14156\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14136\ : std_logic;
signal \N__14133\ : std_logic;
signal \N__14130\ : std_logic;
signal \N__14127\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14120\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14100\ : std_logic;
signal \N__14097\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14066\ : std_logic;
signal \N__14063\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14057\ : std_logic;
signal \N__14054\ : std_logic;
signal \N__14051\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14037\ : std_logic;
signal \N__14034\ : std_logic;
signal \N__14031\ : std_logic;
signal \N__14028\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14022\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14016\ : std_logic;
signal \N__14015\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__13991\ : std_logic;
signal \N__13986\ : std_logic;
signal \N__13983\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13968\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13953\ : std_logic;
signal \N__13950\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13947\ : std_logic;
signal \N__13944\ : std_logic;
signal \N__13937\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13928\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13926\ : std_logic;
signal \N__13925\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13910\ : std_logic;
signal \N__13905\ : std_logic;
signal \N__13902\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13896\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13872\ : std_logic;
signal \N__13869\ : std_logic;
signal \N__13866\ : std_logic;
signal \N__13863\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13857\ : std_logic;
signal \N__13854\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13848\ : std_logic;
signal \N__13845\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13836\ : std_logic;
signal \N__13833\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13824\ : std_logic;
signal \N__13821\ : std_logic;
signal \N__13818\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13815\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13812\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13809\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13802\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13778\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13755\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13746\ : std_logic;
signal \N__13743\ : std_logic;
signal \N__13740\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13738\ : std_logic;
signal \N__13737\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13735\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13731\ : std_logic;
signal \N__13730\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13721\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13709\ : std_logic;
signal \N__13708\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13704\ : std_logic;
signal \N__13701\ : std_logic;
signal \N__13700\ : std_logic;
signal \N__13697\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13647\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13630\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13624\ : std_logic;
signal \N__13621\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13588\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13582\ : std_logic;
signal \N__13579\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13566\ : std_logic;
signal \N__13563\ : std_logic;
signal \N__13560\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13548\ : std_logic;
signal \N__13545\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13528\ : std_logic;
signal \N__13525\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13515\ : std_logic;
signal \N__13512\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13506\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13491\ : std_logic;
signal \N__13488\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13480\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13461\ : std_logic;
signal \N__13458\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13446\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13437\ : std_logic;
signal \N__13434\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13417\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13409\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13377\ : std_logic;
signal \N__13374\ : std_logic;
signal \N__13371\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13366\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13362\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13356\ : std_logic;
signal \N__13353\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13338\ : std_logic;
signal \N__13337\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13335\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13311\ : std_logic;
signal \N__13308\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13302\ : std_logic;
signal \N__13299\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13285\ : std_logic;
signal \N__13282\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13257\ : std_logic;
signal \N__13254\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13248\ : std_logic;
signal \N__13245\ : std_logic;
signal \N__13242\ : std_logic;
signal \N__13239\ : std_logic;
signal \N__13236\ : std_logic;
signal \N__13233\ : std_logic;
signal \N__13230\ : std_logic;
signal \N__13227\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13212\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13206\ : std_logic;
signal \N__13203\ : std_logic;
signal \N__13200\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13191\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13176\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13164\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13158\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13149\ : std_logic;
signal \N__13146\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13108\ : std_logic;
signal \N__13105\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13058\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13047\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13028\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12996\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12984\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12976\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12958\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12939\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12895\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12874\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12868\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12838\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12768\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12714\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12684\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12678\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12605\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12589\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12549\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12388\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12308\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12302\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12289\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11154\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10941\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10707\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10562\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10506\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9807\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8136\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8055\ : std_logic;
signal \N__8052\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7992\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7893\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7827\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7821\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7641\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7578\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7551\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7434\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7260\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6048\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5862\ : std_logic;
signal \wRamRdData_1\ : std_logic;
signal \wRamRdData_6\ : std_logic;
signal \wRamRdData_2\ : std_logic;
signal \wRamRdData_5\ : std_logic;
signal \wRamRdData_4\ : std_logic;
signal \BTN_N_c\ : std_logic;
signal \wRamRdData_7\ : std_logic;
signal \wRamRdData_0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \wRamRdData_3\ : std_logic;
signal \GNDG0\ : std_logic;
signal \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO\ : std_logic;
signal \top_pll_inst.wPllLocked_iso_i\ : std_logic;
signal \DUT.uart_inst0.N_6_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_22_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_22\ : std_logic;
signal \DUT.uart_inst0.g2_3_cascade_\ : std_logic;
signal \DUT.uart_inst0.g2\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_9\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_8\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_6_cascade_\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_7\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_152_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_5\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_7_m1_0_o2_2_2_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_out_6_iv_0_a3_0_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_out_6_iv_0_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_119\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_RNO_0Z0Z_4_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.m25_e_3_cascade_\ : std_logic;
signal \DUT.uart_inst0.m3_0\ : std_logic;
signal \bfn_13_7_0_\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_0\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_1\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_2\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_3\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_4\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_5\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_6\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_7\ : std_logic;
signal \bfn_13_8_0_\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_8\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_9\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_10\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_11\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_12\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_13\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_14\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_15\ : std_logic;
signal \bfn_13_9_0_\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_16\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0\ : std_logic;
signal \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoCount_RNISSQ21Z0Z_1\ : std_logic;
signal \DUT.fifo_tx_inst.N_108_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0\ : std_logic;
signal \DUT.fifo_tx_inst.N_108\ : std_logic;
signal \rTxWriteZ0\ : std_logic;
signal \DUT.fifo_tx_inst.N_104_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_8_i_o2_1_2_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_67\ : std_logic;
signal \DUT.uart_inst0.g0_0_0_a3_0_3_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_159_0\ : std_logic;
signal \DUT.uart_inst0.N_4\ : std_logic;
signal \bfn_14_2_0_\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_0\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_1\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_2\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_3\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_4\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_6\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_5\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_7\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_6\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_7\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_8\ : std_logic;
signal \bfn_14_3_0_\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_9\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_8\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_10\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_9\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_11\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_10\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_12\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_11\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_12\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_13\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remainingZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remainingZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.m9_e_0_3\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remainingZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.m9_e_0_0\ : std_logic;
signal \DUT.uart_inst0.N_152\ : std_logic;
signal \DUT.uart_inst0.tx_state_0_sqmuxa_i_i_a3_c_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_160_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_0_ac0_1\ : std_logic;
signal \DUT.uart_inst0.N_154\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remainingZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.N_72\ : std_logic;
signal \DUT.uart_inst0.N_99\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_RNO_0Z0Z_1\ : std_logic;
signal \DUT.uart_inst0.N_88_i\ : std_logic;
signal \DUT.uart_inst0.N_160\ : std_logic;
signal \DUT.uart_inst0.N_218\ : std_logic;
signal \DUT.uart_inst0.N_218_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_109\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.N_120\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_RNO_1Z0Z_3_cascade_\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_0\ : std_logic;
signal \DUT.uart_inst0.N_164\ : std_logic;
signal \DUT.uart_inst0.N_164_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_RNO_0Z0Z_3\ : std_logic;
signal \DUT.uart_inst0.tx_state_ns_i_i_o2_a0_2_0\ : std_logic;
signal \DUT.uart_inst0.N_159\ : std_logic;
signal \DUT.uart_inst0.N_100\ : std_logic;
signal \DUT.uart_inst0.N_163\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_0_c3\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_30_5\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_7_m1_0_a3_0_2\ : std_logic;
signal \DUT.uart_inst0.N_113\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_7_sm0_0\ : std_logic;
signal \DUT.uart_inst0.N_84\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_17\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_13\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_14\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_15\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_10\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_9\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_11\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_7\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_5\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_6\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_6\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_8\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_12\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.m7_e_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.m7_e_3_cascade_\ : std_logic;
signal \DUT.uart_inst0.m9_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_11_mux\ : std_logic;
signal \DUT.uart_inst0.N_66\ : std_logic;
signal \DUT.uart_inst0.m4_e_0\ : std_logic;
signal \DUT.uart_inst0.m4_e_3\ : std_logic;
signal \DUT.uart_inst0.N_21_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_21_mux_0\ : std_logic;
signal \DUT.uart_inst0.m5_1\ : std_logic;
signal \DUT.uart_inst0.N_6\ : std_logic;
signal \DUT.uart_inst0.N_6_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_18\ : std_logic;
signal \DUT.uart_inst0.N_18_mux_0\ : std_logic;
signal \DUT.uart_inst0.N_30\ : std_logic;
signal \DUT.uart_inst0.g1_i_a4_0_4\ : std_logic;
signal \DUT.uart_inst0.g1_i_a4_0_5_cascade_\ : std_logic;
signal \DUT.uart_inst0.g0_0_0_a3_0_4\ : std_logic;
signal \DUT.uart_inst0.g0_0_0_a3_4_cascade_\ : std_logic;
signal \DUT.uart_inst0.g0_0_0_a3_3\ : std_logic;
signal \DUT.fifo_tx_inst.un1_i11_i_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.N_57_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.un1_i11_i\ : std_logic;
signal \DUT.uart_inst0.m13_2_cascade_\ : std_logic;
signal \DUT.uart_inst0.m13_3\ : std_logic;
signal \DUT.uart_inst0.P19_mux_cascade_\ : std_logic;
signal \DUT.uart_inst0.g0_0_1\ : std_logic;
signal \N_1257_i\ : std_logic;
signal \G_111_cascade_\ : std_logic;
signal \fifo_inst.ftdi_input_inst.SUMZ0Z_2_cascade_\ : std_logic;
signal \G_110_cascade_\ : std_logic;
signal \fifo_inst_ftdi_input_inst_oTxFull_0\ : std_logic;
signal \G_108\ : std_logic;
signal \fifo_inst.ftdi_input_inst.SUMZ0Z_3\ : std_logic;
signal \G_109\ : std_logic;
signal \G_110\ : std_logic;
signal \G_111\ : std_logic;
signal \G_112\ : std_logic;
signal \fifo_inst.ftdi_input_inst.un2_oPacketAvail_iZ0\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_0\ : std_logic;
signal \P1A7_c\ : std_logic;
signal \DUT.uart_inst0.N_116\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_7\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_6\ : std_logic;
signal \DUT.uart_inst0.N_22_i\ : std_logic;
signal \DUT.uart_inst0.N_102\ : std_logic;
signal \DUT.uart_inst0.tx_state_0_sqmuxa_i_i_a3_0_1\ : std_logic;
signal \DUT.tx_state_1\ : std_logic;
signal \DUT.N_114_cascade_\ : std_logic;
signal \DUT.tx_state_0\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_16\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_9_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ1Z_1\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_3\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.m6_3_cascade_\ : std_logic;
signal \top_pll_inst.m12_1_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.G_30_1\ : std_logic;
signal \P18_mux_cascade_\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_11\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_10\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_12\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_13\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_0_cascade_\ : std_logic;
signal \bfn_15_9_0_\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_0_s1\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_1_s1\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_2_s1\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_3_s1\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_4_s1\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.N_20\ : std_logic;
signal \DUT.uart_inst0.N_21_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_21_mux_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_19_mux\ : std_logic;
signal \DUT.uart_inst0.N_13_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_13_0\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_8_i_o2_2_0_2_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.un1_i11_i\ : std_logic;
signal \DUT.uart_inst0.g0_0\ : std_logic;
signal \DUT.uart_inst0.N_49\ : std_logic;
signal \DUT.uart_inst0.m6_1\ : std_logic;
signal \DUT.uart_inst0.N_7\ : std_logic;
signal \DUT.uart_inst0.recv_state_srsts_1_5\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_8_i_o2_2_2\ : std_logic;
signal \DUT.uart_inst0.recv_state_srsts_1_5_cascade_\ : std_logic;
signal \DUT.uart_inst0.recv_state_srsts_1_4\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.N_43_cascade_\ : std_logic;
signal \DUT.uart_inst0.recv_state_RNIL139CZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.m3_e_1_cascade_\ : std_logic;
signal \DUT_uart_inst0_recv_state_2\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remainingZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remainingZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remainingZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remainingZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.recv_state_RNO_4Z0Z_2\ : std_logic;
signal \DUT.uart_inst0.N_19\ : std_logic;
signal \DUT.uart_inst0.G_8_i_a3_0_0\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_8_i_o2_1_1_2\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_\ : std_logic;
signal \DUT.rFifoDatarx_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_\ : std_logic;
signal \DUT.rFifoDatarx_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1_cascade_\ : std_logic;
signal \DUT.rFifoDatarx_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_\ : std_logic;
signal \DUT.rFifoDatarx_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_\ : std_logic;
signal \DUT.rFifoDatarx_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_6\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_\ : std_logic;
signal \DUT.rFifoDatarx_6\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoCountZ0Z_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoCountZ0Z_0\ : std_logic;
signal \DUT.rTransmitZ0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoCountZ0Z_2\ : std_logic;
signal \DUT.fifo_tx_inst.rReadPtr11_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.un1_i11_2_i_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rReadPtr11\ : std_logic;
signal \DUT.fifo_tx_inst.un1_i11_2_i\ : std_logic;
signal \DUT.rFifoDataror_1\ : std_logic;
signal \DUT.rFifoDataror_1_cascade_\ : std_logic;
signal \DUT.rFifoDataror_0_0\ : std_logic;
signal \DUT.rFifoDataror_0\ : std_logic;
signal \G_115\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa\ : std_logic;
signal \DUT.uart_inst0.m6_2\ : std_logic;
signal \G_114\ : std_logic;
signal \G_113\ : std_logic;
signal \fifo_inst.ftdi_input_inst.un1_rWrStateZ0Z_1_cascade_\ : std_logic;
signal \G_118\ : std_logic;
signal \G_118_cascade_\ : std_logic;
signal \G_119\ : std_logic;
signal \G_116\ : std_logic;
signal \fifo_inst.ftdi_input_inst.un1_rWrStateZ0Z_1\ : std_logic;
signal \G_116_cascade_\ : std_logic;
signal \G_117\ : std_logic;
signal \DUT.uart_inst0.g1_i_a4_1_5\ : std_logic;
signal \DUT.uart_inst0.g1_i_a4_1_3\ : std_logic;
signal \DUT.uart_inst0.N_78_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_10_mux_cascade_\ : std_logic;
signal \DUT.uart_inst0.P6_mux\ : std_logic;
signal \DUT.uart_inst0.G_19_0_a5_0_2_cascade_\ : std_logic;
signal \DUT.uart_inst0.G_19_0_1\ : std_logic;
signal \DUT.uart_inst0.G_19_0_a5_0_4_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_8_i_o2_2_0_2\ : std_logic;
signal \DUT.uart_inst0.G_8_i_a3_1\ : std_logic;
signal \DUT_uart_inst0_rx_countdown_3_s1_4\ : std_logic;
signal \DUT_uart_inst0_rx_countdown_3_s1_5\ : std_logic;
signal \DUT_uart_inst0_rx_countdown_3_s1_3\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_3\ : std_logic;
signal \DUT_uart_inst0_rx_countdown_3_s1_2\ : std_logic;
signal \DUT_uart_inst0_rx_countdown_3_s1_1\ : std_logic;
signal \DUT.uart_inst0.G_19_0_a5_4\ : std_logic;
signal \DUT.uart_inst0.N_44\ : std_logic;
signal \DUT.fifo_rx_inst.N_77_mux\ : std_logic;
signal \DUT.uart_inst0.g1_0\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_8_i_a2_0_2\ : std_logic;
signal \DUT.uart_inst0.m10_e_3\ : std_logic;
signal \DUT.uart_inst0.m10_e_2\ : std_logic;
signal \wPllLocked\ : std_logic;
signal \DUT.uart_inst0.N_20_mux_cascade_\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_0\ : std_logic;
signal \DUT.uart_inst0.m7_3_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_28_mux\ : std_logic;
signal \P1A1_c\ : std_logic;
signal \DUT.uart_inst0.m2_e_0\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.m6_e_2\ : std_logic;
signal \DUT.uart_inst0.m6_e_3_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_15_mux\ : std_logic;
signal \DUT.uart_inst0.N_18_mux_1\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ1Z_3\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.G_19_0_a5_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_6\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_\ : std_logic;
signal \DUT.rFifoDatarx_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_2\ : std_logic;
signal \DUT.fifo_tx_inst.rReadPtrZ0Z_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rReadPtrZ0Z_1\ : std_logic;
signal \DUT.rFifoDatarx_3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_6\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_awe0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoDataro_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_awe1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoDataro_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoDataro_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoDataro_3\ : std_logic;
signal \DUT.fifo_rx_inst.N_57\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_6\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_6\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDataro_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDataror_1_0_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_5\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDataro_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDataro_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDataro_2\ : std_logic;
signal \DUT.fifo_rx_inst.rWritePtrZ0Z_0\ : std_logic;
signal \DUT.fifo_rx_inst.rWritePtrZ0Z_1\ : std_logic;
signal \DUT.fifo_tx_inst.rWritePtrZ0Z_0\ : std_logic;
signal \DUT.fifo_tx_inst.rWritePtrZ0Z_1\ : std_logic;
signal \DUT.fifo_tx_inst.N_104\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_awe2\ : std_logic;
signal \DUT.fifo_rx_inst.rWritePtr16_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rWritePtr16\ : std_logic;
signal \DUT.wRcvd\ : std_logic;
signal \DUT.fifo_rx_inst.N_46\ : std_logic;
signal \N_69_mux\ : std_logic;
signal \N_69_mux_cascade_\ : std_logic;
signal \N_1258_i\ : std_logic;
signal \P1A4_c_i\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_6\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_awe3\ : std_logic;
signal \ioFifoData_in_3\ : std_logic;
signal \ioFifoData_in_1\ : std_logic;
signal \ioFifoData_in_5\ : std_logic;
signal \ioFifoData_in_2\ : std_logic;
signal \ioFifoData_in_0\ : std_logic;
signal \ioFifoData_in_6\ : std_logic;
signal \ioFifoData_in_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_5\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_6\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_awe2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDatarx_6\ : std_logic;
signal \wRxFifoData_6\ : std_logic;
signal \rTxByteZ0Z_6\ : std_logic;
signal \wRxFifoData_5\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDatarx_5\ : std_logic;
signal \rTxByteZ0Z_5\ : std_logic;
signal \wRxFifoData_0\ : std_logic;
signal \rTxByteZ0Z_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDatarx_7\ : std_logic;
signal \rTxByteZ0Z_7\ : std_logic;
signal \wRxFifoData_1\ : std_logic;
signal \rTxByteZ0Z_1\ : std_logic;
signal \wRxFifoData_2\ : std_logic;
signal \rTxByteZ0Z_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDatarx_3\ : std_logic;
signal \wRxFifoData_3\ : std_logic;
signal \rTxByteZ0Z_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDataror_0\ : std_logic;
signal \wRxFifoData_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDatarx_4\ : std_logic;
signal \rTxByteZ0Z_4\ : std_logic;
signal \rTxByte_1_sqmuxa_i_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDatarx_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDatarx_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_1\ : std_logic;
signal \DUT.fifo_rx_inst.rReadPtrZ0Z_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rReadPtrZ0Z_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDatarx_2\ : std_logic;
signal \DUT.wRxByte_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_0\ : std_logic;
signal \DUT.wRxByte_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_2\ : std_logic;
signal \DUT.wRxByte_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_3\ : std_logic;
signal \DUT.wRxByte_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_5\ : std_logic;
signal \DUT.wRxByte_6\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_6\ : std_logic;
signal \DUT.wRxByte_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_awe1\ : std_logic;
signal \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoCountZ0Z_0\ : std_logic;
signal \bfn_18_12_0_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoCount_RNIPTFQ1Z0Z_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoCountZ0Z_1\ : std_logic;
signal \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0\ : std_logic;
signal \DUT.fifo_rx_inst.N_4_0\ : std_logic;
signal \rRxReadZ0\ : std_logic;
signal \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoCountZ0Z_2\ : std_logic;
signal \N_1261_i\ : std_logic;
signal \oTx_n_rep4_ess\ : std_logic;
signal \oTx_n_rep1_ess\ : std_logic;
signal \oTx_n_rep0_ess\ : std_logic;
signal \fifo_inst.ftdi_output_inst.N_77_0_cascade_\ : std_logic;
signal \P1A4_c\ : std_logic;
signal \fifo_inst.ftdi_output_inst.oPacketRead_1_sqmuxa_1_cascade_\ : std_logic;
signal \fifo_inst.wRamRdAddr_0\ : std_logic;
signal \fifo_inst.wRamRdAddr_1\ : std_logic;
signal \fifo_inst.ftdi_output_inst.oPacketRead_1_sqmuxa_1\ : std_logic;
signal \fifo_inst.wRamRdAddr_2\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_3\ : std_logic;
signal \P1A2_c\ : std_logic;
signal \P1A3_c\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1\ : std_logic;
signal \iTxE_n_c\ : std_logic;
signal \iRxF_n_c\ : std_logic;
signal \G_120\ : std_logic;
signal \wPllLocked_g\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2\ : std_logic;
signal \fifo_inst.ftdi_output_inst.N_87_cascade_\ : std_logic;
signal \fifo_inst.ftdi_output_inst.N_77_0\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0\ : std_logic;
signal \ioFifoData_in_7\ : std_logic;
signal \wRxFifoData_7\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rFifoState_0_1\ : std_logic;
signal \N_1260_i\ : std_logic;
signal \N_1259_i\ : std_logic;
signal \oTx_n_rep3_ess\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rWrDelayZ0\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4\ : std_logic;
signal \oTx_n_rep2_ess\ : std_logic;
signal \fifo_inst.ftdi_output_inst.N_88_i_0\ : std_logic;
signal \wPllLocked_iso_i_g\ : std_logic;
signal \DUT.wRxByte_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_2\ : std_logic;
signal \DUT.wRxByte_5\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_5\ : std_logic;
signal clk_48mhz : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_awe0\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \iClk_wire\ : std_logic;
signal \P1A8_wire\ : std_logic;
signal \P1A4_wire\ : std_logic;
signal \oRx_n_wire\ : std_logic;
signal \P1A2_wire\ : std_logic;
signal \iRxF_n_wire\ : std_logic;
signal \P1A3_wire\ : std_logic;
signal \P1A7_wire\ : std_logic;
signal \BTN_N_wire\ : std_logic;
signal \oTx_n_wire\ : std_logic;
signal \iTxE_n_wire\ : std_logic;
signal \P1A1_wire\ : std_logic;
signal \P1A9_wire\ : std_logic;
signal \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \top_pll_inst.top_pll_inst_pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \iClk_wire\ <= iClk;
    P1A8 <= \P1A8_wire\;
    P1A4 <= \P1A4_wire\;
    oRx_n <= \oRx_n_wire\;
    P1A2 <= \P1A2_wire\;
    \iRxF_n_wire\ <= iRxF_n;
    P1A3 <= \P1A3_wire\;
    P1A7 <= \P1A7_wire\;
    \BTN_N_wire\ <= BTN_N;
    oTx_n <= \oTx_n_wire\;
    \iTxE_n_wire\ <= iTxE_n;
    \P1A1_wire\ <= P1A1;
    P1A9 <= \P1A9_wire\;
    \wRamRdData_7\ <= \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RDATA_wire\(14);
    \wRamRdData_6\ <= \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RDATA_wire\(12);
    \wRamRdData_5\ <= \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RDATA_wire\(10);
    \wRamRdData_4\ <= \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RDATA_wire\(8);
    \wRamRdData_3\ <= \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RDATA_wire\(6);
    \wRamRdData_2\ <= \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RDATA_wire\(4);
    \wRamRdData_1\ <= \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RDATA_wire\(2);
    \wRamRdData_0\ <= \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RDATA_wire\(0);
    \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__14130\&\N__14157\&\N__14178\;
    \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__9711\&\N__9648\&\N__9684\;
    \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \top_pll_inst.top_pll_inst_pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \fifo_inst.ftdi_input_inst.ram512x8_inst_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RDATA_wire\,
            RADDR => \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RADDR_wire\,
            WADDR => \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_WADDR_wire\,
            MASK => \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_MASK_wire\,
            WDATA => \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \GNDG0\,
            RE => \N__9179\,
            WCLKE => 'H',
            WCLK => \N__15047\,
            WE => \N__9569\
        );

    \top_pll_inst.top_pll_inst_pll\ : PLL40
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "0111111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            PLLOUTGLOBAL => clk_48mhz,
            SDI => \GNDG0\,
            BYPASS => \GNDG0\,
            RESETB => \N__5949\,
            PLLOUTCORE => OPEN,
            LOCK => \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO\,
            SDO => OPEN,
            SCLK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            EXTFEEDBACK => \GNDG0\,
            DYNAMICDELAY => \top_pll_inst.top_pll_inst_pll_DYNAMICDELAY_wire\,
            PLLIN => \N__15651\
        );

    \top_pll_inst.top_pll_inst_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \VCCG0\,
            DIN => '0',
            DOUT => \N__15651\,
            PACKAGEPIN => \iClk_wire\
        );

    \P1A8_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15637\,
            DIN => \N__15636\,
            DOUT => \N__15635\,
            PACKAGEPIN => \P1A8_wire\
        );

    \P1A8_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__15637\,
            PADOUT => \N__15636\,
            PADIN => \N__15635\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15628\,
            DIN => \N__15627\,
            DOUT => \N__15626\,
            PACKAGEPIN => ioFifoData(3)
        );

    \ioFifoData_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__15628\,
            PADOUT => \N__15627\,
            PADIN => \N__15626\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__15447\,
            DIN0 => \ioFifoData_in_3\,
            DOUT0 => \N__5988\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A4_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15619\,
            DIN => \N__15618\,
            DOUT => \N__15617\,
            PACKAGEPIN => \P1A4_wire\
        );

    \P1A4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__15619\,
            PADOUT => \N__15618\,
            PADIN => \N__15617\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14232\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \oRx_n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15610\,
            DIN => \N__15609\,
            DOUT => \N__15608\,
            PACKAGEPIN => \oRx_n_wire\
        );

    \oRx_n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__15610\,
            PADOUT => \N__15609\,
            PADIN => \N__15608\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14723\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15601\,
            DIN => \N__15600\,
            DOUT => \N__15599\,
            PACKAGEPIN => \P1A2_wire\
        );

    \P1A2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__15601\,
            PADOUT => \N__15600\,
            PADIN => \N__15599\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14825\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15592\,
            DIN => \N__15591\,
            DOUT => \N__15590\,
            PACKAGEPIN => ioFifoData(0)
        );

    \ioFifoData_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__15592\,
            PADOUT => \N__15591\,
            PADIN => \N__15590\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7704\,
            DIN0 => \ioFifoData_in_0\,
            DOUT0 => \N__6006\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \iRxF_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15583\,
            DIN => \N__15582\,
            DOUT => \N__15581\,
            PACKAGEPIN => \iRxF_n_wire\
        );

    \iRxF_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15583\,
            PADOUT => \N__15582\,
            PADIN => \N__15581\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \iRxF_n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15574\,
            DIN => \N__15573\,
            DOUT => \N__15572\,
            PACKAGEPIN => \P1A3_wire\
        );

    \P1A3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__15574\,
            PADOUT => \N__15573\,
            PADIN => \N__15572\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14730\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A7_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15565\,
            DIN => \N__15564\,
            DOUT => \N__15563\,
            PACKAGEPIN => \P1A7_wire\
        );

    \P1A7_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__15565\,
            PADOUT => \N__15564\,
            PADIN => \N__15563\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7779\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15556\,
            DIN => \N__15555\,
            DOUT => \N__15554\,
            PACKAGEPIN => ioFifoData(7)
        );

    \ioFifoData_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__15556\,
            PADOUT => \N__15555\,
            PADIN => \N__15554\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__12513\,
            DIN0 => \ioFifoData_in_7\,
            DOUT0 => \N__5934\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BTN_N_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15547\,
            DIN => \N__15546\,
            DOUT => \N__15545\,
            PACKAGEPIN => \BTN_N_wire\
        );

    \BTN_N_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15547\,
            PADOUT => \N__15546\,
            PADIN => \N__15545\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \BTN_N_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15538\,
            DIN => \N__15537\,
            DOUT => \N__15536\,
            PACKAGEPIN => ioFifoData(4)
        );

    \ioFifoData_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__15538\,
            PADOUT => \N__15537\,
            PADIN => \N__15536\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__13872\,
            DIN0 => \ioFifoData_in_4\,
            DOUT0 => \N__5961\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15529\,
            DIN => \N__15528\,
            DOUT => \N__15527\,
            PACKAGEPIN => ioFifoData(1)
        );

    \ioFifoData_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__15529\,
            PADOUT => \N__15528\,
            PADIN => \N__15527\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__12525\,
            DIN0 => \ioFifoData_in_1\,
            DOUT0 => \N__5919\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15520\,
            DIN => \N__15519\,
            DOUT => \N__15518\,
            PACKAGEPIN => ioFifoData(5)
        );

    \ioFifoData_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__15520\,
            PADOUT => \N__15519\,
            PADIN => \N__15518\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__12491\,
            DIN0 => \ioFifoData_in_5\,
            DOUT0 => \N__5871\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \oTx_n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15511\,
            DIN => \N__15510\,
            DOUT => \N__15509\,
            PACKAGEPIN => \oTx_n_wire\
        );

    \oTx_n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__15511\,
            PADOUT => \N__15510\,
            PADIN => \N__15509\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14225\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \iTxE_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15502\,
            DIN => \N__15501\,
            DOUT => \N__15500\,
            PACKAGEPIN => \iTxE_n_wire\
        );

    \iTxE_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15502\,
            PADOUT => \N__15501\,
            PADIN => \N__15500\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \iTxE_n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15493\,
            DIN => \N__15492\,
            DOUT => \N__15491\,
            PACKAGEPIN => \P1A1_wire\
        );

    \P1A1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__15493\,
            PADOUT => \N__15492\,
            PADIN => \N__15491\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \P1A1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15484\,
            DIN => \N__15483\,
            DOUT => \N__15482\,
            PACKAGEPIN => ioFifoData(2)
        );

    \ioFifoData_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__15484\,
            PADOUT => \N__15483\,
            PADIN => \N__15482\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__15441\,
            DIN0 => \ioFifoData_in_2\,
            DOUT0 => \N__5886\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A9_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15475\,
            DIN => \N__15474\,
            DOUT => \N__15473\,
            PACKAGEPIN => \P1A9_wire\
        );

    \P1A9_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__15475\,
            PADOUT => \N__15474\,
            PADIN => \N__15473\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__15466\,
            DIN => \N__15465\,
            DOUT => \N__15464\,
            PACKAGEPIN => ioFifoData(6)
        );

    \ioFifoData_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__15466\,
            PADOUT => \N__15465\,
            PADIN => \N__15464\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__12512\,
            DIN0 => \ioFifoData_in_6\,
            DOUT0 => \N__5901\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__3682\ : IoInMux
    port map (
            O => \N__15447\,
            I => \N__15444\
        );

    \I__3681\ : LocalMux
    port map (
            O => \N__15444\,
            I => \N_1260_i\
        );

    \I__3680\ : IoInMux
    port map (
            O => \N__15441\,
            I => \N__15438\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__15438\,
            I => \N__15435\
        );

    \I__3678\ : Odrv4
    port map (
            O => \N__15435\,
            I => \N_1259_i\
        );

    \I__3677\ : InMux
    port map (
            O => \N__15432\,
            I => \N__15429\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__15429\,
            I => \N__15426\
        );

    \I__3675\ : Odrv12
    port map (
            O => \N__15426\,
            I => \oTx_n_rep3_ess\
        );

    \I__3674\ : CascadeMux
    port map (
            O => \N__15423\,
            I => \N__15418\
        );

    \I__3673\ : CascadeMux
    port map (
            O => \N__15422\,
            I => \N__15414\
        );

    \I__3672\ : CascadeMux
    port map (
            O => \N__15421\,
            I => \N__15411\
        );

    \I__3671\ : InMux
    port map (
            O => \N__15418\,
            I => \N__15403\
        );

    \I__3670\ : InMux
    port map (
            O => \N__15417\,
            I => \N__15403\
        );

    \I__3669\ : InMux
    port map (
            O => \N__15414\,
            I => \N__15396\
        );

    \I__3668\ : InMux
    port map (
            O => \N__15411\,
            I => \N__15396\
        );

    \I__3667\ : InMux
    port map (
            O => \N__15410\,
            I => \N__15396\
        );

    \I__3666\ : CascadeMux
    port map (
            O => \N__15409\,
            I => \N__15393\
        );

    \I__3665\ : CascadeMux
    port map (
            O => \N__15408\,
            I => \N__15389\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__15403\,
            I => \N__15384\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__15396\,
            I => \N__15381\
        );

    \I__3662\ : InMux
    port map (
            O => \N__15393\,
            I => \N__15376\
        );

    \I__3661\ : InMux
    port map (
            O => \N__15392\,
            I => \N__15376\
        );

    \I__3660\ : InMux
    port map (
            O => \N__15389\,
            I => \N__15369\
        );

    \I__3659\ : InMux
    port map (
            O => \N__15388\,
            I => \N__15369\
        );

    \I__3658\ : InMux
    port map (
            O => \N__15387\,
            I => \N__15369\
        );

    \I__3657\ : Odrv4
    port map (
            O => \N__15384\,
            I => \fifo_inst.ftdi_output_inst.rWrDelayZ0\
        );

    \I__3656\ : Odrv4
    port map (
            O => \N__15381\,
            I => \fifo_inst.ftdi_output_inst.rWrDelayZ0\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__15376\,
            I => \fifo_inst.ftdi_output_inst.rWrDelayZ0\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__15369\,
            I => \fifo_inst.ftdi_output_inst.rWrDelayZ0\
        );

    \I__3653\ : InMux
    port map (
            O => \N__15360\,
            I => \N__15351\
        );

    \I__3652\ : InMux
    port map (
            O => \N__15359\,
            I => \N__15351\
        );

    \I__3651\ : InMux
    port map (
            O => \N__15358\,
            I => \N__15344\
        );

    \I__3650\ : InMux
    port map (
            O => \N__15357\,
            I => \N__15344\
        );

    \I__3649\ : InMux
    port map (
            O => \N__15356\,
            I => \N__15344\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__15351\,
            I => \N__15336\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__15344\,
            I => \N__15333\
        );

    \I__3646\ : InMux
    port map (
            O => \N__15343\,
            I => \N__15328\
        );

    \I__3645\ : InMux
    port map (
            O => \N__15342\,
            I => \N__15328\
        );

    \I__3644\ : InMux
    port map (
            O => \N__15341\,
            I => \N__15321\
        );

    \I__3643\ : InMux
    port map (
            O => \N__15340\,
            I => \N__15321\
        );

    \I__3642\ : InMux
    port map (
            O => \N__15339\,
            I => \N__15321\
        );

    \I__3641\ : Odrv4
    port map (
            O => \N__15336\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4\
        );

    \I__3640\ : Odrv4
    port map (
            O => \N__15333\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4\
        );

    \I__3639\ : LocalMux
    port map (
            O => \N__15328\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__15321\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4\
        );

    \I__3637\ : InMux
    port map (
            O => \N__15312\,
            I => \N__15309\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__15309\,
            I => \N__15306\
        );

    \I__3635\ : Odrv4
    port map (
            O => \N__15306\,
            I => \oTx_n_rep2_ess\
        );

    \I__3634\ : CEMux
    port map (
            O => \N__15303\,
            I => \N__15299\
        );

    \I__3633\ : CEMux
    port map (
            O => \N__15302\,
            I => \N__15296\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__15299\,
            I => \fifo_inst.ftdi_output_inst.N_88_i_0\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__15296\,
            I => \fifo_inst.ftdi_output_inst.N_88_i_0\
        );

    \I__3630\ : CascadeMux
    port map (
            O => \N__15291\,
            I => \N__15287\
        );

    \I__3629\ : InMux
    port map (
            O => \N__15290\,
            I => \N__15275\
        );

    \I__3628\ : InMux
    port map (
            O => \N__15287\,
            I => \N__15266\
        );

    \I__3627\ : InMux
    port map (
            O => \N__15286\,
            I => \N__15266\
        );

    \I__3626\ : InMux
    port map (
            O => \N__15285\,
            I => \N__15266\
        );

    \I__3625\ : InMux
    port map (
            O => \N__15284\,
            I => \N__15266\
        );

    \I__3624\ : InMux
    port map (
            O => \N__15283\,
            I => \N__15263\
        );

    \I__3623\ : InMux
    port map (
            O => \N__15282\,
            I => \N__15260\
        );

    \I__3622\ : InMux
    port map (
            O => \N__15281\,
            I => \N__15253\
        );

    \I__3621\ : InMux
    port map (
            O => \N__15280\,
            I => \N__15253\
        );

    \I__3620\ : InMux
    port map (
            O => \N__15279\,
            I => \N__15253\
        );

    \I__3619\ : InMux
    port map (
            O => \N__15278\,
            I => \N__15250\
        );

    \I__3618\ : LocalMux
    port map (
            O => \N__15275\,
            I => \N__15245\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__15266\,
            I => \N__15242\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__15263\,
            I => \N__15237\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__15260\,
            I => \N__15233\
        );

    \I__3614\ : LocalMux
    port map (
            O => \N__15253\,
            I => \N__15226\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__15250\,
            I => \N__15220\
        );

    \I__3612\ : SRMux
    port map (
            O => \N__15249\,
            I => \N__15177\
        );

    \I__3611\ : SRMux
    port map (
            O => \N__15248\,
            I => \N__15177\
        );

    \I__3610\ : Glb2LocalMux
    port map (
            O => \N__15245\,
            I => \N__15177\
        );

    \I__3609\ : Glb2LocalMux
    port map (
            O => \N__15242\,
            I => \N__15177\
        );

    \I__3608\ : SRMux
    port map (
            O => \N__15241\,
            I => \N__15177\
        );

    \I__3607\ : SRMux
    port map (
            O => \N__15240\,
            I => \N__15177\
        );

    \I__3606\ : Glb2LocalMux
    port map (
            O => \N__15237\,
            I => \N__15177\
        );

    \I__3605\ : SRMux
    port map (
            O => \N__15236\,
            I => \N__15177\
        );

    \I__3604\ : Glb2LocalMux
    port map (
            O => \N__15233\,
            I => \N__15177\
        );

    \I__3603\ : SRMux
    port map (
            O => \N__15232\,
            I => \N__15177\
        );

    \I__3602\ : SRMux
    port map (
            O => \N__15231\,
            I => \N__15177\
        );

    \I__3601\ : SRMux
    port map (
            O => \N__15230\,
            I => \N__15177\
        );

    \I__3600\ : SRMux
    port map (
            O => \N__15229\,
            I => \N__15177\
        );

    \I__3599\ : Glb2LocalMux
    port map (
            O => \N__15226\,
            I => \N__15177\
        );

    \I__3598\ : SRMux
    port map (
            O => \N__15225\,
            I => \N__15177\
        );

    \I__3597\ : SRMux
    port map (
            O => \N__15224\,
            I => \N__15177\
        );

    \I__3596\ : SRMux
    port map (
            O => \N__15223\,
            I => \N__15177\
        );

    \I__3595\ : Glb2LocalMux
    port map (
            O => \N__15220\,
            I => \N__15177\
        );

    \I__3594\ : SRMux
    port map (
            O => \N__15219\,
            I => \N__15177\
        );

    \I__3593\ : SRMux
    port map (
            O => \N__15218\,
            I => \N__15177\
        );

    \I__3592\ : GlobalMux
    port map (
            O => \N__15177\,
            I => \N__15174\
        );

    \I__3591\ : gio2CtrlBuf
    port map (
            O => \N__15174\,
            I => \wPllLocked_iso_i_g\
        );

    \I__3590\ : InMux
    port map (
            O => \N__15171\,
            I => \N__15168\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__15168\,
            I => \N__15163\
        );

    \I__3588\ : InMux
    port map (
            O => \N__15167\,
            I => \N__15160\
        );

    \I__3587\ : InMux
    port map (
            O => \N__15166\,
            I => \N__15157\
        );

    \I__3586\ : Span4Mux_h
    port map (
            O => \N__15163\,
            I => \N__15154\
        );

    \I__3585\ : LocalMux
    port map (
            O => \N__15160\,
            I => \N__15151\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__15157\,
            I => \N__15148\
        );

    \I__3583\ : Span4Mux_h
    port map (
            O => \N__15154\,
            I => \N__15143\
        );

    \I__3582\ : Span4Mux_v
    port map (
            O => \N__15151\,
            I => \N__15140\
        );

    \I__3581\ : Span4Mux_h
    port map (
            O => \N__15148\,
            I => \N__15137\
        );

    \I__3580\ : InMux
    port map (
            O => \N__15147\,
            I => \N__15134\
        );

    \I__3579\ : InMux
    port map (
            O => \N__15146\,
            I => \N__15131\
        );

    \I__3578\ : Odrv4
    port map (
            O => \N__15143\,
            I => \DUT.wRxByte_2\
        );

    \I__3577\ : Odrv4
    port map (
            O => \N__15140\,
            I => \DUT.wRxByte_2\
        );

    \I__3576\ : Odrv4
    port map (
            O => \N__15137\,
            I => \DUT.wRxByte_2\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__15134\,
            I => \DUT.wRxByte_2\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__15131\,
            I => \DUT.wRxByte_2\
        );

    \I__3573\ : InMux
    port map (
            O => \N__15120\,
            I => \N__15117\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__15117\,
            I => \N__15114\
        );

    \I__3571\ : Odrv12
    port map (
            O => \N__15114\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_2\
        );

    \I__3570\ : InMux
    port map (
            O => \N__15111\,
            I => \N__15107\
        );

    \I__3569\ : InMux
    port map (
            O => \N__15110\,
            I => \N__15103\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__15107\,
            I => \N__15100\
        );

    \I__3567\ : InMux
    port map (
            O => \N__15106\,
            I => \N__15097\
        );

    \I__3566\ : LocalMux
    port map (
            O => \N__15103\,
            I => \N__15094\
        );

    \I__3565\ : Span4Mux_v
    port map (
            O => \N__15100\,
            I => \N__15089\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__15097\,
            I => \N__15089\
        );

    \I__3563\ : Span4Mux_v
    port map (
            O => \N__15094\,
            I => \N__15086\
        );

    \I__3562\ : Sp12to4
    port map (
            O => \N__15089\,
            I => \N__15083\
        );

    \I__3561\ : Sp12to4
    port map (
            O => \N__15086\,
            I => \N__15076\
        );

    \I__3560\ : Span12Mux_s6_v
    port map (
            O => \N__15083\,
            I => \N__15076\
        );

    \I__3559\ : InMux
    port map (
            O => \N__15082\,
            I => \N__15073\
        );

    \I__3558\ : InMux
    port map (
            O => \N__15081\,
            I => \N__15070\
        );

    \I__3557\ : Odrv12
    port map (
            O => \N__15076\,
            I => \DUT.wRxByte_5\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__15073\,
            I => \DUT.wRxByte_5\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__15070\,
            I => \DUT.wRxByte_5\
        );

    \I__3554\ : InMux
    port map (
            O => \N__15063\,
            I => \N__15060\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__15060\,
            I => \N__15057\
        );

    \I__3552\ : Odrv12
    port map (
            O => \N__15057\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_5\
        );

    \I__3551\ : ClkMux
    port map (
            O => \N__15054\,
            I => \N__14871\
        );

    \I__3550\ : ClkMux
    port map (
            O => \N__15053\,
            I => \N__14871\
        );

    \I__3549\ : ClkMux
    port map (
            O => \N__15052\,
            I => \N__14871\
        );

    \I__3548\ : ClkMux
    port map (
            O => \N__15051\,
            I => \N__14871\
        );

    \I__3547\ : ClkMux
    port map (
            O => \N__15050\,
            I => \N__14871\
        );

    \I__3546\ : ClkMux
    port map (
            O => \N__15049\,
            I => \N__14871\
        );

    \I__3545\ : ClkMux
    port map (
            O => \N__15048\,
            I => \N__14871\
        );

    \I__3544\ : ClkMux
    port map (
            O => \N__15047\,
            I => \N__14871\
        );

    \I__3543\ : ClkMux
    port map (
            O => \N__15046\,
            I => \N__14871\
        );

    \I__3542\ : ClkMux
    port map (
            O => \N__15045\,
            I => \N__14871\
        );

    \I__3541\ : ClkMux
    port map (
            O => \N__15044\,
            I => \N__14871\
        );

    \I__3540\ : ClkMux
    port map (
            O => \N__15043\,
            I => \N__14871\
        );

    \I__3539\ : ClkMux
    port map (
            O => \N__15042\,
            I => \N__14871\
        );

    \I__3538\ : ClkMux
    port map (
            O => \N__15041\,
            I => \N__14871\
        );

    \I__3537\ : ClkMux
    port map (
            O => \N__15040\,
            I => \N__14871\
        );

    \I__3536\ : ClkMux
    port map (
            O => \N__15039\,
            I => \N__14871\
        );

    \I__3535\ : ClkMux
    port map (
            O => \N__15038\,
            I => \N__14871\
        );

    \I__3534\ : ClkMux
    port map (
            O => \N__15037\,
            I => \N__14871\
        );

    \I__3533\ : ClkMux
    port map (
            O => \N__15036\,
            I => \N__14871\
        );

    \I__3532\ : ClkMux
    port map (
            O => \N__15035\,
            I => \N__14871\
        );

    \I__3531\ : ClkMux
    port map (
            O => \N__15034\,
            I => \N__14871\
        );

    \I__3530\ : ClkMux
    port map (
            O => \N__15033\,
            I => \N__14871\
        );

    \I__3529\ : ClkMux
    port map (
            O => \N__15032\,
            I => \N__14871\
        );

    \I__3528\ : ClkMux
    port map (
            O => \N__15031\,
            I => \N__14871\
        );

    \I__3527\ : ClkMux
    port map (
            O => \N__15030\,
            I => \N__14871\
        );

    \I__3526\ : ClkMux
    port map (
            O => \N__15029\,
            I => \N__14871\
        );

    \I__3525\ : ClkMux
    port map (
            O => \N__15028\,
            I => \N__14871\
        );

    \I__3524\ : ClkMux
    port map (
            O => \N__15027\,
            I => \N__14871\
        );

    \I__3523\ : ClkMux
    port map (
            O => \N__15026\,
            I => \N__14871\
        );

    \I__3522\ : ClkMux
    port map (
            O => \N__15025\,
            I => \N__14871\
        );

    \I__3521\ : ClkMux
    port map (
            O => \N__15024\,
            I => \N__14871\
        );

    \I__3520\ : ClkMux
    port map (
            O => \N__15023\,
            I => \N__14871\
        );

    \I__3519\ : ClkMux
    port map (
            O => \N__15022\,
            I => \N__14871\
        );

    \I__3518\ : ClkMux
    port map (
            O => \N__15021\,
            I => \N__14871\
        );

    \I__3517\ : ClkMux
    port map (
            O => \N__15020\,
            I => \N__14871\
        );

    \I__3516\ : ClkMux
    port map (
            O => \N__15019\,
            I => \N__14871\
        );

    \I__3515\ : ClkMux
    port map (
            O => \N__15018\,
            I => \N__14871\
        );

    \I__3514\ : ClkMux
    port map (
            O => \N__15017\,
            I => \N__14871\
        );

    \I__3513\ : ClkMux
    port map (
            O => \N__15016\,
            I => \N__14871\
        );

    \I__3512\ : ClkMux
    port map (
            O => \N__15015\,
            I => \N__14871\
        );

    \I__3511\ : ClkMux
    port map (
            O => \N__15014\,
            I => \N__14871\
        );

    \I__3510\ : ClkMux
    port map (
            O => \N__15013\,
            I => \N__14871\
        );

    \I__3509\ : ClkMux
    port map (
            O => \N__15012\,
            I => \N__14871\
        );

    \I__3508\ : ClkMux
    port map (
            O => \N__15011\,
            I => \N__14871\
        );

    \I__3507\ : ClkMux
    port map (
            O => \N__15010\,
            I => \N__14871\
        );

    \I__3506\ : ClkMux
    port map (
            O => \N__15009\,
            I => \N__14871\
        );

    \I__3505\ : ClkMux
    port map (
            O => \N__15008\,
            I => \N__14871\
        );

    \I__3504\ : ClkMux
    port map (
            O => \N__15007\,
            I => \N__14871\
        );

    \I__3503\ : ClkMux
    port map (
            O => \N__15006\,
            I => \N__14871\
        );

    \I__3502\ : ClkMux
    port map (
            O => \N__15005\,
            I => \N__14871\
        );

    \I__3501\ : ClkMux
    port map (
            O => \N__15004\,
            I => \N__14871\
        );

    \I__3500\ : ClkMux
    port map (
            O => \N__15003\,
            I => \N__14871\
        );

    \I__3499\ : ClkMux
    port map (
            O => \N__15002\,
            I => \N__14871\
        );

    \I__3498\ : ClkMux
    port map (
            O => \N__15001\,
            I => \N__14871\
        );

    \I__3497\ : ClkMux
    port map (
            O => \N__15000\,
            I => \N__14871\
        );

    \I__3496\ : ClkMux
    port map (
            O => \N__14999\,
            I => \N__14871\
        );

    \I__3495\ : ClkMux
    port map (
            O => \N__14998\,
            I => \N__14871\
        );

    \I__3494\ : ClkMux
    port map (
            O => \N__14997\,
            I => \N__14871\
        );

    \I__3493\ : ClkMux
    port map (
            O => \N__14996\,
            I => \N__14871\
        );

    \I__3492\ : ClkMux
    port map (
            O => \N__14995\,
            I => \N__14871\
        );

    \I__3491\ : ClkMux
    port map (
            O => \N__14994\,
            I => \N__14871\
        );

    \I__3490\ : GlobalMux
    port map (
            O => \N__14871\,
            I => clk_48mhz
        );

    \I__3489\ : CEMux
    port map (
            O => \N__14868\,
            I => \N__14863\
        );

    \I__3488\ : CEMux
    port map (
            O => \N__14867\,
            I => \N__14860\
        );

    \I__3487\ : CEMux
    port map (
            O => \N__14866\,
            I => \N__14856\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__14863\,
            I => \N__14853\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__14860\,
            I => \N__14850\
        );

    \I__3484\ : CEMux
    port map (
            O => \N__14859\,
            I => \N__14847\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__14856\,
            I => \N__14844\
        );

    \I__3482\ : Span4Mux_h
    port map (
            O => \N__14853\,
            I => \N__14839\
        );

    \I__3481\ : Span4Mux_h
    port map (
            O => \N__14850\,
            I => \N__14839\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__14847\,
            I => \N__14836\
        );

    \I__3479\ : Span4Mux_v
    port map (
            O => \N__14844\,
            I => \N__14833\
        );

    \I__3478\ : Odrv4
    port map (
            O => \N__14839\,
            I => \DUT.fifo_rx_inst.rFifoData_awe0\
        );

    \I__3477\ : Odrv4
    port map (
            O => \N__14836\,
            I => \DUT.fifo_rx_inst.rFifoData_awe0\
        );

    \I__3476\ : Odrv4
    port map (
            O => \N__14833\,
            I => \DUT.fifo_rx_inst.rFifoData_awe0\
        );

    \I__3475\ : CascadeMux
    port map (
            O => \N__14826\,
            I => \N__14820\
        );

    \I__3474\ : IoInMux
    port map (
            O => \N__14825\,
            I => \N__14809\
        );

    \I__3473\ : InMux
    port map (
            O => \N__14824\,
            I => \N__14806\
        );

    \I__3472\ : InMux
    port map (
            O => \N__14823\,
            I => \N__14789\
        );

    \I__3471\ : InMux
    port map (
            O => \N__14820\,
            I => \N__14789\
        );

    \I__3470\ : InMux
    port map (
            O => \N__14819\,
            I => \N__14789\
        );

    \I__3469\ : InMux
    port map (
            O => \N__14818\,
            I => \N__14789\
        );

    \I__3468\ : InMux
    port map (
            O => \N__14817\,
            I => \N__14789\
        );

    \I__3467\ : InMux
    port map (
            O => \N__14816\,
            I => \N__14789\
        );

    \I__3466\ : InMux
    port map (
            O => \N__14815\,
            I => \N__14789\
        );

    \I__3465\ : InMux
    port map (
            O => \N__14814\,
            I => \N__14789\
        );

    \I__3464\ : InMux
    port map (
            O => \N__14813\,
            I => \N__14786\
        );

    \I__3463\ : InMux
    port map (
            O => \N__14812\,
            I => \N__14783\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__14809\,
            I => \N__14780\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__14806\,
            I => \N__14777\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__14789\,
            I => \N__14774\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__14786\,
            I => \N__14770\
        );

    \I__3458\ : LocalMux
    port map (
            O => \N__14783\,
            I => \N__14767\
        );

    \I__3457\ : Span12Mux_s1_v
    port map (
            O => \N__14780\,
            I => \N__14764\
        );

    \I__3456\ : Span4Mux_h
    port map (
            O => \N__14777\,
            I => \N__14761\
        );

    \I__3455\ : Span4Mux_v
    port map (
            O => \N__14774\,
            I => \N__14758\
        );

    \I__3454\ : InMux
    port map (
            O => \N__14773\,
            I => \N__14755\
        );

    \I__3453\ : Span4Mux_h
    port map (
            O => \N__14770\,
            I => \N__14750\
        );

    \I__3452\ : Span4Mux_h
    port map (
            O => \N__14767\,
            I => \N__14750\
        );

    \I__3451\ : Span12Mux_h
    port map (
            O => \N__14764\,
            I => \N__14747\
        );

    \I__3450\ : Span4Mux_h
    port map (
            O => \N__14761\,
            I => \N__14744\
        );

    \I__3449\ : Span4Mux_h
    port map (
            O => \N__14758\,
            I => \N__14737\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__14755\,
            I => \N__14737\
        );

    \I__3447\ : Span4Mux_v
    port map (
            O => \N__14750\,
            I => \N__14737\
        );

    \I__3446\ : Odrv12
    port map (
            O => \N__14747\,
            I => \P1A2_c\
        );

    \I__3445\ : Odrv4
    port map (
            O => \N__14744\,
            I => \P1A2_c\
        );

    \I__3444\ : Odrv4
    port map (
            O => \N__14737\,
            I => \P1A2_c\
        );

    \I__3443\ : IoInMux
    port map (
            O => \N__14730\,
            I => \N__14727\
        );

    \I__3442\ : LocalMux
    port map (
            O => \N__14727\,
            I => \N__14724\
        );

    \I__3441\ : IoSpan4Mux
    port map (
            O => \N__14724\,
            I => \N__14720\
        );

    \I__3440\ : IoInMux
    port map (
            O => \N__14723\,
            I => \N__14717\
        );

    \I__3439\ : Sp12to4
    port map (
            O => \N__14720\,
            I => \N__14714\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__14717\,
            I => \N__14711\
        );

    \I__3437\ : Span12Mux_s7_v
    port map (
            O => \N__14714\,
            I => \N__14707\
        );

    \I__3436\ : Span12Mux_s7_v
    port map (
            O => \N__14711\,
            I => \N__14704\
        );

    \I__3435\ : InMux
    port map (
            O => \N__14710\,
            I => \N__14701\
        );

    \I__3434\ : Odrv12
    port map (
            O => \N__14707\,
            I => \P1A3_c\
        );

    \I__3433\ : Odrv12
    port map (
            O => \N__14704\,
            I => \P1A3_c\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__14701\,
            I => \P1A3_c\
        );

    \I__3431\ : InMux
    port map (
            O => \N__14694\,
            I => \N__14687\
        );

    \I__3430\ : InMux
    port map (
            O => \N__14693\,
            I => \N__14687\
        );

    \I__3429\ : InMux
    port map (
            O => \N__14692\,
            I => \N__14684\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__14687\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1\
        );

    \I__3427\ : LocalMux
    port map (
            O => \N__14684\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1\
        );

    \I__3426\ : CascadeMux
    port map (
            O => \N__14679\,
            I => \N__14676\
        );

    \I__3425\ : InMux
    port map (
            O => \N__14676\,
            I => \N__14673\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__14673\,
            I => \N__14670\
        );

    \I__3423\ : Span4Mux_v
    port map (
            O => \N__14670\,
            I => \N__14666\
        );

    \I__3422\ : InMux
    port map (
            O => \N__14669\,
            I => \N__14663\
        );

    \I__3421\ : Sp12to4
    port map (
            O => \N__14666\,
            I => \N__14658\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__14663\,
            I => \N__14658\
        );

    \I__3419\ : Span12Mux_s7_h
    port map (
            O => \N__14658\,
            I => \N__14655\
        );

    \I__3418\ : Span12Mux_v
    port map (
            O => \N__14655\,
            I => \N__14652\
        );

    \I__3417\ : Odrv12
    port map (
            O => \N__14652\,
            I => \iTxE_n_c\
        );

    \I__3416\ : CascadeMux
    port map (
            O => \N__14649\,
            I => \N__14644\
        );

    \I__3415\ : InMux
    port map (
            O => \N__14648\,
            I => \N__14637\
        );

    \I__3414\ : InMux
    port map (
            O => \N__14647\,
            I => \N__14637\
        );

    \I__3413\ : InMux
    port map (
            O => \N__14644\,
            I => \N__14637\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__14637\,
            I => \N__14633\
        );

    \I__3411\ : InMux
    port map (
            O => \N__14636\,
            I => \N__14630\
        );

    \I__3410\ : Span4Mux_v
    port map (
            O => \N__14633\,
            I => \N__14627\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__14630\,
            I => \N__14624\
        );

    \I__3408\ : Sp12to4
    port map (
            O => \N__14627\,
            I => \N__14621\
        );

    \I__3407\ : Span4Mux_h
    port map (
            O => \N__14624\,
            I => \N__14618\
        );

    \I__3406\ : Span12Mux_s7_h
    port map (
            O => \N__14621\,
            I => \N__14613\
        );

    \I__3405\ : Sp12to4
    port map (
            O => \N__14618\,
            I => \N__14613\
        );

    \I__3404\ : Span12Mux_v
    port map (
            O => \N__14613\,
            I => \N__14610\
        );

    \I__3403\ : Odrv12
    port map (
            O => \N__14610\,
            I => \iRxF_n_c\
        );

    \I__3402\ : CascadeMux
    port map (
            O => \N__14607\,
            I => \N__14604\
        );

    \I__3401\ : InMux
    port map (
            O => \N__14604\,
            I => \N__14600\
        );

    \I__3400\ : InMux
    port map (
            O => \N__14603\,
            I => \N__14597\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__14600\,
            I => \N__14592\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__14597\,
            I => \N__14592\
        );

    \I__3397\ : Span4Mux_v
    port map (
            O => \N__14592\,
            I => \N__14589\
        );

    \I__3396\ : Span4Mux_h
    port map (
            O => \N__14589\,
            I => \N__14585\
        );

    \I__3395\ : InMux
    port map (
            O => \N__14588\,
            I => \N__14582\
        );

    \I__3394\ : Odrv4
    port map (
            O => \N__14585\,
            I => \G_120\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__14582\,
            I => \G_120\
        );

    \I__3392\ : CascadeMux
    port map (
            O => \N__14577\,
            I => \N__14568\
        );

    \I__3391\ : CascadeMux
    port map (
            O => \N__14576\,
            I => \N__14558\
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__14575\,
            I => \N__14553\
        );

    \I__3389\ : InMux
    port map (
            O => \N__14574\,
            I => \N__14543\
        );

    \I__3388\ : InMux
    port map (
            O => \N__14573\,
            I => \N__14540\
        );

    \I__3387\ : InMux
    port map (
            O => \N__14572\,
            I => \N__14537\
        );

    \I__3386\ : InMux
    port map (
            O => \N__14571\,
            I => \N__14530\
        );

    \I__3385\ : InMux
    port map (
            O => \N__14568\,
            I => \N__14530\
        );

    \I__3384\ : InMux
    port map (
            O => \N__14567\,
            I => \N__14530\
        );

    \I__3383\ : InMux
    port map (
            O => \N__14566\,
            I => \N__14527\
        );

    \I__3382\ : InMux
    port map (
            O => \N__14565\,
            I => \N__14522\
        );

    \I__3381\ : InMux
    port map (
            O => \N__14564\,
            I => \N__14522\
        );

    \I__3380\ : InMux
    port map (
            O => \N__14563\,
            I => \N__14517\
        );

    \I__3379\ : InMux
    port map (
            O => \N__14562\,
            I => \N__14517\
        );

    \I__3378\ : InMux
    port map (
            O => \N__14561\,
            I => \N__14514\
        );

    \I__3377\ : InMux
    port map (
            O => \N__14558\,
            I => \N__14511\
        );

    \I__3376\ : InMux
    port map (
            O => \N__14557\,
            I => \N__14508\
        );

    \I__3375\ : InMux
    port map (
            O => \N__14556\,
            I => \N__14505\
        );

    \I__3374\ : InMux
    port map (
            O => \N__14553\,
            I => \N__14502\
        );

    \I__3373\ : InMux
    port map (
            O => \N__14552\,
            I => \N__14497\
        );

    \I__3372\ : InMux
    port map (
            O => \N__14551\,
            I => \N__14497\
        );

    \I__3371\ : InMux
    port map (
            O => \N__14550\,
            I => \N__14492\
        );

    \I__3370\ : InMux
    port map (
            O => \N__14549\,
            I => \N__14492\
        );

    \I__3369\ : InMux
    port map (
            O => \N__14548\,
            I => \N__14489\
        );

    \I__3368\ : InMux
    port map (
            O => \N__14547\,
            I => \N__14486\
        );

    \I__3367\ : InMux
    port map (
            O => \N__14546\,
            I => \N__14483\
        );

    \I__3366\ : LocalMux
    port map (
            O => \N__14543\,
            I => \N__14480\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__14540\,
            I => \N__14477\
        );

    \I__3364\ : LocalMux
    port map (
            O => \N__14537\,
            I => \N__14474\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__14530\,
            I => \N__14471\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__14527\,
            I => \N__14468\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__14522\,
            I => \N__14465\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__14517\,
            I => \N__14462\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__14514\,
            I => \N__14457\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__14511\,
            I => \N__14453\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__14508\,
            I => \N__14447\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__14505\,
            I => \N__14444\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__14502\,
            I => \N__14440\
        );

    \I__3354\ : LocalMux
    port map (
            O => \N__14497\,
            I => \N__14437\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__14492\,
            I => \N__14432\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__14489\,
            I => \N__14429\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__14486\,
            I => \N__14425\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__14483\,
            I => \N__14422\
        );

    \I__3349\ : Glb2LocalMux
    port map (
            O => \N__14480\,
            I => \N__14364\
        );

    \I__3348\ : Glb2LocalMux
    port map (
            O => \N__14477\,
            I => \N__14364\
        );

    \I__3347\ : Glb2LocalMux
    port map (
            O => \N__14474\,
            I => \N__14364\
        );

    \I__3346\ : Glb2LocalMux
    port map (
            O => \N__14471\,
            I => \N__14364\
        );

    \I__3345\ : Glb2LocalMux
    port map (
            O => \N__14468\,
            I => \N__14364\
        );

    \I__3344\ : Glb2LocalMux
    port map (
            O => \N__14465\,
            I => \N__14364\
        );

    \I__3343\ : Glb2LocalMux
    port map (
            O => \N__14462\,
            I => \N__14364\
        );

    \I__3342\ : CEMux
    port map (
            O => \N__14461\,
            I => \N__14364\
        );

    \I__3341\ : CEMux
    port map (
            O => \N__14460\,
            I => \N__14364\
        );

    \I__3340\ : Glb2LocalMux
    port map (
            O => \N__14457\,
            I => \N__14364\
        );

    \I__3339\ : CEMux
    port map (
            O => \N__14456\,
            I => \N__14364\
        );

    \I__3338\ : Glb2LocalMux
    port map (
            O => \N__14453\,
            I => \N__14364\
        );

    \I__3337\ : CEMux
    port map (
            O => \N__14452\,
            I => \N__14364\
        );

    \I__3336\ : CEMux
    port map (
            O => \N__14451\,
            I => \N__14364\
        );

    \I__3335\ : CEMux
    port map (
            O => \N__14450\,
            I => \N__14364\
        );

    \I__3334\ : Glb2LocalMux
    port map (
            O => \N__14447\,
            I => \N__14364\
        );

    \I__3333\ : Glb2LocalMux
    port map (
            O => \N__14444\,
            I => \N__14364\
        );

    \I__3332\ : CEMux
    port map (
            O => \N__14443\,
            I => \N__14364\
        );

    \I__3331\ : Glb2LocalMux
    port map (
            O => \N__14440\,
            I => \N__14364\
        );

    \I__3330\ : Glb2LocalMux
    port map (
            O => \N__14437\,
            I => \N__14364\
        );

    \I__3329\ : CEMux
    port map (
            O => \N__14436\,
            I => \N__14364\
        );

    \I__3328\ : CEMux
    port map (
            O => \N__14435\,
            I => \N__14364\
        );

    \I__3327\ : Glb2LocalMux
    port map (
            O => \N__14432\,
            I => \N__14364\
        );

    \I__3326\ : Glb2LocalMux
    port map (
            O => \N__14429\,
            I => \N__14364\
        );

    \I__3325\ : CEMux
    port map (
            O => \N__14428\,
            I => \N__14364\
        );

    \I__3324\ : Glb2LocalMux
    port map (
            O => \N__14425\,
            I => \N__14364\
        );

    \I__3323\ : Glb2LocalMux
    port map (
            O => \N__14422\,
            I => \N__14364\
        );

    \I__3322\ : CEMux
    port map (
            O => \N__14421\,
            I => \N__14364\
        );

    \I__3321\ : GlobalMux
    port map (
            O => \N__14364\,
            I => \N__14361\
        );

    \I__3320\ : gio2CtrlBuf
    port map (
            O => \N__14361\,
            I => \wPllLocked_g\
        );

    \I__3319\ : InMux
    port map (
            O => \N__14358\,
            I => \N__14353\
        );

    \I__3318\ : InMux
    port map (
            O => \N__14357\,
            I => \N__14348\
        );

    \I__3317\ : InMux
    port map (
            O => \N__14356\,
            I => \N__14348\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__14353\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__14348\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2\
        );

    \I__3314\ : CascadeMux
    port map (
            O => \N__14343\,
            I => \fifo_inst.ftdi_output_inst.N_87_cascade_\
        );

    \I__3313\ : InMux
    port map (
            O => \N__14340\,
            I => \N__14337\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__14337\,
            I => \N__14333\
        );

    \I__3311\ : InMux
    port map (
            O => \N__14336\,
            I => \N__14330\
        );

    \I__3310\ : Odrv4
    port map (
            O => \N__14333\,
            I => \fifo_inst.ftdi_output_inst.N_77_0\
        );

    \I__3309\ : LocalMux
    port map (
            O => \N__14330\,
            I => \fifo_inst.ftdi_output_inst.N_77_0\
        );

    \I__3308\ : InMux
    port map (
            O => \N__14325\,
            I => \N__14315\
        );

    \I__3307\ : InMux
    port map (
            O => \N__14324\,
            I => \N__14315\
        );

    \I__3306\ : InMux
    port map (
            O => \N__14323\,
            I => \N__14315\
        );

    \I__3305\ : InMux
    port map (
            O => \N__14322\,
            I => \N__14312\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__14315\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__14312\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0\
        );

    \I__3302\ : InMux
    port map (
            O => \N__14307\,
            I => \N__14304\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__14304\,
            I => \N__14301\
        );

    \I__3300\ : Span4Mux_v
    port map (
            O => \N__14301\,
            I => \N__14298\
        );

    \I__3299\ : Sp12to4
    port map (
            O => \N__14298\,
            I => \N__14295\
        );

    \I__3298\ : Span12Mux_s6_h
    port map (
            O => \N__14295\,
            I => \N__14292\
        );

    \I__3297\ : Span12Mux_v
    port map (
            O => \N__14292\,
            I => \N__14289\
        );

    \I__3296\ : Odrv12
    port map (
            O => \N__14289\,
            I => \ioFifoData_in_7\
        );

    \I__3295\ : CascadeMux
    port map (
            O => \N__14286\,
            I => \N__14283\
        );

    \I__3294\ : InMux
    port map (
            O => \N__14283\,
            I => \N__14280\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__14280\,
            I => \N__14277\
        );

    \I__3292\ : Span4Mux_v
    port map (
            O => \N__14277\,
            I => \N__14274\
        );

    \I__3291\ : Span4Mux_h
    port map (
            O => \N__14274\,
            I => \N__14271\
        );

    \I__3290\ : Odrv4
    port map (
            O => \N__14271\,
            I => \wRxFifoData_7\
        );

    \I__3289\ : CEMux
    port map (
            O => \N__14268\,
            I => \N__14263\
        );

    \I__3288\ : CEMux
    port map (
            O => \N__14267\,
            I => \N__14260\
        );

    \I__3287\ : CEMux
    port map (
            O => \N__14266\,
            I => \N__14257\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__14263\,
            I => \N__14254\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__14260\,
            I => \N__14251\
        );

    \I__3284\ : LocalMux
    port map (
            O => \N__14257\,
            I => \N__14248\
        );

    \I__3283\ : Span4Mux_h
    port map (
            O => \N__14254\,
            I => \N__14245\
        );

    \I__3282\ : Span4Mux_h
    port map (
            O => \N__14251\,
            I => \N__14240\
        );

    \I__3281\ : Span4Mux_h
    port map (
            O => \N__14248\,
            I => \N__14240\
        );

    \I__3280\ : Odrv4
    port map (
            O => \N__14245\,
            I => \fifo_inst.ftdi_output_inst.rFifoState_0_1\
        );

    \I__3279\ : Odrv4
    port map (
            O => \N__14240\,
            I => \fifo_inst.ftdi_output_inst.rFifoState_0_1\
        );

    \I__3278\ : CascadeMux
    port map (
            O => \N__14235\,
            I => \fifo_inst.ftdi_output_inst.N_77_0_cascade_\
        );

    \I__3277\ : IoInMux
    port map (
            O => \N__14232\,
            I => \N__14229\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__14229\,
            I => \N__14226\
        );

    \I__3275\ : IoSpan4Mux
    port map (
            O => \N__14226\,
            I => \N__14222\
        );

    \I__3274\ : IoInMux
    port map (
            O => \N__14225\,
            I => \N__14219\
        );

    \I__3273\ : Span4Mux_s2_v
    port map (
            O => \N__14222\,
            I => \N__14216\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__14219\,
            I => \N__14212\
        );

    \I__3271\ : Span4Mux_h
    port map (
            O => \N__14216\,
            I => \N__14209\
        );

    \I__3270\ : InMux
    port map (
            O => \N__14215\,
            I => \N__14206\
        );

    \I__3269\ : Span12Mux_s11_v
    port map (
            O => \N__14212\,
            I => \N__14203\
        );

    \I__3268\ : Span4Mux_h
    port map (
            O => \N__14209\,
            I => \N__14198\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__14206\,
            I => \N__14198\
        );

    \I__3266\ : Span12Mux_v
    port map (
            O => \N__14203\,
            I => \N__14194\
        );

    \I__3265\ : Span4Mux_h
    port map (
            O => \N__14198\,
            I => \N__14191\
        );

    \I__3264\ : InMux
    port map (
            O => \N__14197\,
            I => \N__14188\
        );

    \I__3263\ : Odrv12
    port map (
            O => \N__14194\,
            I => \P1A4_c\
        );

    \I__3262\ : Odrv4
    port map (
            O => \N__14191\,
            I => \P1A4_c\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__14188\,
            I => \P1A4_c\
        );

    \I__3260\ : CascadeMux
    port map (
            O => \N__14181\,
            I => \fifo_inst.ftdi_output_inst.oPacketRead_1_sqmuxa_1_cascade_\
        );

    \I__3259\ : CascadeMux
    port map (
            O => \N__14178\,
            I => \N__14175\
        );

    \I__3258\ : InMux
    port map (
            O => \N__14175\,
            I => \N__14169\
        );

    \I__3257\ : InMux
    port map (
            O => \N__14174\,
            I => \N__14162\
        );

    \I__3256\ : InMux
    port map (
            O => \N__14173\,
            I => \N__14162\
        );

    \I__3255\ : InMux
    port map (
            O => \N__14172\,
            I => \N__14162\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__14169\,
            I => \fifo_inst.wRamRdAddr_0\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__14162\,
            I => \fifo_inst.wRamRdAddr_0\
        );

    \I__3252\ : CascadeMux
    port map (
            O => \N__14157\,
            I => \N__14153\
        );

    \I__3251\ : CascadeMux
    port map (
            O => \N__14156\,
            I => \N__14150\
        );

    \I__3250\ : InMux
    port map (
            O => \N__14153\,
            I => \N__14146\
        );

    \I__3249\ : InMux
    port map (
            O => \N__14150\,
            I => \N__14141\
        );

    \I__3248\ : InMux
    port map (
            O => \N__14149\,
            I => \N__14141\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__14146\,
            I => \fifo_inst.wRamRdAddr_1\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__14141\,
            I => \fifo_inst.wRamRdAddr_1\
        );

    \I__3245\ : InMux
    port map (
            O => \N__14136\,
            I => \N__14133\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__14133\,
            I => \fifo_inst.ftdi_output_inst.oPacketRead_1_sqmuxa_1\
        );

    \I__3243\ : CascadeMux
    port map (
            O => \N__14130\,
            I => \N__14127\
        );

    \I__3242\ : InMux
    port map (
            O => \N__14127\,
            I => \N__14123\
        );

    \I__3241\ : InMux
    port map (
            O => \N__14126\,
            I => \N__14120\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__14123\,
            I => \fifo_inst.wRamRdAddr_2\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__14120\,
            I => \fifo_inst.wRamRdAddr_2\
        );

    \I__3238\ : InMux
    port map (
            O => \N__14115\,
            I => \N__14110\
        );

    \I__3237\ : InMux
    port map (
            O => \N__14114\,
            I => \N__14105\
        );

    \I__3236\ : InMux
    port map (
            O => \N__14113\,
            I => \N__14105\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__14110\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_3\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__14105\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_3\
        );

    \I__3233\ : CascadeMux
    port map (
            O => \N__14100\,
            I => \N__14097\
        );

    \I__3232\ : InMux
    port map (
            O => \N__14097\,
            I => \N__14094\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__14094\,
            I => \N__14091\
        );

    \I__3230\ : Odrv4
    port map (
            O => \N__14091\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_6\
        );

    \I__3229\ : InMux
    port map (
            O => \N__14088\,
            I => \N__14083\
        );

    \I__3228\ : InMux
    port map (
            O => \N__14087\,
            I => \N__14080\
        );

    \I__3227\ : InMux
    port map (
            O => \N__14086\,
            I => \N__14077\
        );

    \I__3226\ : LocalMux
    port map (
            O => \N__14083\,
            I => \N__14074\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__14080\,
            I => \N__14071\
        );

    \I__3224\ : LocalMux
    port map (
            O => \N__14077\,
            I => \N__14068\
        );

    \I__3223\ : Span4Mux_v
    port map (
            O => \N__14074\,
            I => \N__14063\
        );

    \I__3222\ : Span4Mux_h
    port map (
            O => \N__14071\,
            I => \N__14060\
        );

    \I__3221\ : Span4Mux_h
    port map (
            O => \N__14068\,
            I => \N__14057\
        );

    \I__3220\ : InMux
    port map (
            O => \N__14067\,
            I => \N__14054\
        );

    \I__3219\ : InMux
    port map (
            O => \N__14066\,
            I => \N__14051\
        );

    \I__3218\ : Odrv4
    port map (
            O => \N__14063\,
            I => \DUT.wRxByte_7\
        );

    \I__3217\ : Odrv4
    port map (
            O => \N__14060\,
            I => \DUT.wRxByte_7\
        );

    \I__3216\ : Odrv4
    port map (
            O => \N__14057\,
            I => \DUT.wRxByte_7\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__14054\,
            I => \DUT.wRxByte_7\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__14051\,
            I => \DUT.wRxByte_7\
        );

    \I__3213\ : InMux
    port map (
            O => \N__14040\,
            I => \N__14037\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__14037\,
            I => \N__14034\
        );

    \I__3211\ : Span4Mux_h
    port map (
            O => \N__14034\,
            I => \N__14031\
        );

    \I__3210\ : Odrv4
    port map (
            O => \N__14031\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_7\
        );

    \I__3209\ : CEMux
    port map (
            O => \N__14028\,
            I => \N__14025\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__14025\,
            I => \DUT.fifo_rx_inst.rFifoData_awe1\
        );

    \I__3207\ : InMux
    port map (
            O => \N__14022\,
            I => \N__14019\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__14019\,
            I => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0\
        );

    \I__3205\ : CascadeMux
    port map (
            O => \N__14016\,
            I => \N__14012\
        );

    \I__3204\ : CascadeMux
    port map (
            O => \N__14015\,
            I => \N__14008\
        );

    \I__3203\ : InMux
    port map (
            O => \N__14012\,
            I => \N__14002\
        );

    \I__3202\ : InMux
    port map (
            O => \N__14011\,
            I => \N__13991\
        );

    \I__3201\ : InMux
    port map (
            O => \N__14008\,
            I => \N__13991\
        );

    \I__3200\ : InMux
    port map (
            O => \N__14007\,
            I => \N__13991\
        );

    \I__3199\ : InMux
    port map (
            O => \N__14006\,
            I => \N__13991\
        );

    \I__3198\ : InMux
    port map (
            O => \N__14005\,
            I => \N__13991\
        );

    \I__3197\ : LocalMux
    port map (
            O => \N__14002\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_0\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__13991\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_0\
        );

    \I__3195\ : CascadeMux
    port map (
            O => \N__13986\,
            I => \N__13983\
        );

    \I__3194\ : InMux
    port map (
            O => \N__13983\,
            I => \N__13980\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__13980\,
            I => \DUT.fifo_rx_inst.rFifoCount_RNIPTFQ1Z0Z_1\
        );

    \I__3192\ : CascadeMux
    port map (
            O => \N__13977\,
            I => \N__13972\
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__13976\,
            I => \N__13969\
        );

    \I__3190\ : InMux
    port map (
            O => \N__13975\,
            I => \N__13965\
        );

    \I__3189\ : InMux
    port map (
            O => \N__13972\,
            I => \N__13958\
        );

    \I__3188\ : InMux
    port map (
            O => \N__13969\,
            I => \N__13958\
        );

    \I__3187\ : InMux
    port map (
            O => \N__13968\,
            I => \N__13958\
        );

    \I__3186\ : LocalMux
    port map (
            O => \N__13965\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_1\
        );

    \I__3185\ : LocalMux
    port map (
            O => \N__13958\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_1\
        );

    \I__3184\ : InMux
    port map (
            O => \N__13953\,
            I => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0\
        );

    \I__3183\ : InMux
    port map (
            O => \N__13950\,
            I => \N__13944\
        );

    \I__3182\ : InMux
    port map (
            O => \N__13949\,
            I => \N__13937\
        );

    \I__3181\ : InMux
    port map (
            O => \N__13948\,
            I => \N__13937\
        );

    \I__3180\ : InMux
    port map (
            O => \N__13947\,
            I => \N__13937\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__13944\,
            I => \DUT.fifo_rx_inst.N_4_0\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__13937\,
            I => \DUT.fifo_rx_inst.N_4_0\
        );

    \I__3177\ : CascadeMux
    port map (
            O => \N__13932\,
            I => \N__13929\
        );

    \I__3176\ : InMux
    port map (
            O => \N__13929\,
            I => \N__13921\
        );

    \I__3175\ : InMux
    port map (
            O => \N__13928\,
            I => \N__13910\
        );

    \I__3174\ : InMux
    port map (
            O => \N__13927\,
            I => \N__13910\
        );

    \I__3173\ : InMux
    port map (
            O => \N__13926\,
            I => \N__13910\
        );

    \I__3172\ : InMux
    port map (
            O => \N__13925\,
            I => \N__13910\
        );

    \I__3171\ : InMux
    port map (
            O => \N__13924\,
            I => \N__13910\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__13921\,
            I => \rRxReadZ0\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__13910\,
            I => \rRxReadZ0\
        );

    \I__3168\ : InMux
    port map (
            O => \N__13905\,
            I => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1\
        );

    \I__3167\ : InMux
    port map (
            O => \N__13902\,
            I => \N__13898\
        );

    \I__3166\ : InMux
    port map (
            O => \N__13901\,
            I => \N__13891\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__13898\,
            I => \N__13888\
        );

    \I__3164\ : InMux
    port map (
            O => \N__13897\,
            I => \N__13879\
        );

    \I__3163\ : InMux
    port map (
            O => \N__13896\,
            I => \N__13879\
        );

    \I__3162\ : InMux
    port map (
            O => \N__13895\,
            I => \N__13879\
        );

    \I__3161\ : InMux
    port map (
            O => \N__13894\,
            I => \N__13879\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__13891\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\
        );

    \I__3159\ : Odrv12
    port map (
            O => \N__13888\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__13879\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\
        );

    \I__3157\ : IoInMux
    port map (
            O => \N__13872\,
            I => \N__13869\
        );

    \I__3156\ : LocalMux
    port map (
            O => \N__13869\,
            I => \N__13866\
        );

    \I__3155\ : Span4Mux_s2_v
    port map (
            O => \N__13866\,
            I => \N__13863\
        );

    \I__3154\ : Odrv4
    port map (
            O => \N__13863\,
            I => \N_1261_i\
        );

    \I__3153\ : InMux
    port map (
            O => \N__13860\,
            I => \N__13857\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__13857\,
            I => \N__13854\
        );

    \I__3151\ : Odrv4
    port map (
            O => \N__13854\,
            I => \oTx_n_rep4_ess\
        );

    \I__3150\ : InMux
    port map (
            O => \N__13851\,
            I => \N__13848\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__13848\,
            I => \N__13845\
        );

    \I__3148\ : Span4Mux_s1_v
    port map (
            O => \N__13845\,
            I => \N__13842\
        );

    \I__3147\ : Span4Mux_v
    port map (
            O => \N__13842\,
            I => \N__13839\
        );

    \I__3146\ : Odrv4
    port map (
            O => \N__13839\,
            I => \oTx_n_rep1_ess\
        );

    \I__3145\ : InMux
    port map (
            O => \N__13836\,
            I => \N__13833\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__13833\,
            I => \N__13830\
        );

    \I__3143\ : Span4Mux_h
    port map (
            O => \N__13830\,
            I => \N__13827\
        );

    \I__3142\ : Span4Mux_v
    port map (
            O => \N__13827\,
            I => \N__13824\
        );

    \I__3141\ : Odrv4
    port map (
            O => \N__13824\,
            I => \oTx_n_rep0_ess\
        );

    \I__3140\ : CascadeMux
    port map (
            O => \N__13821\,
            I => \N__13818\
        );

    \I__3139\ : InMux
    port map (
            O => \N__13818\,
            I => \N__13802\
        );

    \I__3138\ : InMux
    port map (
            O => \N__13817\,
            I => \N__13802\
        );

    \I__3137\ : InMux
    port map (
            O => \N__13816\,
            I => \N__13795\
        );

    \I__3136\ : InMux
    port map (
            O => \N__13815\,
            I => \N__13795\
        );

    \I__3135\ : InMux
    port map (
            O => \N__13814\,
            I => \N__13795\
        );

    \I__3134\ : InMux
    port map (
            O => \N__13813\,
            I => \N__13792\
        );

    \I__3133\ : InMux
    port map (
            O => \N__13812\,
            I => \N__13785\
        );

    \I__3132\ : InMux
    port map (
            O => \N__13811\,
            I => \N__13785\
        );

    \I__3131\ : InMux
    port map (
            O => \N__13810\,
            I => \N__13785\
        );

    \I__3130\ : InMux
    port map (
            O => \N__13809\,
            I => \N__13778\
        );

    \I__3129\ : InMux
    port map (
            O => \N__13808\,
            I => \N__13778\
        );

    \I__3128\ : InMux
    port map (
            O => \N__13807\,
            I => \N__13778\
        );

    \I__3127\ : LocalMux
    port map (
            O => \N__13802\,
            I => \N__13773\
        );

    \I__3126\ : LocalMux
    port map (
            O => \N__13795\,
            I => \N__13773\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__13792\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__13785\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__13778\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__3122\ : Odrv4
    port map (
            O => \N__13773\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__3121\ : InMux
    port map (
            O => \N__13764\,
            I => \N__13761\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__13761\,
            I => \N__13758\
        );

    \I__3119\ : Span4Mux_v
    port map (
            O => \N__13758\,
            I => \N__13755\
        );

    \I__3118\ : Odrv4
    port map (
            O => \N__13755\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_2\
        );

    \I__3117\ : InMux
    port map (
            O => \N__13752\,
            I => \N__13749\
        );

    \I__3116\ : LocalMux
    port map (
            O => \N__13749\,
            I => \N__13746\
        );

    \I__3115\ : Odrv4
    port map (
            O => \N__13746\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_2\
        );

    \I__3114\ : CascadeMux
    port map (
            O => \N__13743\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2_cascade_\
        );

    \I__3113\ : CascadeMux
    port map (
            O => \N__13740\,
            I => \N__13726\
        );

    \I__3112\ : CascadeMux
    port map (
            O => \N__13739\,
            I => \N__13723\
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__13738\,
            I => \N__13717\
        );

    \I__3110\ : CascadeMux
    port map (
            O => \N__13737\,
            I => \N__13713\
        );

    \I__3109\ : InMux
    port map (
            O => \N__13736\,
            I => \N__13710\
        );

    \I__3108\ : CascadeMux
    port map (
            O => \N__13735\,
            I => \N__13705\
        );

    \I__3107\ : CascadeMux
    port map (
            O => \N__13734\,
            I => \N__13701\
        );

    \I__3106\ : InMux
    port map (
            O => \N__13733\,
            I => \N__13697\
        );

    \I__3105\ : InMux
    port map (
            O => \N__13732\,
            I => \N__13684\
        );

    \I__3104\ : InMux
    port map (
            O => \N__13731\,
            I => \N__13684\
        );

    \I__3103\ : InMux
    port map (
            O => \N__13730\,
            I => \N__13684\
        );

    \I__3102\ : InMux
    port map (
            O => \N__13729\,
            I => \N__13684\
        );

    \I__3101\ : InMux
    port map (
            O => \N__13726\,
            I => \N__13684\
        );

    \I__3100\ : InMux
    port map (
            O => \N__13723\,
            I => \N__13684\
        );

    \I__3099\ : InMux
    port map (
            O => \N__13722\,
            I => \N__13671\
        );

    \I__3098\ : InMux
    port map (
            O => \N__13721\,
            I => \N__13671\
        );

    \I__3097\ : InMux
    port map (
            O => \N__13720\,
            I => \N__13671\
        );

    \I__3096\ : InMux
    port map (
            O => \N__13717\,
            I => \N__13671\
        );

    \I__3095\ : InMux
    port map (
            O => \N__13716\,
            I => \N__13671\
        );

    \I__3094\ : InMux
    port map (
            O => \N__13713\,
            I => \N__13671\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__13710\,
            I => \N__13668\
        );

    \I__3092\ : InMux
    port map (
            O => \N__13709\,
            I => \N__13661\
        );

    \I__3091\ : InMux
    port map (
            O => \N__13708\,
            I => \N__13661\
        );

    \I__3090\ : InMux
    port map (
            O => \N__13705\,
            I => \N__13661\
        );

    \I__3089\ : InMux
    port map (
            O => \N__13704\,
            I => \N__13654\
        );

    \I__3088\ : InMux
    port map (
            O => \N__13701\,
            I => \N__13654\
        );

    \I__3087\ : InMux
    port map (
            O => \N__13700\,
            I => \N__13654\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__13697\,
            I => \N__13647\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__13684\,
            I => \N__13647\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__13671\,
            I => \N__13647\
        );

    \I__3083\ : Odrv4
    port map (
            O => \N__13668\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__13661\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__13654\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__3080\ : Odrv4
    port map (
            O => \N__13647\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__3079\ : InMux
    port map (
            O => \N__13638\,
            I => \N__13635\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__13635\,
            I => \DUT.fifo_rx_inst.rFifoDatarx_2\
        );

    \I__3077\ : InMux
    port map (
            O => \N__13632\,
            I => \N__13627\
        );

    \I__3076\ : InMux
    port map (
            O => \N__13631\,
            I => \N__13624\
        );

    \I__3075\ : InMux
    port map (
            O => \N__13630\,
            I => \N__13621\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__13627\,
            I => \N__13616\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__13624\,
            I => \N__13616\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__13621\,
            I => \N__13613\
        );

    \I__3071\ : Span4Mux_v
    port map (
            O => \N__13616\,
            I => \N__13609\
        );

    \I__3070\ : Span4Mux_h
    port map (
            O => \N__13613\,
            I => \N__13606\
        );

    \I__3069\ : InMux
    port map (
            O => \N__13612\,
            I => \N__13603\
        );

    \I__3068\ : Odrv4
    port map (
            O => \N__13609\,
            I => \DUT.wRxByte_0\
        );

    \I__3067\ : Odrv4
    port map (
            O => \N__13606\,
            I => \DUT.wRxByte_0\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__13603\,
            I => \DUT.wRxByte_0\
        );

    \I__3065\ : InMux
    port map (
            O => \N__13596\,
            I => \N__13593\
        );

    \I__3064\ : LocalMux
    port map (
            O => \N__13593\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_0\
        );

    \I__3063\ : InMux
    port map (
            O => \N__13590\,
            I => \N__13585\
        );

    \I__3062\ : InMux
    port map (
            O => \N__13589\,
            I => \N__13582\
        );

    \I__3061\ : InMux
    port map (
            O => \N__13588\,
            I => \N__13579\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__13585\,
            I => \N__13574\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__13582\,
            I => \N__13574\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__13579\,
            I => \N__13571\
        );

    \I__3057\ : Span4Mux_v
    port map (
            O => \N__13574\,
            I => \N__13566\
        );

    \I__3056\ : Span4Mux_h
    port map (
            O => \N__13571\,
            I => \N__13563\
        );

    \I__3055\ : InMux
    port map (
            O => \N__13570\,
            I => \N__13560\
        );

    \I__3054\ : InMux
    port map (
            O => \N__13569\,
            I => \N__13557\
        );

    \I__3053\ : Odrv4
    port map (
            O => \N__13566\,
            I => \DUT.wRxByte_1\
        );

    \I__3052\ : Odrv4
    port map (
            O => \N__13563\,
            I => \DUT.wRxByte_1\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__13560\,
            I => \DUT.wRxByte_1\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__13557\,
            I => \DUT.wRxByte_1\
        );

    \I__3049\ : InMux
    port map (
            O => \N__13548\,
            I => \N__13545\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__13545\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_1\
        );

    \I__3047\ : InMux
    port map (
            O => \N__13542\,
            I => \N__13539\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__13539\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_2\
        );

    \I__3045\ : InMux
    port map (
            O => \N__13536\,
            I => \N__13531\
        );

    \I__3044\ : InMux
    port map (
            O => \N__13535\,
            I => \N__13528\
        );

    \I__3043\ : InMux
    port map (
            O => \N__13534\,
            I => \N__13525\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__13531\,
            I => \N__13522\
        );

    \I__3041\ : LocalMux
    port map (
            O => \N__13528\,
            I => \N__13517\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__13525\,
            I => \N__13517\
        );

    \I__3039\ : Span4Mux_h
    port map (
            O => \N__13522\,
            I => \N__13512\
        );

    \I__3038\ : Span4Mux_v
    port map (
            O => \N__13517\,
            I => \N__13509\
        );

    \I__3037\ : InMux
    port map (
            O => \N__13516\,
            I => \N__13506\
        );

    \I__3036\ : InMux
    port map (
            O => \N__13515\,
            I => \N__13503\
        );

    \I__3035\ : Odrv4
    port map (
            O => \N__13512\,
            I => \DUT.wRxByte_3\
        );

    \I__3034\ : Odrv4
    port map (
            O => \N__13509\,
            I => \DUT.wRxByte_3\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__13506\,
            I => \DUT.wRxByte_3\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__13503\,
            I => \DUT.wRxByte_3\
        );

    \I__3031\ : InMux
    port map (
            O => \N__13494\,
            I => \N__13491\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__13491\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_3\
        );

    \I__3029\ : InMux
    port map (
            O => \N__13488\,
            I => \N__13484\
        );

    \I__3028\ : InMux
    port map (
            O => \N__13487\,
            I => \N__13481\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__13484\,
            I => \N__13475\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__13481\,
            I => \N__13475\
        );

    \I__3025\ : InMux
    port map (
            O => \N__13480\,
            I => \N__13472\
        );

    \I__3024\ : Span4Mux_v
    port map (
            O => \N__13475\,
            I => \N__13469\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__13472\,
            I => \N__13464\
        );

    \I__3022\ : Sp12to4
    port map (
            O => \N__13469\,
            I => \N__13461\
        );

    \I__3021\ : InMux
    port map (
            O => \N__13468\,
            I => \N__13458\
        );

    \I__3020\ : InMux
    port map (
            O => \N__13467\,
            I => \N__13455\
        );

    \I__3019\ : Odrv4
    port map (
            O => \N__13464\,
            I => \DUT.wRxByte_4\
        );

    \I__3018\ : Odrv12
    port map (
            O => \N__13461\,
            I => \DUT.wRxByte_4\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__13458\,
            I => \DUT.wRxByte_4\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__13455\,
            I => \DUT.wRxByte_4\
        );

    \I__3015\ : InMux
    port map (
            O => \N__13446\,
            I => \N__13443\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__13443\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_4\
        );

    \I__3013\ : InMux
    port map (
            O => \N__13440\,
            I => \N__13437\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__13437\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_5\
        );

    \I__3011\ : InMux
    port map (
            O => \N__13434\,
            I => \N__13430\
        );

    \I__3010\ : InMux
    port map (
            O => \N__13433\,
            I => \N__13427\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__13430\,
            I => \N__13423\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__13427\,
            I => \N__13420\
        );

    \I__3007\ : InMux
    port map (
            O => \N__13426\,
            I => \N__13417\
        );

    \I__3006\ : Span4Mux_v
    port map (
            O => \N__13423\,
            I => \N__13412\
        );

    \I__3005\ : Span4Mux_h
    port map (
            O => \N__13420\,
            I => \N__13409\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__13417\,
            I => \N__13406\
        );

    \I__3003\ : InMux
    port map (
            O => \N__13416\,
            I => \N__13403\
        );

    \I__3002\ : InMux
    port map (
            O => \N__13415\,
            I => \N__13400\
        );

    \I__3001\ : Odrv4
    port map (
            O => \N__13412\,
            I => \DUT.wRxByte_6\
        );

    \I__3000\ : Odrv4
    port map (
            O => \N__13409\,
            I => \DUT.wRxByte_6\
        );

    \I__2999\ : Odrv4
    port map (
            O => \N__13406\,
            I => \DUT.wRxByte_6\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__13403\,
            I => \DUT.wRxByte_6\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__13400\,
            I => \DUT.wRxByte_6\
        );

    \I__2996\ : InMux
    port map (
            O => \N__13389\,
            I => \N__13386\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__13386\,
            I => \DUT.fifo_rx_inst.rFifoDatarx_3\
        );

    \I__2994\ : CascadeMux
    port map (
            O => \N__13383\,
            I => \N__13380\
        );

    \I__2993\ : InMux
    port map (
            O => \N__13380\,
            I => \N__13377\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__13377\,
            I => \N__13374\
        );

    \I__2991\ : Odrv4
    port map (
            O => \N__13374\,
            I => \wRxFifoData_3\
        );

    \I__2990\ : InMux
    port map (
            O => \N__13371\,
            I => \N__13368\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__13368\,
            I => \N__13362\
        );

    \I__2988\ : InMux
    port map (
            O => \N__13367\,
            I => \N__13359\
        );

    \I__2987\ : InMux
    port map (
            O => \N__13366\,
            I => \N__13356\
        );

    \I__2986\ : InMux
    port map (
            O => \N__13365\,
            I => \N__13353\
        );

    \I__2985\ : Span4Mux_h
    port map (
            O => \N__13362\,
            I => \N__13344\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__13359\,
            I => \N__13344\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__13356\,
            I => \N__13344\
        );

    \I__2982\ : LocalMux
    port map (
            O => \N__13353\,
            I => \N__13344\
        );

    \I__2981\ : Span4Mux_v
    port map (
            O => \N__13344\,
            I => \N__13341\
        );

    \I__2980\ : Odrv4
    port map (
            O => \N__13341\,
            I => \rTxByteZ0Z_3\
        );

    \I__2979\ : InMux
    port map (
            O => \N__13338\,
            I => \N__13314\
        );

    \I__2978\ : InMux
    port map (
            O => \N__13337\,
            I => \N__13314\
        );

    \I__2977\ : InMux
    port map (
            O => \N__13336\,
            I => \N__13314\
        );

    \I__2976\ : InMux
    port map (
            O => \N__13335\,
            I => \N__13314\
        );

    \I__2975\ : InMux
    port map (
            O => \N__13334\,
            I => \N__13314\
        );

    \I__2974\ : InMux
    port map (
            O => \N__13333\,
            I => \N__13314\
        );

    \I__2973\ : InMux
    port map (
            O => \N__13332\,
            I => \N__13314\
        );

    \I__2972\ : InMux
    port map (
            O => \N__13331\,
            I => \N__13314\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__13314\,
            I => \DUT.fifo_rx_inst.rFifoDataror_0\
        );

    \I__2970\ : CascadeMux
    port map (
            O => \N__13311\,
            I => \N__13308\
        );

    \I__2969\ : InMux
    port map (
            O => \N__13308\,
            I => \N__13305\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__13305\,
            I => \N__13302\
        );

    \I__2967\ : Odrv12
    port map (
            O => \N__13302\,
            I => \wRxFifoData_4\
        );

    \I__2966\ : InMux
    port map (
            O => \N__13299\,
            I => \N__13296\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__13296\,
            I => \DUT.fifo_rx_inst.rFifoDatarx_4\
        );

    \I__2964\ : InMux
    port map (
            O => \N__13293\,
            I => \N__13289\
        );

    \I__2963\ : InMux
    port map (
            O => \N__13292\,
            I => \N__13286\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__13289\,
            I => \N__13282\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__13286\,
            I => \N__13279\
        );

    \I__2960\ : InMux
    port map (
            O => \N__13285\,
            I => \N__13276\
        );

    \I__2959\ : Span4Mux_v
    port map (
            O => \N__13282\,
            I => \N__13268\
        );

    \I__2958\ : Span4Mux_h
    port map (
            O => \N__13279\,
            I => \N__13268\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__13276\,
            I => \N__13268\
        );

    \I__2956\ : InMux
    port map (
            O => \N__13275\,
            I => \N__13265\
        );

    \I__2955\ : Sp12to4
    port map (
            O => \N__13268\,
            I => \N__13260\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__13265\,
            I => \N__13260\
        );

    \I__2953\ : Odrv12
    port map (
            O => \N__13260\,
            I => \rTxByteZ0Z_4\
        );

    \I__2952\ : CEMux
    port map (
            O => \N__13257\,
            I => \N__13254\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__13254\,
            I => \N__13251\
        );

    \I__2950\ : Span4Mux_v
    port map (
            O => \N__13251\,
            I => \N__13248\
        );

    \I__2949\ : Odrv4
    port map (
            O => \N__13248\,
            I => \rTxByte_1_sqmuxa_i_0\
        );

    \I__2948\ : InMux
    port map (
            O => \N__13245\,
            I => \N__13242\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__13242\,
            I => \N__13239\
        );

    \I__2946\ : Odrv4
    port map (
            O => \N__13239\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_0\
        );

    \I__2945\ : InMux
    port map (
            O => \N__13236\,
            I => \N__13233\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__13233\,
            I => \N__13230\
        );

    \I__2943\ : Span4Mux_h
    port map (
            O => \N__13230\,
            I => \N__13227\
        );

    \I__2942\ : Odrv4
    port map (
            O => \N__13227\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_0\
        );

    \I__2941\ : CascadeMux
    port map (
            O => \N__13224\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_\
        );

    \I__2940\ : InMux
    port map (
            O => \N__13221\,
            I => \N__13218\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__13218\,
            I => \DUT.fifo_rx_inst.rFifoDatarx_0\
        );

    \I__2938\ : InMux
    port map (
            O => \N__13215\,
            I => \N__13212\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__13212\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_0\
        );

    \I__2936\ : InMux
    port map (
            O => \N__13209\,
            I => \N__13206\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__13206\,
            I => \N__13203\
        );

    \I__2934\ : Span4Mux_h
    port map (
            O => \N__13203\,
            I => \N__13200\
        );

    \I__2933\ : Odrv4
    port map (
            O => \N__13200\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_1\
        );

    \I__2932\ : CascadeMux
    port map (
            O => \N__13197\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1_cascade_\
        );

    \I__2931\ : InMux
    port map (
            O => \N__13194\,
            I => \N__13191\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__13191\,
            I => \N__13188\
        );

    \I__2929\ : Odrv4
    port map (
            O => \N__13188\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_1\
        );

    \I__2928\ : InMux
    port map (
            O => \N__13185\,
            I => \N__13182\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__13182\,
            I => \DUT.fifo_rx_inst.rFifoDatarx_1\
        );

    \I__2926\ : CascadeMux
    port map (
            O => \N__13179\,
            I => \N__13176\
        );

    \I__2925\ : InMux
    port map (
            O => \N__13176\,
            I => \N__13173\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__13173\,
            I => \N__13170\
        );

    \I__2923\ : Odrv4
    port map (
            O => \N__13170\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_1\
        );

    \I__2922\ : InMux
    port map (
            O => \N__13167\,
            I => \N__13164\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__13164\,
            I => \N__13161\
        );

    \I__2920\ : Span4Mux_h
    port map (
            O => \N__13161\,
            I => \N__13158\
        );

    \I__2919\ : Odrv4
    port map (
            O => \N__13158\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_5\
        );

    \I__2918\ : InMux
    port map (
            O => \N__13155\,
            I => \N__13152\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__13152\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_6\
        );

    \I__2916\ : InMux
    port map (
            O => \N__13149\,
            I => \N__13146\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__13146\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_7\
        );

    \I__2914\ : CEMux
    port map (
            O => \N__13143\,
            I => \N__13140\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__13140\,
            I => \N__13137\
        );

    \I__2912\ : Span4Mux_v
    port map (
            O => \N__13137\,
            I => \N__13134\
        );

    \I__2911\ : Odrv4
    port map (
            O => \N__13134\,
            I => \DUT.fifo_rx_inst.rFifoData_awe2\
        );

    \I__2910\ : InMux
    port map (
            O => \N__13131\,
            I => \N__13128\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__13128\,
            I => \DUT.fifo_rx_inst.rFifoDatarx_6\
        );

    \I__2908\ : InMux
    port map (
            O => \N__13125\,
            I => \N__13122\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__13122\,
            I => \N__13119\
        );

    \I__2906\ : Odrv12
    port map (
            O => \N__13119\,
            I => \wRxFifoData_6\
        );

    \I__2905\ : InMux
    port map (
            O => \N__13116\,
            I => \N__13112\
        );

    \I__2904\ : InMux
    port map (
            O => \N__13115\,
            I => \N__13109\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__13112\,
            I => \N__13105\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__13109\,
            I => \N__13101\
        );

    \I__2901\ : InMux
    port map (
            O => \N__13108\,
            I => \N__13098\
        );

    \I__2900\ : Span4Mux_h
    port map (
            O => \N__13105\,
            I => \N__13095\
        );

    \I__2899\ : InMux
    port map (
            O => \N__13104\,
            I => \N__13092\
        );

    \I__2898\ : Span4Mux_v
    port map (
            O => \N__13101\,
            I => \N__13087\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__13098\,
            I => \N__13087\
        );

    \I__2896\ : Sp12to4
    port map (
            O => \N__13095\,
            I => \N__13082\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__13092\,
            I => \N__13082\
        );

    \I__2894\ : Odrv4
    port map (
            O => \N__13087\,
            I => \rTxByteZ0Z_6\
        );

    \I__2893\ : Odrv12
    port map (
            O => \N__13082\,
            I => \rTxByteZ0Z_6\
        );

    \I__2892\ : CascadeMux
    port map (
            O => \N__13077\,
            I => \N__13074\
        );

    \I__2891\ : InMux
    port map (
            O => \N__13074\,
            I => \N__13071\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__13071\,
            I => \N__13068\
        );

    \I__2889\ : Odrv4
    port map (
            O => \N__13068\,
            I => \wRxFifoData_5\
        );

    \I__2888\ : InMux
    port map (
            O => \N__13065\,
            I => \N__13062\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__13062\,
            I => \DUT.fifo_rx_inst.rFifoDatarx_5\
        );

    \I__2886\ : InMux
    port map (
            O => \N__13059\,
            I => \N__13055\
        );

    \I__2885\ : InMux
    port map (
            O => \N__13058\,
            I => \N__13052\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__13055\,
            I => \N__13047\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__13052\,
            I => \N__13044\
        );

    \I__2882\ : InMux
    port map (
            O => \N__13051\,
            I => \N__13041\
        );

    \I__2881\ : InMux
    port map (
            O => \N__13050\,
            I => \N__13038\
        );

    \I__2880\ : Span4Mux_v
    port map (
            O => \N__13047\,
            I => \N__13031\
        );

    \I__2879\ : Span4Mux_h
    port map (
            O => \N__13044\,
            I => \N__13031\
        );

    \I__2878\ : LocalMux
    port map (
            O => \N__13041\,
            I => \N__13031\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__13038\,
            I => \N__13028\
        );

    \I__2876\ : Odrv4
    port map (
            O => \N__13031\,
            I => \rTxByteZ0Z_5\
        );

    \I__2875\ : Odrv12
    port map (
            O => \N__13028\,
            I => \rTxByteZ0Z_5\
        );

    \I__2874\ : CascadeMux
    port map (
            O => \N__13023\,
            I => \N__13020\
        );

    \I__2873\ : InMux
    port map (
            O => \N__13020\,
            I => \N__13017\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__13017\,
            I => \N__13014\
        );

    \I__2871\ : Odrv4
    port map (
            O => \N__13014\,
            I => \wRxFifoData_0\
        );

    \I__2870\ : InMux
    port map (
            O => \N__13011\,
            I => \N__13008\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__13008\,
            I => \N__13004\
        );

    \I__2868\ : InMux
    port map (
            O => \N__13007\,
            I => \N__13001\
        );

    \I__2867\ : Span4Mux_h
    port map (
            O => \N__13004\,
            I => \N__12996\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__13001\,
            I => \N__12993\
        );

    \I__2865\ : InMux
    port map (
            O => \N__13000\,
            I => \N__12990\
        );

    \I__2864\ : InMux
    port map (
            O => \N__12999\,
            I => \N__12987\
        );

    \I__2863\ : Span4Mux_v
    port map (
            O => \N__12996\,
            I => \N__12984\
        );

    \I__2862\ : Span4Mux_v
    port map (
            O => \N__12993\,
            I => \N__12979\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__12990\,
            I => \N__12979\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__12987\,
            I => \N__12976\
        );

    \I__2859\ : Odrv4
    port map (
            O => \N__12984\,
            I => \rTxByteZ0Z_0\
        );

    \I__2858\ : Odrv4
    port map (
            O => \N__12979\,
            I => \rTxByteZ0Z_0\
        );

    \I__2857\ : Odrv12
    port map (
            O => \N__12976\,
            I => \rTxByteZ0Z_0\
        );

    \I__2856\ : InMux
    port map (
            O => \N__12969\,
            I => \N__12966\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__12966\,
            I => \DUT.fifo_rx_inst.rFifoDatarx_7\
        );

    \I__2854\ : InMux
    port map (
            O => \N__12963\,
            I => \N__12960\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__12960\,
            I => \N__12955\
        );

    \I__2852\ : InMux
    port map (
            O => \N__12959\,
            I => \N__12952\
        );

    \I__2851\ : InMux
    port map (
            O => \N__12958\,
            I => \N__12949\
        );

    \I__2850\ : Span4Mux_h
    port map (
            O => \N__12955\,
            I => \N__12945\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__12952\,
            I => \N__12942\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__12949\,
            I => \N__12939\
        );

    \I__2847\ : InMux
    port map (
            O => \N__12948\,
            I => \N__12936\
        );

    \I__2846\ : Span4Mux_v
    port map (
            O => \N__12945\,
            I => \N__12933\
        );

    \I__2845\ : Span4Mux_v
    port map (
            O => \N__12942\,
            I => \N__12930\
        );

    \I__2844\ : Span4Mux_h
    port map (
            O => \N__12939\,
            I => \N__12927\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__12936\,
            I => \N__12924\
        );

    \I__2842\ : Odrv4
    port map (
            O => \N__12933\,
            I => \rTxByteZ0Z_7\
        );

    \I__2841\ : Odrv4
    port map (
            O => \N__12930\,
            I => \rTxByteZ0Z_7\
        );

    \I__2840\ : Odrv4
    port map (
            O => \N__12927\,
            I => \rTxByteZ0Z_7\
        );

    \I__2839\ : Odrv12
    port map (
            O => \N__12924\,
            I => \rTxByteZ0Z_7\
        );

    \I__2838\ : CascadeMux
    port map (
            O => \N__12915\,
            I => \N__12912\
        );

    \I__2837\ : InMux
    port map (
            O => \N__12912\,
            I => \N__12909\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__12909\,
            I => \N__12906\
        );

    \I__2835\ : Odrv4
    port map (
            O => \N__12906\,
            I => \wRxFifoData_1\
        );

    \I__2834\ : InMux
    port map (
            O => \N__12903\,
            I => \N__12899\
        );

    \I__2833\ : InMux
    port map (
            O => \N__12902\,
            I => \N__12896\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__12899\,
            I => \N__12891\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__12896\,
            I => \N__12888\
        );

    \I__2830\ : InMux
    port map (
            O => \N__12895\,
            I => \N__12885\
        );

    \I__2829\ : InMux
    port map (
            O => \N__12894\,
            I => \N__12882\
        );

    \I__2828\ : Span4Mux_h
    port map (
            O => \N__12891\,
            I => \N__12879\
        );

    \I__2827\ : Span4Mux_h
    port map (
            O => \N__12888\,
            I => \N__12874\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__12885\,
            I => \N__12874\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__12882\,
            I => \N__12871\
        );

    \I__2824\ : Span4Mux_v
    port map (
            O => \N__12879\,
            I => \N__12868\
        );

    \I__2823\ : Span4Mux_v
    port map (
            O => \N__12874\,
            I => \N__12865\
        );

    \I__2822\ : Span4Mux_h
    port map (
            O => \N__12871\,
            I => \N__12862\
        );

    \I__2821\ : Odrv4
    port map (
            O => \N__12868\,
            I => \rTxByteZ0Z_1\
        );

    \I__2820\ : Odrv4
    port map (
            O => \N__12865\,
            I => \rTxByteZ0Z_1\
        );

    \I__2819\ : Odrv4
    port map (
            O => \N__12862\,
            I => \rTxByteZ0Z_1\
        );

    \I__2818\ : CascadeMux
    port map (
            O => \N__12855\,
            I => \N__12852\
        );

    \I__2817\ : InMux
    port map (
            O => \N__12852\,
            I => \N__12849\
        );

    \I__2816\ : LocalMux
    port map (
            O => \N__12849\,
            I => \N__12846\
        );

    \I__2815\ : Odrv4
    port map (
            O => \N__12846\,
            I => \wRxFifoData_2\
        );

    \I__2814\ : InMux
    port map (
            O => \N__12843\,
            I => \N__12840\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__12840\,
            I => \N__12834\
        );

    \I__2812\ : InMux
    port map (
            O => \N__12839\,
            I => \N__12831\
        );

    \I__2811\ : InMux
    port map (
            O => \N__12838\,
            I => \N__12828\
        );

    \I__2810\ : InMux
    port map (
            O => \N__12837\,
            I => \N__12825\
        );

    \I__2809\ : Span4Mux_h
    port map (
            O => \N__12834\,
            I => \N__12816\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__12831\,
            I => \N__12816\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__12828\,
            I => \N__12816\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__12825\,
            I => \N__12816\
        );

    \I__2805\ : Span4Mux_v
    port map (
            O => \N__12816\,
            I => \N__12813\
        );

    \I__2804\ : Odrv4
    port map (
            O => \N__12813\,
            I => \rTxByteZ0Z_2\
        );

    \I__2803\ : InMux
    port map (
            O => \N__12810\,
            I => \N__12807\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__12807\,
            I => \N__12804\
        );

    \I__2801\ : Span12Mux_h
    port map (
            O => \N__12804\,
            I => \N__12801\
        );

    \I__2800\ : Odrv12
    port map (
            O => \N__12801\,
            I => \ioFifoData_in_2\
        );

    \I__2799\ : InMux
    port map (
            O => \N__12798\,
            I => \N__12795\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__12795\,
            I => \N__12792\
        );

    \I__2797\ : Span12Mux_h
    port map (
            O => \N__12792\,
            I => \N__12789\
        );

    \I__2796\ : Odrv12
    port map (
            O => \N__12789\,
            I => \ioFifoData_in_0\
        );

    \I__2795\ : InMux
    port map (
            O => \N__12786\,
            I => \N__12783\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__12783\,
            I => \N__12780\
        );

    \I__2793\ : Sp12to4
    port map (
            O => \N__12780\,
            I => \N__12777\
        );

    \I__2792\ : Span12Mux_v
    port map (
            O => \N__12777\,
            I => \N__12774\
        );

    \I__2791\ : Odrv12
    port map (
            O => \N__12774\,
            I => \ioFifoData_in_6\
        );

    \I__2790\ : InMux
    port map (
            O => \N__12771\,
            I => \N__12768\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__12768\,
            I => \N__12765\
        );

    \I__2788\ : Span4Mux_v
    port map (
            O => \N__12765\,
            I => \N__12762\
        );

    \I__2787\ : Odrv4
    port map (
            O => \N__12762\,
            I => \ioFifoData_in_4\
        );

    \I__2786\ : InMux
    port map (
            O => \N__12759\,
            I => \N__12756\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__12756\,
            I => \N__12753\
        );

    \I__2784\ : Span4Mux_v
    port map (
            O => \N__12753\,
            I => \N__12750\
        );

    \I__2783\ : Odrv4
    port map (
            O => \N__12750\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_3\
        );

    \I__2782\ : InMux
    port map (
            O => \N__12747\,
            I => \N__12744\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__12744\,
            I => \N__12741\
        );

    \I__2780\ : Odrv4
    port map (
            O => \N__12741\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_4\
        );

    \I__2779\ : InMux
    port map (
            O => \N__12738\,
            I => \N__12735\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__12735\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_2\
        );

    \I__2777\ : InMux
    port map (
            O => \N__12732\,
            I => \N__12729\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__12729\,
            I => \N__12726\
        );

    \I__2775\ : Odrv4
    port map (
            O => \N__12726\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_3\
        );

    \I__2774\ : InMux
    port map (
            O => \N__12723\,
            I => \N__12720\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__12720\,
            I => \N__12717\
        );

    \I__2772\ : Span4Mux_h
    port map (
            O => \N__12717\,
            I => \N__12714\
        );

    \I__2771\ : Odrv4
    port map (
            O => \N__12714\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_4\
        );

    \I__2770\ : InMux
    port map (
            O => \N__12711\,
            I => \N__12708\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__12708\,
            I => \N__12705\
        );

    \I__2768\ : Span4Mux_h
    port map (
            O => \N__12705\,
            I => \N__12702\
        );

    \I__2767\ : Odrv4
    port map (
            O => \N__12702\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_5\
        );

    \I__2766\ : InMux
    port map (
            O => \N__12699\,
            I => \N__12696\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__12696\,
            I => \N__12693\
        );

    \I__2764\ : Odrv12
    port map (
            O => \N__12693\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_6\
        );

    \I__2763\ : InMux
    port map (
            O => \N__12690\,
            I => \N__12687\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__12687\,
            I => \N__12684\
        );

    \I__2761\ : Span4Mux_h
    port map (
            O => \N__12684\,
            I => \N__12681\
        );

    \I__2760\ : Odrv4
    port map (
            O => \N__12681\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_7\
        );

    \I__2759\ : CEMux
    port map (
            O => \N__12678\,
            I => \N__12675\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__12675\,
            I => \N__12672\
        );

    \I__2757\ : Span4Mux_v
    port map (
            O => \N__12672\,
            I => \N__12668\
        );

    \I__2756\ : InMux
    port map (
            O => \N__12671\,
            I => \N__12665\
        );

    \I__2755\ : Span4Mux_h
    port map (
            O => \N__12668\,
            I => \N__12660\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__12665\,
            I => \N__12660\
        );

    \I__2753\ : Span4Mux_h
    port map (
            O => \N__12660\,
            I => \N__12656\
        );

    \I__2752\ : InMux
    port map (
            O => \N__12659\,
            I => \N__12653\
        );

    \I__2751\ : Odrv4
    port map (
            O => \N__12656\,
            I => \DUT.fifo_tx_inst.rFifoData_awe3\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__12653\,
            I => \DUT.fifo_tx_inst.rFifoData_awe3\
        );

    \I__2749\ : InMux
    port map (
            O => \N__12648\,
            I => \N__12645\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__12645\,
            I => \N__12642\
        );

    \I__2747\ : Span4Mux_h
    port map (
            O => \N__12642\,
            I => \N__12639\
        );

    \I__2746\ : Span4Mux_v
    port map (
            O => \N__12639\,
            I => \N__12636\
        );

    \I__2745\ : Odrv4
    port map (
            O => \N__12636\,
            I => \ioFifoData_in_3\
        );

    \I__2744\ : InMux
    port map (
            O => \N__12633\,
            I => \N__12630\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__12630\,
            I => \N__12627\
        );

    \I__2742\ : Span4Mux_h
    port map (
            O => \N__12627\,
            I => \N__12624\
        );

    \I__2741\ : Span4Mux_v
    port map (
            O => \N__12624\,
            I => \N__12621\
        );

    \I__2740\ : Odrv4
    port map (
            O => \N__12621\,
            I => \ioFifoData_in_1\
        );

    \I__2739\ : InMux
    port map (
            O => \N__12618\,
            I => \N__12615\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__12615\,
            I => \N__12612\
        );

    \I__2737\ : Odrv12
    port map (
            O => \N__12612\,
            I => \ioFifoData_in_5\
        );

    \I__2736\ : CascadeMux
    port map (
            O => \N__12609\,
            I => \N__12605\
        );

    \I__2735\ : InMux
    port map (
            O => \N__12608\,
            I => \N__12601\
        );

    \I__2734\ : InMux
    port map (
            O => \N__12605\,
            I => \N__12596\
        );

    \I__2733\ : InMux
    port map (
            O => \N__12604\,
            I => \N__12596\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__12601\,
            I => \N__12593\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__12596\,
            I => \N__12589\
        );

    \I__2730\ : Span4Mux_v
    port map (
            O => \N__12593\,
            I => \N__12586\
        );

    \I__2729\ : InMux
    port map (
            O => \N__12592\,
            I => \N__12583\
        );

    \I__2728\ : Span4Mux_h
    port map (
            O => \N__12589\,
            I => \N__12580\
        );

    \I__2727\ : Odrv4
    port map (
            O => \N__12586\,
            I => \DUT.wRcvd\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__12583\,
            I => \DUT.wRcvd\
        );

    \I__2725\ : Odrv4
    port map (
            O => \N__12580\,
            I => \DUT.wRcvd\
        );

    \I__2724\ : InMux
    port map (
            O => \N__12573\,
            I => \N__12567\
        );

    \I__2723\ : InMux
    port map (
            O => \N__12572\,
            I => \N__12567\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__12567\,
            I => \N__12563\
        );

    \I__2721\ : CascadeMux
    port map (
            O => \N__12566\,
            I => \N__12560\
        );

    \I__2720\ : Span4Mux_h
    port map (
            O => \N__12563\,
            I => \N__12557\
        );

    \I__2719\ : InMux
    port map (
            O => \N__12560\,
            I => \N__12554\
        );

    \I__2718\ : Odrv4
    port map (
            O => \N__12557\,
            I => \DUT.fifo_rx_inst.N_46\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__12554\,
            I => \DUT.fifo_rx_inst.N_46\
        );

    \I__2716\ : InMux
    port map (
            O => \N__12549\,
            I => \N__12546\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__12546\,
            I => \N__12543\
        );

    \I__2714\ : Span4Mux_h
    port map (
            O => \N__12543\,
            I => \N__12540\
        );

    \I__2713\ : Span4Mux_h
    port map (
            O => \N__12540\,
            I => \N__12536\
        );

    \I__2712\ : InMux
    port map (
            O => \N__12539\,
            I => \N__12533\
        );

    \I__2711\ : Odrv4
    port map (
            O => \N__12536\,
            I => \N_69_mux\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__12533\,
            I => \N_69_mux\
        );

    \I__2709\ : CascadeMux
    port map (
            O => \N__12528\,
            I => \N_69_mux_cascade_\
        );

    \I__2708\ : IoInMux
    port map (
            O => \N__12525\,
            I => \N__12522\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__12522\,
            I => \N__12519\
        );

    \I__2706\ : IoSpan4Mux
    port map (
            O => \N__12519\,
            I => \N__12516\
        );

    \I__2705\ : Odrv4
    port map (
            O => \N__12516\,
            I => \N_1258_i\
        );

    \I__2704\ : IoInMux
    port map (
            O => \N__12513\,
            I => \N__12509\
        );

    \I__2703\ : IoInMux
    port map (
            O => \N__12512\,
            I => \N__12506\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__12509\,
            I => \N__12501\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__12506\,
            I => \N__12501\
        );

    \I__2700\ : Span4Mux_s1_v
    port map (
            O => \N__12501\,
            I => \N__12498\
        );

    \I__2699\ : Sp12to4
    port map (
            O => \N__12498\,
            I => \N__12495\
        );

    \I__2698\ : Span12Mux_s7_h
    port map (
            O => \N__12495\,
            I => \N__12492\
        );

    \I__2697\ : Span12Mux_v
    port map (
            O => \N__12492\,
            I => \N__12488\
        );

    \I__2696\ : IoInMux
    port map (
            O => \N__12491\,
            I => \N__12485\
        );

    \I__2695\ : Span12Mux_v
    port map (
            O => \N__12488\,
            I => \N__12482\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__12485\,
            I => \N__12479\
        );

    \I__2693\ : Odrv12
    port map (
            O => \N__12482\,
            I => \P1A4_c_i\
        );

    \I__2692\ : Odrv4
    port map (
            O => \N__12479\,
            I => \P1A4_c_i\
        );

    \I__2691\ : InMux
    port map (
            O => \N__12474\,
            I => \N__12471\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__12471\,
            I => \N__12468\
        );

    \I__2689\ : Span4Mux_v
    port map (
            O => \N__12468\,
            I => \N__12465\
        );

    \I__2688\ : Odrv4
    port map (
            O => \N__12465\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_0\
        );

    \I__2687\ : InMux
    port map (
            O => \N__12462\,
            I => \N__12459\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__12459\,
            I => \N__12456\
        );

    \I__2685\ : Span4Mux_v
    port map (
            O => \N__12456\,
            I => \N__12453\
        );

    \I__2684\ : Odrv4
    port map (
            O => \N__12453\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_1\
        );

    \I__2683\ : InMux
    port map (
            O => \N__12450\,
            I => \N__12446\
        );

    \I__2682\ : InMux
    port map (
            O => \N__12449\,
            I => \N__12443\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__12446\,
            I => \N__12440\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__12443\,
            I => \DUT.fifo_rx_inst.rFifoDataro_0\
        );

    \I__2679\ : Odrv4
    port map (
            O => \N__12440\,
            I => \DUT.fifo_rx_inst.rFifoDataro_0\
        );

    \I__2678\ : CascadeMux
    port map (
            O => \N__12435\,
            I => \N__12431\
        );

    \I__2677\ : InMux
    port map (
            O => \N__12434\,
            I => \N__12428\
        );

    \I__2676\ : InMux
    port map (
            O => \N__12431\,
            I => \N__12425\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__12428\,
            I => \N__12422\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__12425\,
            I => \DUT.fifo_rx_inst.rFifoDataro_1\
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__12422\,
            I => \DUT.fifo_rx_inst.rFifoDataro_1\
        );

    \I__2672\ : InMux
    port map (
            O => \N__12417\,
            I => \N__12413\
        );

    \I__2671\ : InMux
    port map (
            O => \N__12416\,
            I => \N__12410\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__12413\,
            I => \N__12407\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__12410\,
            I => \DUT.fifo_rx_inst.rFifoDataro_2\
        );

    \I__2668\ : Odrv4
    port map (
            O => \N__12407\,
            I => \DUT.fifo_rx_inst.rFifoDataro_2\
        );

    \I__2667\ : CascadeMux
    port map (
            O => \N__12402\,
            I => \N__12397\
        );

    \I__2666\ : CascadeMux
    port map (
            O => \N__12401\,
            I => \N__12393\
        );

    \I__2665\ : CascadeMux
    port map (
            O => \N__12400\,
            I => \N__12390\
        );

    \I__2664\ : InMux
    port map (
            O => \N__12397\,
            I => \N__12375\
        );

    \I__2663\ : InMux
    port map (
            O => \N__12396\,
            I => \N__12375\
        );

    \I__2662\ : InMux
    port map (
            O => \N__12393\,
            I => \N__12375\
        );

    \I__2661\ : InMux
    port map (
            O => \N__12390\,
            I => \N__12375\
        );

    \I__2660\ : InMux
    port map (
            O => \N__12389\,
            I => \N__12375\
        );

    \I__2659\ : InMux
    port map (
            O => \N__12388\,
            I => \N__12375\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__12375\,
            I => \N__12371\
        );

    \I__2657\ : CascadeMux
    port map (
            O => \N__12374\,
            I => \N__12366\
        );

    \I__2656\ : Span4Mux_v
    port map (
            O => \N__12371\,
            I => \N__12363\
        );

    \I__2655\ : InMux
    port map (
            O => \N__12370\,
            I => \N__12356\
        );

    \I__2654\ : InMux
    port map (
            O => \N__12369\,
            I => \N__12356\
        );

    \I__2653\ : InMux
    port map (
            O => \N__12366\,
            I => \N__12356\
        );

    \I__2652\ : Odrv4
    port map (
            O => \N__12363\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_0\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__12356\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_0\
        );

    \I__2650\ : InMux
    port map (
            O => \N__12351\,
            I => \N__12333\
        );

    \I__2649\ : InMux
    port map (
            O => \N__12350\,
            I => \N__12333\
        );

    \I__2648\ : InMux
    port map (
            O => \N__12349\,
            I => \N__12333\
        );

    \I__2647\ : InMux
    port map (
            O => \N__12348\,
            I => \N__12333\
        );

    \I__2646\ : InMux
    port map (
            O => \N__12347\,
            I => \N__12333\
        );

    \I__2645\ : InMux
    port map (
            O => \N__12346\,
            I => \N__12333\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__12333\,
            I => \N__12330\
        );

    \I__2643\ : Span4Mux_v
    port map (
            O => \N__12330\,
            I => \N__12325\
        );

    \I__2642\ : InMux
    port map (
            O => \N__12329\,
            I => \N__12320\
        );

    \I__2641\ : InMux
    port map (
            O => \N__12328\,
            I => \N__12320\
        );

    \I__2640\ : Odrv4
    port map (
            O => \N__12325\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_1\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__12320\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_1\
        );

    \I__2638\ : InMux
    port map (
            O => \N__12315\,
            I => \N__12308\
        );

    \I__2637\ : InMux
    port map (
            O => \N__12314\,
            I => \N__12305\
        );

    \I__2636\ : InMux
    port map (
            O => \N__12313\,
            I => \N__12302\
        );

    \I__2635\ : InMux
    port map (
            O => \N__12312\,
            I => \N__12296\
        );

    \I__2634\ : InMux
    port map (
            O => \N__12311\,
            I => \N__12296\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__12308\,
            I => \N__12289\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__12305\,
            I => \N__12289\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__12302\,
            I => \N__12289\
        );

    \I__2630\ : InMux
    port map (
            O => \N__12301\,
            I => \N__12286\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__12296\,
            I => \N__12283\
        );

    \I__2628\ : Odrv4
    port map (
            O => \N__12289\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_0\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__12286\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_0\
        );

    \I__2626\ : Odrv4
    port map (
            O => \N__12283\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_0\
        );

    \I__2625\ : InMux
    port map (
            O => \N__12276\,
            I => \N__12273\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__12273\,
            I => \N__12268\
        );

    \I__2623\ : InMux
    port map (
            O => \N__12272\,
            I => \N__12265\
        );

    \I__2622\ : InMux
    port map (
            O => \N__12271\,
            I => \N__12260\
        );

    \I__2621\ : Span4Mux_h
    port map (
            O => \N__12268\,
            I => \N__12255\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__12265\,
            I => \N__12255\
        );

    \I__2619\ : InMux
    port map (
            O => \N__12264\,
            I => \N__12250\
        );

    \I__2618\ : InMux
    port map (
            O => \N__12263\,
            I => \N__12250\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__12260\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_1\
        );

    \I__2616\ : Odrv4
    port map (
            O => \N__12255\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_1\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__12250\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_1\
        );

    \I__2614\ : InMux
    port map (
            O => \N__12243\,
            I => \N__12235\
        );

    \I__2613\ : InMux
    port map (
            O => \N__12242\,
            I => \N__12232\
        );

    \I__2612\ : InMux
    port map (
            O => \N__12241\,
            I => \N__12229\
        );

    \I__2611\ : InMux
    port map (
            O => \N__12240\,
            I => \N__12226\
        );

    \I__2610\ : InMux
    port map (
            O => \N__12239\,
            I => \N__12221\
        );

    \I__2609\ : InMux
    port map (
            O => \N__12238\,
            I => \N__12221\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__12235\,
            I => \N__12214\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__12232\,
            I => \N__12214\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__12229\,
            I => \N__12214\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__12226\,
            I => \DUT.fifo_tx_inst.N_104\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__12221\,
            I => \DUT.fifo_tx_inst.N_104\
        );

    \I__2603\ : Odrv12
    port map (
            O => \N__12214\,
            I => \DUT.fifo_tx_inst.N_104\
        );

    \I__2602\ : CEMux
    port map (
            O => \N__12207\,
            I => \N__12204\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__12204\,
            I => \N__12200\
        );

    \I__2600\ : InMux
    port map (
            O => \N__12203\,
            I => \N__12197\
        );

    \I__2599\ : Span4Mux_v
    port map (
            O => \N__12200\,
            I => \N__12194\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__12197\,
            I => \N__12191\
        );

    \I__2597\ : Odrv4
    port map (
            O => \N__12194\,
            I => \DUT.fifo_tx_inst.rFifoData_awe2\
        );

    \I__2596\ : Odrv12
    port map (
            O => \N__12191\,
            I => \DUT.fifo_tx_inst.rFifoData_awe2\
        );

    \I__2595\ : CascadeMux
    port map (
            O => \N__12186\,
            I => \DUT.fifo_rx_inst.rWritePtr16_cascade_\
        );

    \I__2594\ : CascadeMux
    port map (
            O => \N__12183\,
            I => \N__12180\
        );

    \I__2593\ : InMux
    port map (
            O => \N__12180\,
            I => \N__12174\
        );

    \I__2592\ : InMux
    port map (
            O => \N__12179\,
            I => \N__12174\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__12174\,
            I => \N__12171\
        );

    \I__2590\ : Span4Mux_h
    port map (
            O => \N__12171\,
            I => \N__12161\
        );

    \I__2589\ : InMux
    port map (
            O => \N__12170\,
            I => \N__12158\
        );

    \I__2588\ : InMux
    port map (
            O => \N__12169\,
            I => \N__12145\
        );

    \I__2587\ : InMux
    port map (
            O => \N__12168\,
            I => \N__12145\
        );

    \I__2586\ : InMux
    port map (
            O => \N__12167\,
            I => \N__12145\
        );

    \I__2585\ : InMux
    port map (
            O => \N__12166\,
            I => \N__12145\
        );

    \I__2584\ : InMux
    port map (
            O => \N__12165\,
            I => \N__12145\
        );

    \I__2583\ : InMux
    port map (
            O => \N__12164\,
            I => \N__12145\
        );

    \I__2582\ : Odrv4
    port map (
            O => \N__12161\,
            I => \DUT.fifo_rx_inst.rWritePtr16\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__12158\,
            I => \DUT.fifo_rx_inst.rWritePtr16\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__12145\,
            I => \DUT.fifo_rx_inst.rWritePtr16\
        );

    \I__2579\ : CascadeMux
    port map (
            O => \N__12138\,
            I => \DUT.fifo_rx_inst.rFifoDataror_1_0_cascade_\
        );

    \I__2578\ : InMux
    port map (
            O => \N__12135\,
            I => \N__12132\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__12132\,
            I => \N__12129\
        );

    \I__2576\ : Odrv4
    port map (
            O => \N__12129\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_3\
        );

    \I__2575\ : CascadeMux
    port map (
            O => \N__12126\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_\
        );

    \I__2574\ : InMux
    port map (
            O => \N__12123\,
            I => \N__12120\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__12120\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_3\
        );

    \I__2572\ : InMux
    port map (
            O => \N__12117\,
            I => \N__12114\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__12114\,
            I => \N__12111\
        );

    \I__2570\ : Odrv4
    port map (
            O => \N__12111\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_4\
        );

    \I__2569\ : CascadeMux
    port map (
            O => \N__12108\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4_cascade_\
        );

    \I__2568\ : CascadeMux
    port map (
            O => \N__12105\,
            I => \N__12102\
        );

    \I__2567\ : InMux
    port map (
            O => \N__12102\,
            I => \N__12099\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__12099\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_4\
        );

    \I__2565\ : InMux
    port map (
            O => \N__12096\,
            I => \N__12093\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__12093\,
            I => \N__12090\
        );

    \I__2563\ : Odrv12
    port map (
            O => \N__12090\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_5\
        );

    \I__2562\ : CascadeMux
    port map (
            O => \N__12087\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_\
        );

    \I__2561\ : CEMux
    port map (
            O => \N__12084\,
            I => \N__12080\
        );

    \I__2560\ : InMux
    port map (
            O => \N__12083\,
            I => \N__12077\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__12080\,
            I => \N__12074\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__12077\,
            I => \N__12071\
        );

    \I__2557\ : Span4Mux_v
    port map (
            O => \N__12074\,
            I => \N__12068\
        );

    \I__2556\ : Span4Mux_h
    port map (
            O => \N__12071\,
            I => \N__12065\
        );

    \I__2555\ : Span4Mux_h
    port map (
            O => \N__12068\,
            I => \N__12060\
        );

    \I__2554\ : Span4Mux_v
    port map (
            O => \N__12065\,
            I => \N__12060\
        );

    \I__2553\ : Odrv4
    port map (
            O => \N__12060\,
            I => \DUT.fifo_rx_inst.N_57\
        );

    \I__2552\ : InMux
    port map (
            O => \N__12057\,
            I => \N__12054\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__12054\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_6\
        );

    \I__2550\ : CascadeMux
    port map (
            O => \N__12051\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6_cascade_\
        );

    \I__2549\ : InMux
    port map (
            O => \N__12048\,
            I => \N__12045\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__12045\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_6\
        );

    \I__2547\ : InMux
    port map (
            O => \N__12042\,
            I => \N__12039\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__12039\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_7\
        );

    \I__2545\ : CascadeMux
    port map (
            O => \N__12036\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7_cascade_\
        );

    \I__2544\ : InMux
    port map (
            O => \N__12033\,
            I => \N__12030\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__12030\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_7\
        );

    \I__2542\ : InMux
    port map (
            O => \N__12027\,
            I => \N__12023\
        );

    \I__2541\ : InMux
    port map (
            O => \N__12026\,
            I => \N__12020\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__12023\,
            I => \N__12017\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__12020\,
            I => \DUT.fifo_rx_inst.rFifoDataro_3\
        );

    \I__2538\ : Odrv4
    port map (
            O => \N__12017\,
            I => \DUT.fifo_rx_inst.rFifoDataro_3\
        );

    \I__2537\ : InMux
    port map (
            O => \N__12012\,
            I => \N__12008\
        );

    \I__2536\ : InMux
    port map (
            O => \N__12011\,
            I => \N__12005\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__12008\,
            I => \N__12002\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__12005\,
            I => \DUT.fifo_tx_inst.rFifoDataro_0\
        );

    \I__2533\ : Odrv4
    port map (
            O => \N__12002\,
            I => \DUT.fifo_tx_inst.rFifoDataro_0\
        );

    \I__2532\ : CEMux
    port map (
            O => \N__11997\,
            I => \N__11994\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__11994\,
            I => \N__11990\
        );

    \I__2530\ : InMux
    port map (
            O => \N__11993\,
            I => \N__11987\
        );

    \I__2529\ : Span4Mux_v
    port map (
            O => \N__11990\,
            I => \N__11984\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__11987\,
            I => \N__11981\
        );

    \I__2527\ : Span4Mux_v
    port map (
            O => \N__11984\,
            I => \N__11978\
        );

    \I__2526\ : Span4Mux_h
    port map (
            O => \N__11981\,
            I => \N__11975\
        );

    \I__2525\ : Span4Mux_h
    port map (
            O => \N__11978\,
            I => \N__11972\
        );

    \I__2524\ : Span4Mux_v
    port map (
            O => \N__11975\,
            I => \N__11969\
        );

    \I__2523\ : Odrv4
    port map (
            O => \N__11972\,
            I => \DUT.fifo_tx_inst.rFifoData_awe1\
        );

    \I__2522\ : Odrv4
    port map (
            O => \N__11969\,
            I => \DUT.fifo_tx_inst.rFifoData_awe1\
        );

    \I__2521\ : CascadeMux
    port map (
            O => \N__11964\,
            I => \N__11960\
        );

    \I__2520\ : InMux
    port map (
            O => \N__11963\,
            I => \N__11957\
        );

    \I__2519\ : InMux
    port map (
            O => \N__11960\,
            I => \N__11954\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__11957\,
            I => \DUT.fifo_tx_inst.rFifoDataro_1\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__11954\,
            I => \DUT.fifo_tx_inst.rFifoDataro_1\
        );

    \I__2516\ : InMux
    port map (
            O => \N__11949\,
            I => \N__11945\
        );

    \I__2515\ : InMux
    port map (
            O => \N__11948\,
            I => \N__11942\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__11945\,
            I => \DUT.fifo_tx_inst.rFifoDataro_2\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__11942\,
            I => \DUT.fifo_tx_inst.rFifoDataro_2\
        );

    \I__2512\ : InMux
    port map (
            O => \N__11937\,
            I => \N__11933\
        );

    \I__2511\ : InMux
    port map (
            O => \N__11936\,
            I => \N__11930\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__11933\,
            I => \DUT.fifo_tx_inst.rFifoDataro_3\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__11930\,
            I => \DUT.fifo_tx_inst.rFifoDataro_3\
        );

    \I__2508\ : InMux
    port map (
            O => \N__11925\,
            I => \N__11922\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__11922\,
            I => \N__11919\
        );

    \I__2506\ : Span4Mux_h
    port map (
            O => \N__11919\,
            I => \N__11916\
        );

    \I__2505\ : Odrv4
    port map (
            O => \N__11916\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_0\
        );

    \I__2504\ : InMux
    port map (
            O => \N__11913\,
            I => \N__11910\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__11910\,
            I => \N__11907\
        );

    \I__2502\ : Span4Mux_h
    port map (
            O => \N__11907\,
            I => \N__11904\
        );

    \I__2501\ : Odrv4
    port map (
            O => \N__11904\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_1\
        );

    \I__2500\ : InMux
    port map (
            O => \N__11901\,
            I => \N__11898\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__11898\,
            I => \N__11895\
        );

    \I__2498\ : Odrv4
    port map (
            O => \N__11895\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_2\
        );

    \I__2497\ : InMux
    port map (
            O => \N__11892\,
            I => \N__11889\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__11889\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_3\
        );

    \I__2495\ : InMux
    port map (
            O => \N__11886\,
            I => \N__11883\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__11883\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_4\
        );

    \I__2493\ : InMux
    port map (
            O => \N__11880\,
            I => \N__11877\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__11877\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_5\
        );

    \I__2491\ : InMux
    port map (
            O => \N__11874\,
            I => \N__11871\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__11871\,
            I => \N__11868\
        );

    \I__2489\ : Odrv4
    port map (
            O => \N__11868\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_6\
        );

    \I__2488\ : InMux
    port map (
            O => \N__11865\,
            I => \N__11862\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__11862\,
            I => \N__11859\
        );

    \I__2486\ : Span4Mux_h
    port map (
            O => \N__11859\,
            I => \N__11856\
        );

    \I__2485\ : Odrv4
    port map (
            O => \N__11856\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_7\
        );

    \I__2484\ : CEMux
    port map (
            O => \N__11853\,
            I => \N__11849\
        );

    \I__2483\ : CEMux
    port map (
            O => \N__11852\,
            I => \N__11845\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__11849\,
            I => \N__11842\
        );

    \I__2481\ : CEMux
    port map (
            O => \N__11848\,
            I => \N__11839\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__11845\,
            I => \N__11835\
        );

    \I__2479\ : Span4Mux_s2_v
    port map (
            O => \N__11842\,
            I => \N__11829\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__11839\,
            I => \N__11829\
        );

    \I__2477\ : InMux
    port map (
            O => \N__11838\,
            I => \N__11826\
        );

    \I__2476\ : Span4Mux_v
    port map (
            O => \N__11835\,
            I => \N__11823\
        );

    \I__2475\ : CEMux
    port map (
            O => \N__11834\,
            I => \N__11820\
        );

    \I__2474\ : Span4Mux_v
    port map (
            O => \N__11829\,
            I => \N__11815\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__11826\,
            I => \N__11815\
        );

    \I__2472\ : Span4Mux_h
    port map (
            O => \N__11823\,
            I => \N__11812\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__11820\,
            I => \N__11809\
        );

    \I__2470\ : Span4Mux_h
    port map (
            O => \N__11815\,
            I => \N__11806\
        );

    \I__2469\ : Odrv4
    port map (
            O => \N__11812\,
            I => \DUT.fifo_tx_inst.rFifoData_awe0\
        );

    \I__2468\ : Odrv12
    port map (
            O => \N__11809\,
            I => \DUT.fifo_tx_inst.rFifoData_awe0\
        );

    \I__2467\ : Odrv4
    port map (
            O => \N__11806\,
            I => \DUT.fifo_tx_inst.rFifoData_awe0\
        );

    \I__2466\ : InMux
    port map (
            O => \N__11799\,
            I => \N__11796\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__11796\,
            I => \N__11793\
        );

    \I__2464\ : Odrv4
    port map (
            O => \N__11793\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_5\
        );

    \I__2463\ : CascadeMux
    port map (
            O => \N__11790\,
            I => \N__11787\
        );

    \I__2462\ : InMux
    port map (
            O => \N__11787\,
            I => \N__11784\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__11784\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_6\
        );

    \I__2460\ : InMux
    port map (
            O => \N__11781\,
            I => \N__11778\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__11778\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_7\
        );

    \I__2458\ : CascadeMux
    port map (
            O => \N__11775\,
            I => \N__11772\
        );

    \I__2457\ : InMux
    port map (
            O => \N__11772\,
            I => \N__11769\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__11769\,
            I => \N__11766\
        );

    \I__2455\ : Odrv4
    port map (
            O => \N__11766\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_2\
        );

    \I__2454\ : CascadeMux
    port map (
            O => \N__11763\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_\
        );

    \I__2453\ : InMux
    port map (
            O => \N__11760\,
            I => \N__11757\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__11757\,
            I => \N__11754\
        );

    \I__2451\ : Odrv4
    port map (
            O => \N__11754\,
            I => \DUT.rFifoDatarx_2\
        );

    \I__2450\ : InMux
    port map (
            O => \N__11751\,
            I => \N__11748\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__11748\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_2\
        );

    \I__2448\ : InMux
    port map (
            O => \N__11745\,
            I => \N__11732\
        );

    \I__2447\ : InMux
    port map (
            O => \N__11744\,
            I => \N__11732\
        );

    \I__2446\ : InMux
    port map (
            O => \N__11743\,
            I => \N__11732\
        );

    \I__2445\ : InMux
    port map (
            O => \N__11742\,
            I => \N__11723\
        );

    \I__2444\ : InMux
    port map (
            O => \N__11741\,
            I => \N__11716\
        );

    \I__2443\ : InMux
    port map (
            O => \N__11740\,
            I => \N__11716\
        );

    \I__2442\ : InMux
    port map (
            O => \N__11739\,
            I => \N__11716\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__11732\,
            I => \N__11713\
        );

    \I__2440\ : InMux
    port map (
            O => \N__11731\,
            I => \N__11708\
        );

    \I__2439\ : InMux
    port map (
            O => \N__11730\,
            I => \N__11708\
        );

    \I__2438\ : InMux
    port map (
            O => \N__11729\,
            I => \N__11699\
        );

    \I__2437\ : InMux
    port map (
            O => \N__11728\,
            I => \N__11699\
        );

    \I__2436\ : InMux
    port map (
            O => \N__11727\,
            I => \N__11699\
        );

    \I__2435\ : InMux
    port map (
            O => \N__11726\,
            I => \N__11699\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__11723\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__11716\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__2432\ : Odrv4
    port map (
            O => \N__11713\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__11708\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__11699\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__2429\ : InMux
    port map (
            O => \N__11688\,
            I => \N__11685\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__11685\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_3\
        );

    \I__2427\ : CascadeMux
    port map (
            O => \N__11682\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_\
        );

    \I__2426\ : CascadeMux
    port map (
            O => \N__11679\,
            I => \N__11670\
        );

    \I__2425\ : CascadeMux
    port map (
            O => \N__11678\,
            I => \N__11667\
        );

    \I__2424\ : CascadeMux
    port map (
            O => \N__11677\,
            I => \N__11659\
        );

    \I__2423\ : CascadeMux
    port map (
            O => \N__11676\,
            I => \N__11651\
        );

    \I__2422\ : InMux
    port map (
            O => \N__11675\,
            I => \N__11638\
        );

    \I__2421\ : InMux
    port map (
            O => \N__11674\,
            I => \N__11638\
        );

    \I__2420\ : InMux
    port map (
            O => \N__11673\,
            I => \N__11638\
        );

    \I__2419\ : InMux
    port map (
            O => \N__11670\,
            I => \N__11638\
        );

    \I__2418\ : InMux
    port map (
            O => \N__11667\,
            I => \N__11638\
        );

    \I__2417\ : InMux
    port map (
            O => \N__11666\,
            I => \N__11638\
        );

    \I__2416\ : CascadeMux
    port map (
            O => \N__11665\,
            I => \N__11632\
        );

    \I__2415\ : InMux
    port map (
            O => \N__11664\,
            I => \N__11619\
        );

    \I__2414\ : InMux
    port map (
            O => \N__11663\,
            I => \N__11619\
        );

    \I__2413\ : InMux
    port map (
            O => \N__11662\,
            I => \N__11619\
        );

    \I__2412\ : InMux
    port map (
            O => \N__11659\,
            I => \N__11619\
        );

    \I__2411\ : InMux
    port map (
            O => \N__11658\,
            I => \N__11619\
        );

    \I__2410\ : InMux
    port map (
            O => \N__11657\,
            I => \N__11619\
        );

    \I__2409\ : InMux
    port map (
            O => \N__11656\,
            I => \N__11610\
        );

    \I__2408\ : InMux
    port map (
            O => \N__11655\,
            I => \N__11610\
        );

    \I__2407\ : InMux
    port map (
            O => \N__11654\,
            I => \N__11610\
        );

    \I__2406\ : InMux
    port map (
            O => \N__11651\,
            I => \N__11610\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__11638\,
            I => \N__11607\
        );

    \I__2404\ : InMux
    port map (
            O => \N__11637\,
            I => \N__11598\
        );

    \I__2403\ : InMux
    port map (
            O => \N__11636\,
            I => \N__11598\
        );

    \I__2402\ : InMux
    port map (
            O => \N__11635\,
            I => \N__11598\
        );

    \I__2401\ : InMux
    port map (
            O => \N__11632\,
            I => \N__11598\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__11619\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__11610\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__2398\ : Odrv4
    port map (
            O => \N__11607\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__11598\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__2396\ : InMux
    port map (
            O => \N__11589\,
            I => \N__11586\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__11586\,
            I => \N__11583\
        );

    \I__2394\ : Odrv12
    port map (
            O => \N__11583\,
            I => \DUT.rFifoDatarx_3\
        );

    \I__2393\ : InMux
    port map (
            O => \N__11580\,
            I => \N__11577\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__11577\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_3\
        );

    \I__2391\ : CascadeMux
    port map (
            O => \N__11574\,
            I => \N__11569\
        );

    \I__2390\ : CascadeMux
    port map (
            O => \N__11573\,
            I => \N__11565\
        );

    \I__2389\ : CascadeMux
    port map (
            O => \N__11572\,
            I => \N__11559\
        );

    \I__2388\ : InMux
    port map (
            O => \N__11569\,
            I => \N__11552\
        );

    \I__2387\ : InMux
    port map (
            O => \N__11568\,
            I => \N__11552\
        );

    \I__2386\ : InMux
    port map (
            O => \N__11565\,
            I => \N__11552\
        );

    \I__2385\ : InMux
    port map (
            O => \N__11564\,
            I => \N__11549\
        );

    \I__2384\ : InMux
    port map (
            O => \N__11563\,
            I => \N__11539\
        );

    \I__2383\ : InMux
    port map (
            O => \N__11562\,
            I => \N__11539\
        );

    \I__2382\ : InMux
    port map (
            O => \N__11559\,
            I => \N__11536\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__11552\,
            I => \N__11533\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__11549\,
            I => \N__11530\
        );

    \I__2379\ : InMux
    port map (
            O => \N__11548\,
            I => \N__11523\
        );

    \I__2378\ : InMux
    port map (
            O => \N__11547\,
            I => \N__11523\
        );

    \I__2377\ : InMux
    port map (
            O => \N__11546\,
            I => \N__11523\
        );

    \I__2376\ : InMux
    port map (
            O => \N__11545\,
            I => \N__11520\
        );

    \I__2375\ : InMux
    port map (
            O => \N__11544\,
            I => \N__11517\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__11539\,
            I => \N__11510\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__11536\,
            I => \N__11510\
        );

    \I__2372\ : Span4Mux_h
    port map (
            O => \N__11533\,
            I => \N__11510\
        );

    \I__2371\ : Odrv12
    port map (
            O => \N__11530\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_5\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__11523\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_5\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__11520\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_5\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__11517\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_5\
        );

    \I__2367\ : Odrv4
    port map (
            O => \N__11510\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_5\
        );

    \I__2366\ : CascadeMux
    port map (
            O => \N__11499\,
            I => \N__11494\
        );

    \I__2365\ : InMux
    port map (
            O => \N__11498\,
            I => \N__11484\
        );

    \I__2364\ : CascadeMux
    port map (
            O => \N__11497\,
            I => \N__11481\
        );

    \I__2363\ : InMux
    port map (
            O => \N__11494\,
            I => \N__11475\
        );

    \I__2362\ : InMux
    port map (
            O => \N__11493\,
            I => \N__11475\
        );

    \I__2361\ : InMux
    port map (
            O => \N__11492\,
            I => \N__11468\
        );

    \I__2360\ : InMux
    port map (
            O => \N__11491\,
            I => \N__11468\
        );

    \I__2359\ : InMux
    port map (
            O => \N__11490\,
            I => \N__11468\
        );

    \I__2358\ : InMux
    port map (
            O => \N__11489\,
            I => \N__11462\
        );

    \I__2357\ : InMux
    port map (
            O => \N__11488\,
            I => \N__11462\
        );

    \I__2356\ : CascadeMux
    port map (
            O => \N__11487\,
            I => \N__11459\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__11484\,
            I => \N__11456\
        );

    \I__2354\ : InMux
    port map (
            O => \N__11481\,
            I => \N__11452\
        );

    \I__2353\ : InMux
    port map (
            O => \N__11480\,
            I => \N__11449\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__11475\,
            I => \N__11444\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__11468\,
            I => \N__11444\
        );

    \I__2350\ : CascadeMux
    port map (
            O => \N__11467\,
            I => \N__11441\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__11462\,
            I => \N__11438\
        );

    \I__2348\ : InMux
    port map (
            O => \N__11459\,
            I => \N__11435\
        );

    \I__2347\ : Span4Mux_v
    port map (
            O => \N__11456\,
            I => \N__11432\
        );

    \I__2346\ : InMux
    port map (
            O => \N__11455\,
            I => \N__11429\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__11452\,
            I => \N__11426\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__11449\,
            I => \N__11421\
        );

    \I__2343\ : Span4Mux_v
    port map (
            O => \N__11444\,
            I => \N__11421\
        );

    \I__2342\ : InMux
    port map (
            O => \N__11441\,
            I => \N__11418\
        );

    \I__2341\ : Span4Mux_v
    port map (
            O => \N__11438\,
            I => \N__11415\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__11435\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_4\
        );

    \I__2339\ : Odrv4
    port map (
            O => \N__11432\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_4\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__11429\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_4\
        );

    \I__2337\ : Odrv4
    port map (
            O => \N__11426\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_4\
        );

    \I__2336\ : Odrv4
    port map (
            O => \N__11421\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_4\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__11418\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_4\
        );

    \I__2334\ : Odrv4
    port map (
            O => \N__11415\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_4\
        );

    \I__2333\ : InMux
    port map (
            O => \N__11400\,
            I => \N__11394\
        );

    \I__2332\ : InMux
    port map (
            O => \N__11399\,
            I => \N__11389\
        );

    \I__2331\ : InMux
    port map (
            O => \N__11398\,
            I => \N__11384\
        );

    \I__2330\ : InMux
    port map (
            O => \N__11397\,
            I => \N__11384\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__11394\,
            I => \N__11381\
        );

    \I__2328\ : CascadeMux
    port map (
            O => \N__11393\,
            I => \N__11374\
        );

    \I__2327\ : InMux
    port map (
            O => \N__11392\,
            I => \N__11371\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__11389\,
            I => \N__11368\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__11384\,
            I => \N__11363\
        );

    \I__2324\ : Span4Mux_h
    port map (
            O => \N__11381\,
            I => \N__11363\
        );

    \I__2323\ : InMux
    port map (
            O => \N__11380\,
            I => \N__11356\
        );

    \I__2322\ : InMux
    port map (
            O => \N__11379\,
            I => \N__11356\
        );

    \I__2321\ : InMux
    port map (
            O => \N__11378\,
            I => \N__11356\
        );

    \I__2320\ : InMux
    port map (
            O => \N__11377\,
            I => \N__11353\
        );

    \I__2319\ : InMux
    port map (
            O => \N__11374\,
            I => \N__11350\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__11371\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_1\
        );

    \I__2317\ : Odrv4
    port map (
            O => \N__11368\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_1\
        );

    \I__2316\ : Odrv4
    port map (
            O => \N__11363\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_1\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__11356\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_1\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__11353\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_1\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__11350\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_1\
        );

    \I__2312\ : InMux
    port map (
            O => \N__11337\,
            I => \N__11333\
        );

    \I__2311\ : CascadeMux
    port map (
            O => \N__11336\,
            I => \N__11329\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__11333\,
            I => \N__11326\
        );

    \I__2309\ : InMux
    port map (
            O => \N__11332\,
            I => \N__11323\
        );

    \I__2308\ : InMux
    port map (
            O => \N__11329\,
            I => \N__11318\
        );

    \I__2307\ : Span4Mux_v
    port map (
            O => \N__11326\,
            I => \N__11313\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__11323\,
            I => \N__11313\
        );

    \I__2305\ : InMux
    port map (
            O => \N__11322\,
            I => \N__11308\
        );

    \I__2304\ : InMux
    port map (
            O => \N__11321\,
            I => \N__11308\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__11318\,
            I => \DUT.uart_inst0.recv_stateZ0Z_3\
        );

    \I__2302\ : Odrv4
    port map (
            O => \N__11313\,
            I => \DUT.uart_inst0.recv_stateZ0Z_3\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__11308\,
            I => \DUT.uart_inst0.recv_stateZ0Z_3\
        );

    \I__2300\ : InMux
    port map (
            O => \N__11301\,
            I => \N__11298\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__11298\,
            I => \N__11295\
        );

    \I__2298\ : Span4Mux_v
    port map (
            O => \N__11295\,
            I => \N__11292\
        );

    \I__2297\ : Odrv4
    port map (
            O => \N__11292\,
            I => \DUT.uart_inst0.m6_e_2\
        );

    \I__2296\ : CascadeMux
    port map (
            O => \N__11289\,
            I => \DUT.uart_inst0.m6_e_3_cascade_\
        );

    \I__2295\ : InMux
    port map (
            O => \N__11286\,
            I => \N__11282\
        );

    \I__2294\ : InMux
    port map (
            O => \N__11285\,
            I => \N__11279\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__11282\,
            I => \N__11276\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__11279\,
            I => \DUT.uart_inst0.N_15_mux\
        );

    \I__2291\ : Odrv4
    port map (
            O => \N__11276\,
            I => \DUT.uart_inst0.N_15_mux\
        );

    \I__2290\ : InMux
    port map (
            O => \N__11271\,
            I => \N__11268\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__11268\,
            I => \DUT.uart_inst0.N_18_mux_1\
        );

    \I__2288\ : CascadeMux
    port map (
            O => \N__11265\,
            I => \N__11258\
        );

    \I__2287\ : InMux
    port map (
            O => \N__11264\,
            I => \N__11251\
        );

    \I__2286\ : InMux
    port map (
            O => \N__11263\,
            I => \N__11251\
        );

    \I__2285\ : InMux
    port map (
            O => \N__11262\,
            I => \N__11246\
        );

    \I__2284\ : InMux
    port map (
            O => \N__11261\,
            I => \N__11246\
        );

    \I__2283\ : InMux
    port map (
            O => \N__11258\,
            I => \N__11241\
        );

    \I__2282\ : InMux
    port map (
            O => \N__11257\,
            I => \N__11238\
        );

    \I__2281\ : InMux
    port map (
            O => \N__11256\,
            I => \N__11235\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__11251\,
            I => \N__11230\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__11246\,
            I => \N__11230\
        );

    \I__2278\ : InMux
    port map (
            O => \N__11245\,
            I => \N__11225\
        );

    \I__2277\ : InMux
    port map (
            O => \N__11244\,
            I => \N__11225\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__11241\,
            I => \N__11221\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__11238\,
            I => \N__11213\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__11235\,
            I => \N__11213\
        );

    \I__2273\ : Span4Mux_h
    port map (
            O => \N__11230\,
            I => \N__11208\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__11225\,
            I => \N__11208\
        );

    \I__2271\ : CascadeMux
    port map (
            O => \N__11224\,
            I => \N__11205\
        );

    \I__2270\ : Span4Mux_v
    port map (
            O => \N__11221\,
            I => \N__11202\
        );

    \I__2269\ : InMux
    port map (
            O => \N__11220\,
            I => \N__11197\
        );

    \I__2268\ : InMux
    port map (
            O => \N__11219\,
            I => \N__11197\
        );

    \I__2267\ : InMux
    port map (
            O => \N__11218\,
            I => \N__11194\
        );

    \I__2266\ : Span4Mux_v
    port map (
            O => \N__11213\,
            I => \N__11189\
        );

    \I__2265\ : Span4Mux_v
    port map (
            O => \N__11208\,
            I => \N__11189\
        );

    \I__2264\ : InMux
    port map (
            O => \N__11205\,
            I => \N__11186\
        );

    \I__2263\ : Odrv4
    port map (
            O => \N__11202\,
            I => \DUT.uart_inst0.rx_countdownZ1Z_3\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__11197\,
            I => \DUT.uart_inst0.rx_countdownZ1Z_3\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__11194\,
            I => \DUT.uart_inst0.rx_countdownZ1Z_3\
        );

    \I__2260\ : Odrv4
    port map (
            O => \N__11189\,
            I => \DUT.uart_inst0.rx_countdownZ1Z_3\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__11186\,
            I => \DUT.uart_inst0.rx_countdownZ1Z_3\
        );

    \I__2258\ : InMux
    port map (
            O => \N__11175\,
            I => \N__11170\
        );

    \I__2257\ : InMux
    port map (
            O => \N__11174\,
            I => \N__11167\
        );

    \I__2256\ : InMux
    port map (
            O => \N__11173\,
            I => \N__11164\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__11170\,
            I => \DUT.uart_inst0.recv_stateZ0Z_4\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__11167\,
            I => \DUT.uart_inst0.recv_stateZ0Z_4\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__11164\,
            I => \DUT.uart_inst0.recv_stateZ0Z_4\
        );

    \I__2252\ : InMux
    port map (
            O => \N__11157\,
            I => \N__11150\
        );

    \I__2251\ : CascadeMux
    port map (
            O => \N__11156\,
            I => \N__11146\
        );

    \I__2250\ : InMux
    port map (
            O => \N__11155\,
            I => \N__11141\
        );

    \I__2249\ : InMux
    port map (
            O => \N__11154\,
            I => \N__11141\
        );

    \I__2248\ : InMux
    port map (
            O => \N__11153\,
            I => \N__11136\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__11150\,
            I => \N__11133\
        );

    \I__2246\ : InMux
    port map (
            O => \N__11149\,
            I => \N__11128\
        );

    \I__2245\ : InMux
    port map (
            O => \N__11146\,
            I => \N__11128\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__11141\,
            I => \N__11125\
        );

    \I__2243\ : InMux
    port map (
            O => \N__11140\,
            I => \N__11120\
        );

    \I__2242\ : InMux
    port map (
            O => \N__11139\,
            I => \N__11120\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__11136\,
            I => \N__11109\
        );

    \I__2240\ : Span4Mux_v
    port map (
            O => \N__11133\,
            I => \N__11109\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__11128\,
            I => \N__11109\
        );

    \I__2238\ : Span4Mux_h
    port map (
            O => \N__11125\,
            I => \N__11104\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__11120\,
            I => \N__11104\
        );

    \I__2236\ : InMux
    port map (
            O => \N__11119\,
            I => \N__11095\
        );

    \I__2235\ : InMux
    port map (
            O => \N__11118\,
            I => \N__11095\
        );

    \I__2234\ : InMux
    port map (
            O => \N__11117\,
            I => \N__11095\
        );

    \I__2233\ : InMux
    port map (
            O => \N__11116\,
            I => \N__11095\
        );

    \I__2232\ : Span4Mux_h
    port map (
            O => \N__11109\,
            I => \N__11092\
        );

    \I__2231\ : Odrv4
    port map (
            O => \N__11104\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_2\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__11095\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_2\
        );

    \I__2229\ : Odrv4
    port map (
            O => \N__11092\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_2\
        );

    \I__2228\ : CascadeMux
    port map (
            O => \N__11085\,
            I => \N__11082\
        );

    \I__2227\ : InMux
    port map (
            O => \N__11082\,
            I => \N__11079\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__11079\,
            I => \N__11076\
        );

    \I__2225\ : Odrv4
    port map (
            O => \N__11076\,
            I => \DUT.uart_inst0.G_19_0_a5_2\
        );

    \I__2224\ : CascadeMux
    port map (
            O => \N__11073\,
            I => \N__11070\
        );

    \I__2223\ : InMux
    port map (
            O => \N__11070\,
            I => \N__11067\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__11067\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_0\
        );

    \I__2221\ : InMux
    port map (
            O => \N__11064\,
            I => \N__11061\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__11061\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_1\
        );

    \I__2219\ : CascadeMux
    port map (
            O => \N__11058\,
            I => \N__11055\
        );

    \I__2218\ : InMux
    port map (
            O => \N__11055\,
            I => \N__11052\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__11052\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_4\
        );

    \I__2216\ : InMux
    port map (
            O => \N__11049\,
            I => \N__11043\
        );

    \I__2215\ : InMux
    port map (
            O => \N__11048\,
            I => \N__11043\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__11043\,
            I => \DUT.fifo_rx_inst.N_77_mux\
        );

    \I__2213\ : InMux
    port map (
            O => \N__11040\,
            I => \N__11036\
        );

    \I__2212\ : InMux
    port map (
            O => \N__11039\,
            I => \N__11032\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__11036\,
            I => \N__11029\
        );

    \I__2210\ : InMux
    port map (
            O => \N__11035\,
            I => \N__11026\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__11032\,
            I => \N__11023\
        );

    \I__2208\ : Odrv4
    port map (
            O => \N__11029\,
            I => \DUT.uart_inst0.g1_0\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__11026\,
            I => \DUT.uart_inst0.g1_0\
        );

    \I__2206\ : Odrv4
    port map (
            O => \N__11023\,
            I => \DUT.uart_inst0.g1_0\
        );

    \I__2205\ : CascadeMux
    port map (
            O => \N__11016\,
            I => \N__11006\
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__11015\,
            I => \N__11001\
        );

    \I__2203\ : CascadeMux
    port map (
            O => \N__11014\,
            I => \N__10998\
        );

    \I__2202\ : InMux
    port map (
            O => \N__11013\,
            I => \N__10990\
        );

    \I__2201\ : InMux
    port map (
            O => \N__11012\,
            I => \N__10985\
        );

    \I__2200\ : InMux
    port map (
            O => \N__11011\,
            I => \N__10985\
        );

    \I__2199\ : InMux
    port map (
            O => \N__11010\,
            I => \N__10976\
        );

    \I__2198\ : InMux
    port map (
            O => \N__11009\,
            I => \N__10976\
        );

    \I__2197\ : InMux
    port map (
            O => \N__11006\,
            I => \N__10976\
        );

    \I__2196\ : InMux
    port map (
            O => \N__11005\,
            I => \N__10976\
        );

    \I__2195\ : InMux
    port map (
            O => \N__11004\,
            I => \N__10961\
        );

    \I__2194\ : InMux
    port map (
            O => \N__11001\,
            I => \N__10961\
        );

    \I__2193\ : InMux
    port map (
            O => \N__10998\,
            I => \N__10961\
        );

    \I__2192\ : InMux
    port map (
            O => \N__10997\,
            I => \N__10961\
        );

    \I__2191\ : InMux
    port map (
            O => \N__10996\,
            I => \N__10961\
        );

    \I__2190\ : InMux
    port map (
            O => \N__10995\,
            I => \N__10961\
        );

    \I__2189\ : InMux
    port map (
            O => \N__10994\,
            I => \N__10961\
        );

    \I__2188\ : CascadeMux
    port map (
            O => \N__10993\,
            I => \N__10956\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__10990\,
            I => \N__10949\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__10985\,
            I => \N__10946\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__10976\,
            I => \N__10941\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__10961\,
            I => \N__10941\
        );

    \I__2183\ : InMux
    port map (
            O => \N__10960\,
            I => \N__10928\
        );

    \I__2182\ : InMux
    port map (
            O => \N__10959\,
            I => \N__10928\
        );

    \I__2181\ : InMux
    port map (
            O => \N__10956\,
            I => \N__10928\
        );

    \I__2180\ : InMux
    port map (
            O => \N__10955\,
            I => \N__10928\
        );

    \I__2179\ : InMux
    port map (
            O => \N__10954\,
            I => \N__10928\
        );

    \I__2178\ : InMux
    port map (
            O => \N__10953\,
            I => \N__10928\
        );

    \I__2177\ : InMux
    port map (
            O => \N__10952\,
            I => \N__10922\
        );

    \I__2176\ : Span4Mux_h
    port map (
            O => \N__10949\,
            I => \N__10919\
        );

    \I__2175\ : Span4Mux_h
    port map (
            O => \N__10946\,
            I => \N__10916\
        );

    \I__2174\ : Span4Mux_v
    port map (
            O => \N__10941\,
            I => \N__10913\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__10928\,
            I => \N__10910\
        );

    \I__2172\ : InMux
    port map (
            O => \N__10927\,
            I => \N__10903\
        );

    \I__2171\ : InMux
    port map (
            O => \N__10926\,
            I => \N__10903\
        );

    \I__2170\ : InMux
    port map (
            O => \N__10925\,
            I => \N__10903\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__10922\,
            I => \DUT.uart_inst0.recv_stateZ0Z_0\
        );

    \I__2168\ : Odrv4
    port map (
            O => \N__10919\,
            I => \DUT.uart_inst0.recv_stateZ0Z_0\
        );

    \I__2167\ : Odrv4
    port map (
            O => \N__10916\,
            I => \DUT.uart_inst0.recv_stateZ0Z_0\
        );

    \I__2166\ : Odrv4
    port map (
            O => \N__10913\,
            I => \DUT.uart_inst0.recv_stateZ0Z_0\
        );

    \I__2165\ : Odrv4
    port map (
            O => \N__10910\,
            I => \DUT.uart_inst0.recv_stateZ0Z_0\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__10903\,
            I => \DUT.uart_inst0.recv_stateZ0Z_0\
        );

    \I__2163\ : CascadeMux
    port map (
            O => \N__10890\,
            I => \N__10886\
        );

    \I__2162\ : InMux
    port map (
            O => \N__10889\,
            I => \N__10883\
        );

    \I__2161\ : InMux
    port map (
            O => \N__10886\,
            I => \N__10880\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__10883\,
            I => \N__10873\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__10880\,
            I => \N__10870\
        );

    \I__2158\ : InMux
    port map (
            O => \N__10879\,
            I => \N__10865\
        );

    \I__2157\ : InMux
    port map (
            O => \N__10878\,
            I => \N__10865\
        );

    \I__2156\ : InMux
    port map (
            O => \N__10877\,
            I => \N__10860\
        );

    \I__2155\ : InMux
    port map (
            O => \N__10876\,
            I => \N__10860\
        );

    \I__2154\ : Odrv4
    port map (
            O => \N__10873\,
            I => \DUT.uart_inst0.recv_stateZ0Z_5\
        );

    \I__2153\ : Odrv4
    port map (
            O => \N__10870\,
            I => \DUT.uart_inst0.recv_stateZ0Z_5\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__10865\,
            I => \DUT.uart_inst0.recv_stateZ0Z_5\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__10860\,
            I => \DUT.uart_inst0.recv_stateZ0Z_5\
        );

    \I__2150\ : CascadeMux
    port map (
            O => \N__10851\,
            I => \N__10848\
        );

    \I__2149\ : InMux
    port map (
            O => \N__10848\,
            I => \N__10845\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__10845\,
            I => \N__10842\
        );

    \I__2147\ : Span4Mux_v
    port map (
            O => \N__10842\,
            I => \N__10839\
        );

    \I__2146\ : Odrv4
    port map (
            O => \N__10839\,
            I => \DUT.uart_inst0.rx_countdown_8_i_a2_0_2\
        );

    \I__2145\ : InMux
    port map (
            O => \N__10836\,
            I => \N__10833\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__10833\,
            I => \DUT.uart_inst0.m10_e_3\
        );

    \I__2143\ : InMux
    port map (
            O => \N__10830\,
            I => \N__10827\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__10827\,
            I => \DUT.uart_inst0.m10_e_2\
        );

    \I__2141\ : InMux
    port map (
            O => \N__10824\,
            I => \N__10818\
        );

    \I__2140\ : CascadeMux
    port map (
            O => \N__10823\,
            I => \N__10815\
        );

    \I__2139\ : IoInMux
    port map (
            O => \N__10822\,
            I => \N__10809\
        );

    \I__2138\ : InMux
    port map (
            O => \N__10821\,
            I => \N__10806\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__10818\,
            I => \N__10803\
        );

    \I__2136\ : InMux
    port map (
            O => \N__10815\,
            I => \N__10800\
        );

    \I__2135\ : InMux
    port map (
            O => \N__10814\,
            I => \N__10795\
        );

    \I__2134\ : InMux
    port map (
            O => \N__10813\,
            I => \N__10795\
        );

    \I__2133\ : InMux
    port map (
            O => \N__10812\,
            I => \N__10792\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__10809\,
            I => \N__10788\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__10806\,
            I => \N__10784\
        );

    \I__2130\ : Span4Mux_v
    port map (
            O => \N__10803\,
            I => \N__10779\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__10800\,
            I => \N__10779\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__10795\,
            I => \N__10776\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__10792\,
            I => \N__10773\
        );

    \I__2126\ : InMux
    port map (
            O => \N__10791\,
            I => \N__10770\
        );

    \I__2125\ : Span4Mux_s1_v
    port map (
            O => \N__10788\,
            I => \N__10767\
        );

    \I__2124\ : InMux
    port map (
            O => \N__10787\,
            I => \N__10764\
        );

    \I__2123\ : Span4Mux_v
    port map (
            O => \N__10784\,
            I => \N__10759\
        );

    \I__2122\ : Span4Mux_v
    port map (
            O => \N__10779\,
            I => \N__10759\
        );

    \I__2121\ : Span4Mux_h
    port map (
            O => \N__10776\,
            I => \N__10752\
        );

    \I__2120\ : Span4Mux_v
    port map (
            O => \N__10773\,
            I => \N__10752\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__10770\,
            I => \N__10752\
        );

    \I__2118\ : Span4Mux_v
    port map (
            O => \N__10767\,
            I => \N__10749\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__10764\,
            I => \N__10746\
        );

    \I__2116\ : Sp12to4
    port map (
            O => \N__10759\,
            I => \N__10743\
        );

    \I__2115\ : Span4Mux_v
    port map (
            O => \N__10752\,
            I => \N__10740\
        );

    \I__2114\ : Sp12to4
    port map (
            O => \N__10749\,
            I => \N__10735\
        );

    \I__2113\ : Span12Mux_s5_v
    port map (
            O => \N__10746\,
            I => \N__10735\
        );

    \I__2112\ : Span12Mux_h
    port map (
            O => \N__10743\,
            I => \N__10730\
        );

    \I__2111\ : Sp12to4
    port map (
            O => \N__10740\,
            I => \N__10730\
        );

    \I__2110\ : Span12Mux_h
    port map (
            O => \N__10735\,
            I => \N__10727\
        );

    \I__2109\ : Span12Mux_h
    port map (
            O => \N__10730\,
            I => \N__10724\
        );

    \I__2108\ : Span12Mux_v
    port map (
            O => \N__10727\,
            I => \N__10721\
        );

    \I__2107\ : Span12Mux_v
    port map (
            O => \N__10724\,
            I => \N__10718\
        );

    \I__2106\ : Odrv12
    port map (
            O => \N__10721\,
            I => \wPllLocked\
        );

    \I__2105\ : Odrv12
    port map (
            O => \N__10718\,
            I => \wPllLocked\
        );

    \I__2104\ : CascadeMux
    port map (
            O => \N__10713\,
            I => \DUT.uart_inst0.N_20_mux_cascade_\
        );

    \I__2103\ : InMux
    port map (
            O => \N__10710\,
            I => \N__10703\
        );

    \I__2102\ : CascadeMux
    port map (
            O => \N__10709\,
            I => \N__10696\
        );

    \I__2101\ : InMux
    port map (
            O => \N__10708\,
            I => \N__10687\
        );

    \I__2100\ : InMux
    port map (
            O => \N__10707\,
            I => \N__10687\
        );

    \I__2099\ : CascadeMux
    port map (
            O => \N__10706\,
            I => \N__10679\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__10703\,
            I => \N__10672\
        );

    \I__2097\ : InMux
    port map (
            O => \N__10702\,
            I => \N__10667\
        );

    \I__2096\ : InMux
    port map (
            O => \N__10701\,
            I => \N__10667\
        );

    \I__2095\ : InMux
    port map (
            O => \N__10700\,
            I => \N__10664\
        );

    \I__2094\ : InMux
    port map (
            O => \N__10699\,
            I => \N__10659\
        );

    \I__2093\ : InMux
    port map (
            O => \N__10696\,
            I => \N__10659\
        );

    \I__2092\ : InMux
    port map (
            O => \N__10695\,
            I => \N__10656\
        );

    \I__2091\ : InMux
    port map (
            O => \N__10694\,
            I => \N__10653\
        );

    \I__2090\ : InMux
    port map (
            O => \N__10693\,
            I => \N__10648\
        );

    \I__2089\ : InMux
    port map (
            O => \N__10692\,
            I => \N__10648\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__10687\,
            I => \N__10645\
        );

    \I__2087\ : InMux
    port map (
            O => \N__10686\,
            I => \N__10642\
        );

    \I__2086\ : InMux
    port map (
            O => \N__10685\,
            I => \N__10637\
        );

    \I__2085\ : InMux
    port map (
            O => \N__10684\,
            I => \N__10637\
        );

    \I__2084\ : InMux
    port map (
            O => \N__10683\,
            I => \N__10632\
        );

    \I__2083\ : InMux
    port map (
            O => \N__10682\,
            I => \N__10632\
        );

    \I__2082\ : InMux
    port map (
            O => \N__10679\,
            I => \N__10627\
        );

    \I__2081\ : InMux
    port map (
            O => \N__10678\,
            I => \N__10627\
        );

    \I__2080\ : InMux
    port map (
            O => \N__10677\,
            I => \N__10622\
        );

    \I__2079\ : InMux
    port map (
            O => \N__10676\,
            I => \N__10622\
        );

    \I__2078\ : InMux
    port map (
            O => \N__10675\,
            I => \N__10619\
        );

    \I__2077\ : Span4Mux_v
    port map (
            O => \N__10672\,
            I => \N__10608\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__10667\,
            I => \N__10608\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__10664\,
            I => \N__10608\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__10659\,
            I => \N__10608\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__10656\,
            I => \N__10608\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__10653\,
            I => \N__10603\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__10648\,
            I => \N__10603\
        );

    \I__2070\ : Span4Mux_v
    port map (
            O => \N__10645\,
            I => \N__10600\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__10642\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__10637\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__10632\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__10627\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__10622\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__10619\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__2063\ : Odrv4
    port map (
            O => \N__10608\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__2062\ : Odrv4
    port map (
            O => \N__10603\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__2061\ : Odrv4
    port map (
            O => \N__10600\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__2060\ : CascadeMux
    port map (
            O => \N__10581\,
            I => \DUT.uart_inst0.m7_3_cascade_\
        );

    \I__2059\ : InMux
    port map (
            O => \N__10578\,
            I => \N__10575\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__10575\,
            I => \N__10572\
        );

    \I__2057\ : Odrv12
    port map (
            O => \N__10572\,
            I => \DUT.uart_inst0.N_28_mux\
        );

    \I__2056\ : CascadeMux
    port map (
            O => \N__10569\,
            I => \N__10552\
        );

    \I__2055\ : CascadeMux
    port map (
            O => \N__10568\,
            I => \N__10549\
        );

    \I__2054\ : CascadeMux
    port map (
            O => \N__10567\,
            I => \N__10544\
        );

    \I__2053\ : InMux
    port map (
            O => \N__10566\,
            I => \N__10537\
        );

    \I__2052\ : InMux
    port map (
            O => \N__10565\,
            I => \N__10537\
        );

    \I__2051\ : InMux
    port map (
            O => \N__10564\,
            I => \N__10537\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__10563\,
            I => \N__10532\
        );

    \I__2049\ : CascadeMux
    port map (
            O => \N__10562\,
            I => \N__10528\
        );

    \I__2048\ : CascadeMux
    port map (
            O => \N__10561\,
            I => \N__10523\
        );

    \I__2047\ : CascadeMux
    port map (
            O => \N__10560\,
            I => \N__10520\
        );

    \I__2046\ : CascadeMux
    port map (
            O => \N__10559\,
            I => \N__10514\
        );

    \I__2045\ : CascadeMux
    port map (
            O => \N__10558\,
            I => \N__10510\
        );

    \I__2044\ : CascadeMux
    port map (
            O => \N__10557\,
            I => \N__10506\
        );

    \I__2043\ : InMux
    port map (
            O => \N__10556\,
            I => \N__10499\
        );

    \I__2042\ : InMux
    port map (
            O => \N__10555\,
            I => \N__10494\
        );

    \I__2041\ : InMux
    port map (
            O => \N__10552\,
            I => \N__10494\
        );

    \I__2040\ : InMux
    port map (
            O => \N__10549\,
            I => \N__10491\
        );

    \I__2039\ : InMux
    port map (
            O => \N__10548\,
            I => \N__10488\
        );

    \I__2038\ : InMux
    port map (
            O => \N__10547\,
            I => \N__10483\
        );

    \I__2037\ : InMux
    port map (
            O => \N__10544\,
            I => \N__10483\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__10537\,
            I => \N__10479\
        );

    \I__2035\ : InMux
    port map (
            O => \N__10536\,
            I => \N__10474\
        );

    \I__2034\ : InMux
    port map (
            O => \N__10535\,
            I => \N__10474\
        );

    \I__2033\ : InMux
    port map (
            O => \N__10532\,
            I => \N__10463\
        );

    \I__2032\ : InMux
    port map (
            O => \N__10531\,
            I => \N__10463\
        );

    \I__2031\ : InMux
    port map (
            O => \N__10528\,
            I => \N__10463\
        );

    \I__2030\ : InMux
    port map (
            O => \N__10527\,
            I => \N__10463\
        );

    \I__2029\ : InMux
    port map (
            O => \N__10526\,
            I => \N__10463\
        );

    \I__2028\ : InMux
    port map (
            O => \N__10523\,
            I => \N__10456\
        );

    \I__2027\ : InMux
    port map (
            O => \N__10520\,
            I => \N__10456\
        );

    \I__2026\ : InMux
    port map (
            O => \N__10519\,
            I => \N__10456\
        );

    \I__2025\ : InMux
    port map (
            O => \N__10518\,
            I => \N__10453\
        );

    \I__2024\ : InMux
    port map (
            O => \N__10517\,
            I => \N__10450\
        );

    \I__2023\ : InMux
    port map (
            O => \N__10514\,
            I => \N__10443\
        );

    \I__2022\ : InMux
    port map (
            O => \N__10513\,
            I => \N__10443\
        );

    \I__2021\ : InMux
    port map (
            O => \N__10510\,
            I => \N__10443\
        );

    \I__2020\ : InMux
    port map (
            O => \N__10509\,
            I => \N__10430\
        );

    \I__2019\ : InMux
    port map (
            O => \N__10506\,
            I => \N__10430\
        );

    \I__2018\ : InMux
    port map (
            O => \N__10505\,
            I => \N__10430\
        );

    \I__2017\ : InMux
    port map (
            O => \N__10504\,
            I => \N__10430\
        );

    \I__2016\ : InMux
    port map (
            O => \N__10503\,
            I => \N__10430\
        );

    \I__2015\ : InMux
    port map (
            O => \N__10502\,
            I => \N__10430\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__10499\,
            I => \N__10425\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__10494\,
            I => \N__10425\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__10491\,
            I => \N__10417\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__10488\,
            I => \N__10417\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__10483\,
            I => \N__10417\
        );

    \I__2009\ : CascadeMux
    port map (
            O => \N__10482\,
            I => \N__10414\
        );

    \I__2008\ : Span4Mux_v
    port map (
            O => \N__10479\,
            I => \N__10409\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__10474\,
            I => \N__10409\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__10463\,
            I => \N__10406\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__10456\,
            I => \N__10403\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__10453\,
            I => \N__10400\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__10450\,
            I => \N__10393\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__10443\,
            I => \N__10393\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__10430\,
            I => \N__10393\
        );

    \I__2000\ : Span4Mux_v
    port map (
            O => \N__10425\,
            I => \N__10390\
        );

    \I__1999\ : InMux
    port map (
            O => \N__10424\,
            I => \N__10387\
        );

    \I__1998\ : Span4Mux_v
    port map (
            O => \N__10417\,
            I => \N__10384\
        );

    \I__1997\ : InMux
    port map (
            O => \N__10414\,
            I => \N__10381\
        );

    \I__1996\ : Span4Mux_h
    port map (
            O => \N__10409\,
            I => \N__10376\
        );

    \I__1995\ : Span4Mux_h
    port map (
            O => \N__10406\,
            I => \N__10376\
        );

    \I__1994\ : Span4Mux_h
    port map (
            O => \N__10403\,
            I => \N__10369\
        );

    \I__1993\ : Span4Mux_v
    port map (
            O => \N__10400\,
            I => \N__10369\
        );

    \I__1992\ : Span4Mux_h
    port map (
            O => \N__10393\,
            I => \N__10369\
        );

    \I__1991\ : Sp12to4
    port map (
            O => \N__10390\,
            I => \N__10360\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__10387\,
            I => \N__10360\
        );

    \I__1989\ : Sp12to4
    port map (
            O => \N__10384\,
            I => \N__10360\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__10381\,
            I => \N__10360\
        );

    \I__1987\ : Span4Mux_h
    port map (
            O => \N__10376\,
            I => \N__10357\
        );

    \I__1986\ : Span4Mux_h
    port map (
            O => \N__10369\,
            I => \N__10354\
        );

    \I__1985\ : Span12Mux_h
    port map (
            O => \N__10360\,
            I => \N__10351\
        );

    \I__1984\ : Span4Mux_v
    port map (
            O => \N__10357\,
            I => \N__10348\
        );

    \I__1983\ : Span4Mux_v
    port map (
            O => \N__10354\,
            I => \N__10345\
        );

    \I__1982\ : Odrv12
    port map (
            O => \N__10351\,
            I => \P1A1_c\
        );

    \I__1981\ : Odrv4
    port map (
            O => \N__10348\,
            I => \P1A1_c\
        );

    \I__1980\ : Odrv4
    port map (
            O => \N__10345\,
            I => \P1A1_c\
        );

    \I__1979\ : CascadeMux
    port map (
            O => \N__10338\,
            I => \N__10335\
        );

    \I__1978\ : InMux
    port map (
            O => \N__10335\,
            I => \N__10332\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__10332\,
            I => \DUT.uart_inst0.m2_e_0\
        );

    \I__1976\ : InMux
    port map (
            O => \N__10329\,
            I => \N__10326\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__10326\,
            I => \N__10323\
        );

    \I__1974\ : Span4Mux_v
    port map (
            O => \N__10323\,
            I => \N__10320\
        );

    \I__1973\ : Odrv4
    port map (
            O => \N__10320\,
            I => \DUT.uart_inst0.G_19_0_1\
        );

    \I__1972\ : CascadeMux
    port map (
            O => \N__10317\,
            I => \DUT.uart_inst0.G_19_0_a5_0_4_cascade_\
        );

    \I__1971\ : InMux
    port map (
            O => \N__10314\,
            I => \N__10310\
        );

    \I__1970\ : InMux
    port map (
            O => \N__10313\,
            I => \N__10307\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__10310\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_2_0_2\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__10307\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_2_0_2\
        );

    \I__1967\ : InMux
    port map (
            O => \N__10302\,
            I => \N__10299\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__10299\,
            I => \DUT.uart_inst0.G_8_i_a3_1\
        );

    \I__1965\ : InMux
    port map (
            O => \N__10296\,
            I => \N__10293\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__10293\,
            I => \N__10286\
        );

    \I__1963\ : InMux
    port map (
            O => \N__10292\,
            I => \N__10283\
        );

    \I__1962\ : InMux
    port map (
            O => \N__10291\,
            I => \N__10278\
        );

    \I__1961\ : InMux
    port map (
            O => \N__10290\,
            I => \N__10278\
        );

    \I__1960\ : InMux
    port map (
            O => \N__10289\,
            I => \N__10268\
        );

    \I__1959\ : Span4Mux_h
    port map (
            O => \N__10286\,
            I => \N__10261\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__10283\,
            I => \N__10261\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__10278\,
            I => \N__10261\
        );

    \I__1956\ : InMux
    port map (
            O => \N__10277\,
            I => \N__10258\
        );

    \I__1955\ : InMux
    port map (
            O => \N__10276\,
            I => \N__10253\
        );

    \I__1954\ : InMux
    port map (
            O => \N__10275\,
            I => \N__10253\
        );

    \I__1953\ : InMux
    port map (
            O => \N__10274\,
            I => \N__10246\
        );

    \I__1952\ : InMux
    port map (
            O => \N__10273\,
            I => \N__10246\
        );

    \I__1951\ : InMux
    port map (
            O => \N__10272\,
            I => \N__10246\
        );

    \I__1950\ : InMux
    port map (
            O => \N__10271\,
            I => \N__10243\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__10268\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_4\
        );

    \I__1948\ : Odrv4
    port map (
            O => \N__10261\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_4\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__10258\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_4\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__10253\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_4\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__10246\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_4\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__10243\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_4\
        );

    \I__1943\ : InMux
    port map (
            O => \N__10230\,
            I => \N__10225\
        );

    \I__1942\ : InMux
    port map (
            O => \N__10229\,
            I => \N__10222\
        );

    \I__1941\ : InMux
    port map (
            O => \N__10228\,
            I => \N__10211\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__10225\,
            I => \N__10206\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__10222\,
            I => \N__10206\
        );

    \I__1938\ : InMux
    port map (
            O => \N__10221\,
            I => \N__10201\
        );

    \I__1937\ : InMux
    port map (
            O => \N__10220\,
            I => \N__10201\
        );

    \I__1936\ : InMux
    port map (
            O => \N__10219\,
            I => \N__10198\
        );

    \I__1935\ : InMux
    port map (
            O => \N__10218\,
            I => \N__10193\
        );

    \I__1934\ : InMux
    port map (
            O => \N__10217\,
            I => \N__10193\
        );

    \I__1933\ : InMux
    port map (
            O => \N__10216\,
            I => \N__10190\
        );

    \I__1932\ : InMux
    port map (
            O => \N__10215\,
            I => \N__10185\
        );

    \I__1931\ : InMux
    port map (
            O => \N__10214\,
            I => \N__10185\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__10211\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_5\
        );

    \I__1929\ : Odrv4
    port map (
            O => \N__10206\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_5\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__10201\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_5\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__10198\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_5\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__10193\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_5\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__10190\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_5\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__10185\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_5\
        );

    \I__1923\ : InMux
    port map (
            O => \N__10170\,
            I => \N__10165\
        );

    \I__1922\ : CascadeMux
    port map (
            O => \N__10169\,
            I => \N__10160\
        );

    \I__1921\ : CascadeMux
    port map (
            O => \N__10168\,
            I => \N__10154\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__10165\,
            I => \N__10148\
        );

    \I__1919\ : InMux
    port map (
            O => \N__10164\,
            I => \N__10143\
        );

    \I__1918\ : InMux
    port map (
            O => \N__10163\,
            I => \N__10143\
        );

    \I__1917\ : InMux
    port map (
            O => \N__10160\,
            I => \N__10139\
        );

    \I__1916\ : InMux
    port map (
            O => \N__10159\,
            I => \N__10136\
        );

    \I__1915\ : InMux
    port map (
            O => \N__10158\,
            I => \N__10129\
        );

    \I__1914\ : InMux
    port map (
            O => \N__10157\,
            I => \N__10129\
        );

    \I__1913\ : InMux
    port map (
            O => \N__10154\,
            I => \N__10129\
        );

    \I__1912\ : InMux
    port map (
            O => \N__10153\,
            I => \N__10122\
        );

    \I__1911\ : InMux
    port map (
            O => \N__10152\,
            I => \N__10122\
        );

    \I__1910\ : InMux
    port map (
            O => \N__10151\,
            I => \N__10122\
        );

    \I__1909\ : Span4Mux_h
    port map (
            O => \N__10148\,
            I => \N__10117\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__10143\,
            I => \N__10117\
        );

    \I__1907\ : InMux
    port map (
            O => \N__10142\,
            I => \N__10114\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__10139\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_3\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__10136\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_3\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__10129\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_3\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__10122\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_3\
        );

    \I__1902\ : Odrv4
    port map (
            O => \N__10117\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_3\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__10114\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_3\
        );

    \I__1900\ : InMux
    port map (
            O => \N__10101\,
            I => \N__10094\
        );

    \I__1899\ : CascadeMux
    port map (
            O => \N__10100\,
            I => \N__10090\
        );

    \I__1898\ : InMux
    port map (
            O => \N__10099\,
            I => \N__10087\
        );

    \I__1897\ : InMux
    port map (
            O => \N__10098\,
            I => \N__10082\
        );

    \I__1896\ : InMux
    port map (
            O => \N__10097\,
            I => \N__10082\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__10094\,
            I => \N__10077\
        );

    \I__1894\ : InMux
    port map (
            O => \N__10093\,
            I => \N__10072\
        );

    \I__1893\ : InMux
    port map (
            O => \N__10090\,
            I => \N__10072\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__10087\,
            I => \N__10066\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__10082\,
            I => \N__10066\
        );

    \I__1890\ : InMux
    port map (
            O => \N__10081\,
            I => \N__10061\
        );

    \I__1889\ : InMux
    port map (
            O => \N__10080\,
            I => \N__10058\
        );

    \I__1888\ : Span4Mux_v
    port map (
            O => \N__10077\,
            I => \N__10052\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__10072\,
            I => \N__10052\
        );

    \I__1886\ : InMux
    port map (
            O => \N__10071\,
            I => \N__10046\
        );

    \I__1885\ : Span4Mux_v
    port map (
            O => \N__10066\,
            I => \N__10043\
        );

    \I__1884\ : InMux
    port map (
            O => \N__10065\,
            I => \N__10038\
        );

    \I__1883\ : InMux
    port map (
            O => \N__10064\,
            I => \N__10038\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__10061\,
            I => \N__10033\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__10058\,
            I => \N__10033\
        );

    \I__1880\ : InMux
    port map (
            O => \N__10057\,
            I => \N__10030\
        );

    \I__1879\ : Span4Mux_h
    port map (
            O => \N__10052\,
            I => \N__10027\
        );

    \I__1878\ : InMux
    port map (
            O => \N__10051\,
            I => \N__10022\
        );

    \I__1877\ : InMux
    port map (
            O => \N__10050\,
            I => \N__10022\
        );

    \I__1876\ : InMux
    port map (
            O => \N__10049\,
            I => \N__10019\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__10046\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__1874\ : Odrv4
    port map (
            O => \N__10043\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__10038\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__1872\ : Odrv4
    port map (
            O => \N__10033\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__10030\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__1870\ : Odrv4
    port map (
            O => \N__10027\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__10022\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__10019\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__1867\ : CascadeMux
    port map (
            O => \N__10002\,
            I => \N__9998\
        );

    \I__1866\ : InMux
    port map (
            O => \N__10001\,
            I => \N__9992\
        );

    \I__1865\ : InMux
    port map (
            O => \N__9998\,
            I => \N__9989\
        );

    \I__1864\ : InMux
    port map (
            O => \N__9997\,
            I => \N__9986\
        );

    \I__1863\ : CascadeMux
    port map (
            O => \N__9996\,
            I => \N__9978\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__9995\,
            I => \N__9974\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__9992\,
            I => \N__9969\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__9989\,
            I => \N__9969\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__9986\,
            I => \N__9966\
        );

    \I__1858\ : InMux
    port map (
            O => \N__9985\,
            I => \N__9963\
        );

    \I__1857\ : InMux
    port map (
            O => \N__9984\,
            I => \N__9958\
        );

    \I__1856\ : InMux
    port map (
            O => \N__9983\,
            I => \N__9958\
        );

    \I__1855\ : InMux
    port map (
            O => \N__9982\,
            I => \N__9955\
        );

    \I__1854\ : InMux
    port map (
            O => \N__9981\,
            I => \N__9948\
        );

    \I__1853\ : InMux
    port map (
            O => \N__9978\,
            I => \N__9948\
        );

    \I__1852\ : InMux
    port map (
            O => \N__9977\,
            I => \N__9948\
        );

    \I__1851\ : InMux
    port map (
            O => \N__9974\,
            I => \N__9945\
        );

    \I__1850\ : Span4Mux_v
    port map (
            O => \N__9969\,
            I => \N__9940\
        );

    \I__1849\ : Span4Mux_v
    port map (
            O => \N__9966\,
            I => \N__9940\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__9963\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_2\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__9958\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_2\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__9955\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_2\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__9948\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_2\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__9945\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_2\
        );

    \I__1843\ : Odrv4
    port map (
            O => \N__9940\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_2\
        );

    \I__1842\ : InMux
    port map (
            O => \N__9927\,
            I => \N__9922\
        );

    \I__1841\ : InMux
    port map (
            O => \N__9926\,
            I => \N__9914\
        );

    \I__1840\ : InMux
    port map (
            O => \N__9925\,
            I => \N__9914\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__9922\,
            I => \N__9910\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__9921\,
            I => \N__9904\
        );

    \I__1837\ : CascadeMux
    port map (
            O => \N__9920\,
            I => \N__9900\
        );

    \I__1836\ : InMux
    port map (
            O => \N__9919\,
            I => \N__9896\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__9914\,
            I => \N__9893\
        );

    \I__1834\ : InMux
    port map (
            O => \N__9913\,
            I => \N__9890\
        );

    \I__1833\ : Span4Mux_v
    port map (
            O => \N__9910\,
            I => \N__9887\
        );

    \I__1832\ : InMux
    port map (
            O => \N__9909\,
            I => \N__9884\
        );

    \I__1831\ : InMux
    port map (
            O => \N__9908\,
            I => \N__9881\
        );

    \I__1830\ : InMux
    port map (
            O => \N__9907\,
            I => \N__9878\
        );

    \I__1829\ : InMux
    port map (
            O => \N__9904\,
            I => \N__9873\
        );

    \I__1828\ : InMux
    port map (
            O => \N__9903\,
            I => \N__9873\
        );

    \I__1827\ : InMux
    port map (
            O => \N__9900\,
            I => \N__9868\
        );

    \I__1826\ : InMux
    port map (
            O => \N__9899\,
            I => \N__9868\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__9896\,
            I => \N__9861\
        );

    \I__1824\ : Span4Mux_h
    port map (
            O => \N__9893\,
            I => \N__9861\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__9890\,
            I => \N__9861\
        );

    \I__1822\ : Odrv4
    port map (
            O => \N__9887\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_1\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__9884\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_1\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__9881\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_1\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__9878\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_1\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__9873\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_1\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__9868\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_1\
        );

    \I__1816\ : Odrv4
    port map (
            O => \N__9861\,
            I => \DUT_uart_inst0_rx_countdown_3_s1_1\
        );

    \I__1815\ : InMux
    port map (
            O => \N__9846\,
            I => \N__9843\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__9843\,
            I => \DUT.uart_inst0.G_19_0_a5_4\
        );

    \I__1813\ : InMux
    port map (
            O => \N__9840\,
            I => \N__9833\
        );

    \I__1812\ : InMux
    port map (
            O => \N__9839\,
            I => \N__9833\
        );

    \I__1811\ : InMux
    port map (
            O => \N__9838\,
            I => \N__9830\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__9833\,
            I => \N__9827\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__9830\,
            I => \N__9822\
        );

    \I__1808\ : Span4Mux_h
    port map (
            O => \N__9827\,
            I => \N__9822\
        );

    \I__1807\ : Odrv4
    port map (
            O => \N__9822\,
            I => \DUT.uart_inst0.N_44\
        );

    \I__1806\ : InMux
    port map (
            O => \N__9819\,
            I => \N__9816\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__9816\,
            I => \N__9813\
        );

    \I__1804\ : Span4Mux_h
    port map (
            O => \N__9813\,
            I => \N__9810\
        );

    \I__1803\ : Odrv4
    port map (
            O => \N__9810\,
            I => \DUT.uart_inst0.g1_i_a4_1_5\
        );

    \I__1802\ : CascadeMux
    port map (
            O => \N__9807\,
            I => \N__9804\
        );

    \I__1801\ : InMux
    port map (
            O => \N__9804\,
            I => \N__9801\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__9801\,
            I => \DUT.uart_inst0.g1_i_a4_1_3\
        );

    \I__1799\ : CascadeMux
    port map (
            O => \N__9798\,
            I => \DUT.uart_inst0.N_78_cascade_\
        );

    \I__1798\ : CascadeMux
    port map (
            O => \N__9795\,
            I => \DUT.uart_inst0.N_10_mux_cascade_\
        );

    \I__1797\ : InMux
    port map (
            O => \N__9792\,
            I => \N__9789\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__9789\,
            I => \DUT.uart_inst0.P6_mux\
        );

    \I__1795\ : CascadeMux
    port map (
            O => \N__9786\,
            I => \DUT.uart_inst0.G_19_0_a5_0_2_cascade_\
        );

    \I__1794\ : CEMux
    port map (
            O => \N__9783\,
            I => \N__9780\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__9780\,
            I => \N__9777\
        );

    \I__1792\ : Span4Mux_v
    port map (
            O => \N__9777\,
            I => \N__9774\
        );

    \I__1791\ : Odrv4
    port map (
            O => \N__9774\,
            I => \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa\
        );

    \I__1790\ : InMux
    port map (
            O => \N__9771\,
            I => \N__9768\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__9768\,
            I => \DUT.uart_inst0.m6_2\
        );

    \I__1788\ : CascadeMux
    port map (
            O => \N__9765\,
            I => \N__9761\
        );

    \I__1787\ : InMux
    port map (
            O => \N__9764\,
            I => \N__9758\
        );

    \I__1786\ : InMux
    port map (
            O => \N__9761\,
            I => \N__9755\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__9758\,
            I => \N__9749\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__9755\,
            I => \N__9749\
        );

    \I__1783\ : InMux
    port map (
            O => \N__9754\,
            I => \N__9746\
        );

    \I__1782\ : Span4Mux_v
    port map (
            O => \N__9749\,
            I => \N__9743\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__9746\,
            I => \N__9740\
        );

    \I__1780\ : Odrv4
    port map (
            O => \N__9743\,
            I => \G_114\
        );

    \I__1779\ : Odrv12
    port map (
            O => \N__9740\,
            I => \G_114\
        );

    \I__1778\ : InMux
    port map (
            O => \N__9735\,
            I => \N__9732\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__9732\,
            I => \N__9727\
        );

    \I__1776\ : InMux
    port map (
            O => \N__9731\,
            I => \N__9724\
        );

    \I__1775\ : InMux
    port map (
            O => \N__9730\,
            I => \N__9721\
        );

    \I__1774\ : Odrv4
    port map (
            O => \N__9727\,
            I => \G_113\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__9724\,
            I => \G_113\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__9721\,
            I => \G_113\
        );

    \I__1771\ : CascadeMux
    port map (
            O => \N__9714\,
            I => \fifo_inst.ftdi_input_inst.un1_rWrStateZ0Z_1_cascade_\
        );

    \I__1770\ : CascadeMux
    port map (
            O => \N__9711\,
            I => \N__9708\
        );

    \I__1769\ : InMux
    port map (
            O => \N__9708\,
            I => \N__9705\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__9705\,
            I => \N__9701\
        );

    \I__1767\ : InMux
    port map (
            O => \N__9704\,
            I => \N__9698\
        );

    \I__1766\ : Odrv4
    port map (
            O => \N__9701\,
            I => \G_118\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__9698\,
            I => \G_118\
        );

    \I__1764\ : CascadeMux
    port map (
            O => \N__9693\,
            I => \G_118_cascade_\
        );

    \I__1763\ : InMux
    port map (
            O => \N__9690\,
            I => \N__9687\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__9687\,
            I => \G_119\
        );

    \I__1761\ : CascadeMux
    port map (
            O => \N__9684\,
            I => \N__9681\
        );

    \I__1760\ : InMux
    port map (
            O => \N__9681\,
            I => \N__9678\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__9678\,
            I => \N__9673\
        );

    \I__1758\ : InMux
    port map (
            O => \N__9677\,
            I => \N__9670\
        );

    \I__1757\ : InMux
    port map (
            O => \N__9676\,
            I => \N__9667\
        );

    \I__1756\ : Odrv12
    port map (
            O => \N__9673\,
            I => \G_116\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__9670\,
            I => \G_116\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__9667\,
            I => \G_116\
        );

    \I__1753\ : InMux
    port map (
            O => \N__9660\,
            I => \N__9654\
        );

    \I__1752\ : InMux
    port map (
            O => \N__9659\,
            I => \N__9654\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__9654\,
            I => \fifo_inst.ftdi_input_inst.un1_rWrStateZ0Z_1\
        );

    \I__1750\ : CascadeMux
    port map (
            O => \N__9651\,
            I => \G_116_cascade_\
        );

    \I__1749\ : CascadeMux
    port map (
            O => \N__9648\,
            I => \N__9645\
        );

    \I__1748\ : InMux
    port map (
            O => \N__9645\,
            I => \N__9642\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__9642\,
            I => \N__9637\
        );

    \I__1746\ : InMux
    port map (
            O => \N__9641\,
            I => \N__9634\
        );

    \I__1745\ : InMux
    port map (
            O => \N__9640\,
            I => \N__9631\
        );

    \I__1744\ : Odrv12
    port map (
            O => \N__9637\,
            I => \G_117\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__9634\,
            I => \G_117\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__9631\,
            I => \G_117\
        );

    \I__1741\ : CascadeMux
    port map (
            O => \N__9624\,
            I => \N__9621\
        );

    \I__1740\ : InMux
    port map (
            O => \N__9621\,
            I => \N__9618\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__9618\,
            I => \N__9615\
        );

    \I__1738\ : Odrv4
    port map (
            O => \N__9615\,
            I => \DUT.rFifoDataror_1\
        );

    \I__1737\ : CascadeMux
    port map (
            O => \N__9612\,
            I => \DUT.rFifoDataror_1_cascade_\
        );

    \I__1736\ : InMux
    port map (
            O => \N__9609\,
            I => \N__9606\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__9606\,
            I => \N__9602\
        );

    \I__1734\ : InMux
    port map (
            O => \N__9605\,
            I => \N__9599\
        );

    \I__1733\ : Odrv4
    port map (
            O => \N__9602\,
            I => \DUT.rFifoDataror_0_0\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__9599\,
            I => \DUT.rFifoDataror_0_0\
        );

    \I__1731\ : InMux
    port map (
            O => \N__9594\,
            I => \N__9573\
        );

    \I__1730\ : InMux
    port map (
            O => \N__9593\,
            I => \N__9573\
        );

    \I__1729\ : InMux
    port map (
            O => \N__9592\,
            I => \N__9573\
        );

    \I__1728\ : InMux
    port map (
            O => \N__9591\,
            I => \N__9573\
        );

    \I__1727\ : InMux
    port map (
            O => \N__9590\,
            I => \N__9573\
        );

    \I__1726\ : InMux
    port map (
            O => \N__9589\,
            I => \N__9573\
        );

    \I__1725\ : InMux
    port map (
            O => \N__9588\,
            I => \N__9573\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__9573\,
            I => \DUT.rFifoDataror_0\
        );

    \I__1723\ : InMux
    port map (
            O => \N__9570\,
            I => \N__9566\
        );

    \I__1722\ : SRMux
    port map (
            O => \N__9569\,
            I => \N__9563\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__9566\,
            I => \N__9560\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__9563\,
            I => \N__9557\
        );

    \I__1719\ : Span4Mux_s3_v
    port map (
            O => \N__9560\,
            I => \N__9551\
        );

    \I__1718\ : Span4Mux_h
    port map (
            O => \N__9557\,
            I => \N__9551\
        );

    \I__1717\ : InMux
    port map (
            O => \N__9556\,
            I => \N__9548\
        );

    \I__1716\ : Odrv4
    port map (
            O => \N__9551\,
            I => \G_115\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__9548\,
            I => \G_115\
        );

    \I__1714\ : InMux
    port map (
            O => \N__9543\,
            I => \N__9540\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__9540\,
            I => \DUT.rFifoDatarx_5\
        );

    \I__1712\ : InMux
    port map (
            O => \N__9537\,
            I => \N__9534\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__9534\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_5\
        );

    \I__1710\ : InMux
    port map (
            O => \N__9531\,
            I => \N__9528\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__9528\,
            I => \N__9525\
        );

    \I__1708\ : Odrv12
    port map (
            O => \N__9525\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_6\
        );

    \I__1707\ : CascadeMux
    port map (
            O => \N__9522\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_\
        );

    \I__1706\ : InMux
    port map (
            O => \N__9519\,
            I => \N__9516\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__9516\,
            I => \DUT.rFifoDatarx_6\
        );

    \I__1704\ : InMux
    port map (
            O => \N__9513\,
            I => \N__9508\
        );

    \I__1703\ : InMux
    port map (
            O => \N__9512\,
            I => \N__9505\
        );

    \I__1702\ : CascadeMux
    port map (
            O => \N__9511\,
            I => \N__9502\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__9508\,
            I => \N__9497\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__9505\,
            I => \N__9497\
        );

    \I__1699\ : InMux
    port map (
            O => \N__9502\,
            I => \N__9492\
        );

    \I__1698\ : Span4Mux_h
    port map (
            O => \N__9497\,
            I => \N__9489\
        );

    \I__1697\ : InMux
    port map (
            O => \N__9496\,
            I => \N__9484\
        );

    \I__1696\ : InMux
    port map (
            O => \N__9495\,
            I => \N__9484\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__9492\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_1\
        );

    \I__1694\ : Odrv4
    port map (
            O => \N__9489\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_1\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__9484\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_1\
        );

    \I__1692\ : InMux
    port map (
            O => \N__9477\,
            I => \N__9473\
        );

    \I__1691\ : InMux
    port map (
            O => \N__9476\,
            I => \N__9470\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__9473\,
            I => \N__9464\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__9470\,
            I => \N__9464\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__9469\,
            I => \N__9461\
        );

    \I__1687\ : Span4Mux_h
    port map (
            O => \N__9464\,
            I => \N__9458\
        );

    \I__1686\ : InMux
    port map (
            O => \N__9461\,
            I => \N__9452\
        );

    \I__1685\ : Span4Mux_v
    port map (
            O => \N__9458\,
            I => \N__9449\
        );

    \I__1684\ : InMux
    port map (
            O => \N__9457\,
            I => \N__9442\
        );

    \I__1683\ : InMux
    port map (
            O => \N__9456\,
            I => \N__9442\
        );

    \I__1682\ : InMux
    port map (
            O => \N__9455\,
            I => \N__9442\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__9452\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_0\
        );

    \I__1680\ : Odrv4
    port map (
            O => \N__9449\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_0\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__9442\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_0\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__9435\,
            I => \N__9431\
        );

    \I__1677\ : CascadeMux
    port map (
            O => \N__9434\,
            I => \N__9426\
        );

    \I__1676\ : InMux
    port map (
            O => \N__9431\,
            I => \N__9422\
        );

    \I__1675\ : InMux
    port map (
            O => \N__9430\,
            I => \N__9417\
        );

    \I__1674\ : InMux
    port map (
            O => \N__9429\,
            I => \N__9417\
        );

    \I__1673\ : InMux
    port map (
            O => \N__9426\,
            I => \N__9413\
        );

    \I__1672\ : InMux
    port map (
            O => \N__9425\,
            I => \N__9409\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__9422\,
            I => \N__9403\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__9417\,
            I => \N__9403\
        );

    \I__1669\ : InMux
    port map (
            O => \N__9416\,
            I => \N__9400\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__9413\,
            I => \N__9394\
        );

    \I__1667\ : CascadeMux
    port map (
            O => \N__9412\,
            I => \N__9391\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__9409\,
            I => \N__9388\
        );

    \I__1665\ : InMux
    port map (
            O => \N__9408\,
            I => \N__9385\
        );

    \I__1664\ : Span4Mux_h
    port map (
            O => \N__9403\,
            I => \N__9382\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__9400\,
            I => \N__9379\
        );

    \I__1662\ : InMux
    port map (
            O => \N__9399\,
            I => \N__9374\
        );

    \I__1661\ : InMux
    port map (
            O => \N__9398\,
            I => \N__9374\
        );

    \I__1660\ : InMux
    port map (
            O => \N__9397\,
            I => \N__9369\
        );

    \I__1659\ : Span4Mux_v
    port map (
            O => \N__9394\,
            I => \N__9366\
        );

    \I__1658\ : InMux
    port map (
            O => \N__9391\,
            I => \N__9363\
        );

    \I__1657\ : Span4Mux_h
    port map (
            O => \N__9388\,
            I => \N__9360\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__9385\,
            I => \N__9351\
        );

    \I__1655\ : Span4Mux_v
    port map (
            O => \N__9382\,
            I => \N__9351\
        );

    \I__1654\ : Span4Mux_s2_v
    port map (
            O => \N__9379\,
            I => \N__9351\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__9374\,
            I => \N__9351\
        );

    \I__1652\ : InMux
    port map (
            O => \N__9373\,
            I => \N__9346\
        );

    \I__1651\ : InMux
    port map (
            O => \N__9372\,
            I => \N__9346\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__9369\,
            I => \DUT.rTransmitZ0\
        );

    \I__1649\ : Odrv4
    port map (
            O => \N__9366\,
            I => \DUT.rTransmitZ0\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__9363\,
            I => \DUT.rTransmitZ0\
        );

    \I__1647\ : Odrv4
    port map (
            O => \N__9360\,
            I => \DUT.rTransmitZ0\
        );

    \I__1646\ : Odrv4
    port map (
            O => \N__9351\,
            I => \DUT.rTransmitZ0\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__9346\,
            I => \DUT.rTransmitZ0\
        );

    \I__1644\ : InMux
    port map (
            O => \N__9333\,
            I => \N__9329\
        );

    \I__1643\ : InMux
    port map (
            O => \N__9332\,
            I => \N__9326\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__9329\,
            I => \N__9320\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__9326\,
            I => \N__9320\
        );

    \I__1640\ : InMux
    port map (
            O => \N__9325\,
            I => \N__9314\
        );

    \I__1639\ : Span4Mux_h
    port map (
            O => \N__9320\,
            I => \N__9311\
        );

    \I__1638\ : InMux
    port map (
            O => \N__9319\,
            I => \N__9304\
        );

    \I__1637\ : InMux
    port map (
            O => \N__9318\,
            I => \N__9304\
        );

    \I__1636\ : InMux
    port map (
            O => \N__9317\,
            I => \N__9304\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__9314\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_2\
        );

    \I__1634\ : Odrv4
    port map (
            O => \N__9311\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_2\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__9304\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_2\
        );

    \I__1632\ : CascadeMux
    port map (
            O => \N__9297\,
            I => \DUT.fifo_tx_inst.rReadPtr11_cascade_\
        );

    \I__1631\ : CascadeMux
    port map (
            O => \N__9294\,
            I => \DUT.fifo_tx_inst.un1_i11_2_i_cascade_\
        );

    \I__1630\ : InMux
    port map (
            O => \N__9291\,
            I => \N__9285\
        );

    \I__1629\ : InMux
    port map (
            O => \N__9290\,
            I => \N__9285\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__9285\,
            I => \DUT.fifo_tx_inst.rReadPtr11\
        );

    \I__1627\ : InMux
    port map (
            O => \N__9282\,
            I => \N__9279\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__9279\,
            I => \DUT.fifo_tx_inst.un1_i11_2_i\
        );

    \I__1625\ : CascadeMux
    port map (
            O => \N__9276\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_\
        );

    \I__1624\ : InMux
    port map (
            O => \N__9273\,
            I => \N__9270\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__9270\,
            I => \N__9267\
        );

    \I__1622\ : Odrv4
    port map (
            O => \N__9267\,
            I => \DUT.rFifoDatarx_0\
        );

    \I__1621\ : InMux
    port map (
            O => \N__9264\,
            I => \N__9261\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__9261\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_0\
        );

    \I__1619\ : InMux
    port map (
            O => \N__9258\,
            I => \N__9255\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__9255\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_1\
        );

    \I__1617\ : CascadeMux
    port map (
            O => \N__9252\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1_cascade_\
        );

    \I__1616\ : InMux
    port map (
            O => \N__9249\,
            I => \N__9246\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__9246\,
            I => \DUT.rFifoDatarx_1\
        );

    \I__1614\ : CascadeMux
    port map (
            O => \N__9243\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_\
        );

    \I__1613\ : InMux
    port map (
            O => \N__9240\,
            I => \N__9237\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__9237\,
            I => \DUT.rFifoDatarx_4\
        );

    \I__1611\ : InMux
    port map (
            O => \N__9234\,
            I => \N__9231\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__9231\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_4\
        );

    \I__1609\ : CascadeMux
    port map (
            O => \N__9228\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_\
        );

    \I__1608\ : InMux
    port map (
            O => \N__9225\,
            I => \N__9222\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__9222\,
            I => \N__9219\
        );

    \I__1606\ : Odrv4
    port map (
            O => \N__9219\,
            I => \DUT.uart_inst0.N_19\
        );

    \I__1605\ : InMux
    port map (
            O => \N__9216\,
            I => \N__9213\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__9213\,
            I => \DUT.uart_inst0.G_8_i_a3_0_0\
        );

    \I__1603\ : CascadeMux
    port map (
            O => \N__9210\,
            I => \N__9207\
        );

    \I__1602\ : InMux
    port map (
            O => \N__9207\,
            I => \N__9204\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__9204\,
            I => \N__9201\
        );

    \I__1600\ : Span4Mux_h
    port map (
            O => \N__9201\,
            I => \N__9198\
        );

    \I__1599\ : Odrv4
    port map (
            O => \N__9198\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_1_1_2\
        );

    \I__1598\ : CascadeMux
    port map (
            O => \N__9195\,
            I => \N__9174\
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__9194\,
            I => \N__9171\
        );

    \I__1596\ : CascadeMux
    port map (
            O => \N__9193\,
            I => \N__9168\
        );

    \I__1595\ : CascadeMux
    port map (
            O => \N__9192\,
            I => \N__9165\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__9191\,
            I => \N__9162\
        );

    \I__1593\ : CascadeMux
    port map (
            O => \N__9190\,
            I => \N__9159\
        );

    \I__1592\ : CascadeMux
    port map (
            O => \N__9189\,
            I => \N__9156\
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__9188\,
            I => \N__9153\
        );

    \I__1590\ : CascadeMux
    port map (
            O => \N__9187\,
            I => \N__9150\
        );

    \I__1589\ : CascadeMux
    port map (
            O => \N__9186\,
            I => \N__9147\
        );

    \I__1588\ : CascadeMux
    port map (
            O => \N__9185\,
            I => \N__9144\
        );

    \I__1587\ : CascadeMux
    port map (
            O => \N__9184\,
            I => \N__9141\
        );

    \I__1586\ : CascadeMux
    port map (
            O => \N__9183\,
            I => \N__9138\
        );

    \I__1585\ : CascadeMux
    port map (
            O => \N__9182\,
            I => \N__9135\
        );

    \I__1584\ : CascadeMux
    port map (
            O => \N__9181\,
            I => \N__9132\
        );

    \I__1583\ : CascadeMux
    port map (
            O => \N__9180\,
            I => \N__9129\
        );

    \I__1582\ : SRMux
    port map (
            O => \N__9179\,
            I => \N__9121\
        );

    \I__1581\ : InMux
    port map (
            O => \N__9178\,
            I => \N__9116\
        );

    \I__1580\ : InMux
    port map (
            O => \N__9177\,
            I => \N__9116\
        );

    \I__1579\ : InMux
    port map (
            O => \N__9174\,
            I => \N__9110\
        );

    \I__1578\ : InMux
    port map (
            O => \N__9171\,
            I => \N__9101\
        );

    \I__1577\ : InMux
    port map (
            O => \N__9168\,
            I => \N__9101\
        );

    \I__1576\ : InMux
    port map (
            O => \N__9165\,
            I => \N__9101\
        );

    \I__1575\ : InMux
    port map (
            O => \N__9162\,
            I => \N__9101\
        );

    \I__1574\ : InMux
    port map (
            O => \N__9159\,
            I => \N__9094\
        );

    \I__1573\ : InMux
    port map (
            O => \N__9156\,
            I => \N__9094\
        );

    \I__1572\ : InMux
    port map (
            O => \N__9153\,
            I => \N__9094\
        );

    \I__1571\ : InMux
    port map (
            O => \N__9150\,
            I => \N__9085\
        );

    \I__1570\ : InMux
    port map (
            O => \N__9147\,
            I => \N__9085\
        );

    \I__1569\ : InMux
    port map (
            O => \N__9144\,
            I => \N__9085\
        );

    \I__1568\ : InMux
    port map (
            O => \N__9141\,
            I => \N__9085\
        );

    \I__1567\ : InMux
    port map (
            O => \N__9138\,
            I => \N__9076\
        );

    \I__1566\ : InMux
    port map (
            O => \N__9135\,
            I => \N__9076\
        );

    \I__1565\ : InMux
    port map (
            O => \N__9132\,
            I => \N__9076\
        );

    \I__1564\ : InMux
    port map (
            O => \N__9129\,
            I => \N__9076\
        );

    \I__1563\ : CascadeMux
    port map (
            O => \N__9128\,
            I => \N__9073\
        );

    \I__1562\ : CascadeMux
    port map (
            O => \N__9127\,
            I => \N__9070\
        );

    \I__1561\ : CascadeMux
    port map (
            O => \N__9126\,
            I => \N__9067\
        );

    \I__1560\ : CascadeMux
    port map (
            O => \N__9125\,
            I => \N__9064\
        );

    \I__1559\ : CascadeMux
    port map (
            O => \N__9124\,
            I => \N__9061\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__9121\,
            I => \N__9051\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__9116\,
            I => \N__9048\
        );

    \I__1556\ : InMux
    port map (
            O => \N__9115\,
            I => \N__9041\
        );

    \I__1555\ : InMux
    port map (
            O => \N__9114\,
            I => \N__9041\
        );

    \I__1554\ : InMux
    port map (
            O => \N__9113\,
            I => \N__9041\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__9110\,
            I => \N__9034\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__9101\,
            I => \N__9034\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__9094\,
            I => \N__9034\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__9085\,
            I => \N__9029\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__9076\,
            I => \N__9029\
        );

    \I__1548\ : InMux
    port map (
            O => \N__9073\,
            I => \N__9024\
        );

    \I__1547\ : InMux
    port map (
            O => \N__9070\,
            I => \N__9024\
        );

    \I__1546\ : InMux
    port map (
            O => \N__9067\,
            I => \N__9017\
        );

    \I__1545\ : InMux
    port map (
            O => \N__9064\,
            I => \N__9017\
        );

    \I__1544\ : InMux
    port map (
            O => \N__9061\,
            I => \N__9017\
        );

    \I__1543\ : CascadeMux
    port map (
            O => \N__9060\,
            I => \N__9014\
        );

    \I__1542\ : CascadeMux
    port map (
            O => \N__9059\,
            I => \N__9011\
        );

    \I__1541\ : CascadeMux
    port map (
            O => \N__9058\,
            I => \N__9008\
        );

    \I__1540\ : CascadeMux
    port map (
            O => \N__9057\,
            I => \N__9005\
        );

    \I__1539\ : CascadeMux
    port map (
            O => \N__9056\,
            I => \N__9002\
        );

    \I__1538\ : CascadeMux
    port map (
            O => \N__9055\,
            I => \N__8999\
        );

    \I__1537\ : CascadeMux
    port map (
            O => \N__9054\,
            I => \N__8996\
        );

    \I__1536\ : Span4Mux_v
    port map (
            O => \N__9051\,
            I => \N__8993\
        );

    \I__1535\ : Span4Mux_h
    port map (
            O => \N__9048\,
            I => \N__8990\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__9041\,
            I => \N__8987\
        );

    \I__1533\ : Span4Mux_v
    port map (
            O => \N__9034\,
            I => \N__8978\
        );

    \I__1532\ : Span4Mux_v
    port map (
            O => \N__9029\,
            I => \N__8978\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__9024\,
            I => \N__8978\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__9017\,
            I => \N__8978\
        );

    \I__1529\ : InMux
    port map (
            O => \N__9014\,
            I => \N__8971\
        );

    \I__1528\ : InMux
    port map (
            O => \N__9011\,
            I => \N__8971\
        );

    \I__1527\ : InMux
    port map (
            O => \N__9008\,
            I => \N__8971\
        );

    \I__1526\ : InMux
    port map (
            O => \N__9005\,
            I => \N__8962\
        );

    \I__1525\ : InMux
    port map (
            O => \N__9002\,
            I => \N__8962\
        );

    \I__1524\ : InMux
    port map (
            O => \N__8999\,
            I => \N__8962\
        );

    \I__1523\ : InMux
    port map (
            O => \N__8996\,
            I => \N__8962\
        );

    \I__1522\ : Span4Mux_h
    port map (
            O => \N__8993\,
            I => \N__8955\
        );

    \I__1521\ : Span4Mux_v
    port map (
            O => \N__8990\,
            I => \N__8955\
        );

    \I__1520\ : Span4Mux_v
    port map (
            O => \N__8987\,
            I => \N__8955\
        );

    \I__1519\ : Span4Mux_v
    port map (
            O => \N__8978\,
            I => \N__8948\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__8971\,
            I => \N__8948\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__8962\,
            I => \N__8948\
        );

    \I__1516\ : Odrv4
    port map (
            O => \N__8955\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1515\ : Odrv4
    port map (
            O => \N__8948\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1514\ : CascadeMux
    port map (
            O => \N__8943\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_\
        );

    \I__1513\ : InMux
    port map (
            O => \N__8940\,
            I => \N__8937\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__8937\,
            I => \DUT.rFifoDatarx_7\
        );

    \I__1511\ : InMux
    port map (
            O => \N__8934\,
            I => \N__8931\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__8931\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_7\
        );

    \I__1509\ : InMux
    port map (
            O => \N__8928\,
            I => \N__8925\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__8925\,
            I => \DUT.uart_inst0.m6_1\
        );

    \I__1507\ : InMux
    port map (
            O => \N__8922\,
            I => \N__8916\
        );

    \I__1506\ : InMux
    port map (
            O => \N__8921\,
            I => \N__8916\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__8916\,
            I => \DUT.uart_inst0.N_7\
        );

    \I__1504\ : InMux
    port map (
            O => \N__8913\,
            I => \N__8910\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__8910\,
            I => \DUT.uart_inst0.recv_state_srsts_1_5\
        );

    \I__1502\ : InMux
    port map (
            O => \N__8907\,
            I => \N__8902\
        );

    \I__1501\ : InMux
    port map (
            O => \N__8906\,
            I => \N__8897\
        );

    \I__1500\ : InMux
    port map (
            O => \N__8905\,
            I => \N__8897\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__8902\,
            I => \N__8894\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__8897\,
            I => \N__8891\
        );

    \I__1497\ : Span4Mux_v
    port map (
            O => \N__8894\,
            I => \N__8888\
        );

    \I__1496\ : Odrv4
    port map (
            O => \N__8891\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_2_2\
        );

    \I__1495\ : Odrv4
    port map (
            O => \N__8888\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_2_2\
        );

    \I__1494\ : CascadeMux
    port map (
            O => \N__8883\,
            I => \DUT.uart_inst0.recv_state_srsts_1_5_cascade_\
        );

    \I__1493\ : InMux
    port map (
            O => \N__8880\,
            I => \N__8877\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__8877\,
            I => \DUT.uart_inst0.recv_state_srsts_1_4\
        );

    \I__1491\ : InMux
    port map (
            O => \N__8874\,
            I => \N__8870\
        );

    \I__1490\ : InMux
    port map (
            O => \N__8873\,
            I => \N__8860\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__8870\,
            I => \N__8857\
        );

    \I__1488\ : InMux
    port map (
            O => \N__8869\,
            I => \N__8854\
        );

    \I__1487\ : InMux
    port map (
            O => \N__8868\,
            I => \N__8847\
        );

    \I__1486\ : InMux
    port map (
            O => \N__8867\,
            I => \N__8847\
        );

    \I__1485\ : InMux
    port map (
            O => \N__8866\,
            I => \N__8847\
        );

    \I__1484\ : InMux
    port map (
            O => \N__8865\,
            I => \N__8840\
        );

    \I__1483\ : InMux
    port map (
            O => \N__8864\,
            I => \N__8840\
        );

    \I__1482\ : InMux
    port map (
            O => \N__8863\,
            I => \N__8840\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__8860\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__1480\ : Odrv4
    port map (
            O => \N__8857\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__8854\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__8847\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__8840\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__1476\ : CascadeMux
    port map (
            O => \N__8829\,
            I => \DUT.uart_inst0.N_43_cascade_\
        );

    \I__1475\ : CEMux
    port map (
            O => \N__8826\,
            I => \N__8822\
        );

    \I__1474\ : CEMux
    port map (
            O => \N__8825\,
            I => \N__8819\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__8822\,
            I => \N__8816\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__8819\,
            I => \DUT.uart_inst0.recv_state_RNIL139CZ0Z_1\
        );

    \I__1471\ : Odrv4
    port map (
            O => \N__8816\,
            I => \DUT.uart_inst0.recv_state_RNIL139CZ0Z_1\
        );

    \I__1470\ : CascadeMux
    port map (
            O => \N__8811\,
            I => \DUT.uart_inst0.m3_e_1_cascade_\
        );

    \I__1469\ : CascadeMux
    port map (
            O => \N__8808\,
            I => \N__8805\
        );

    \I__1468\ : InMux
    port map (
            O => \N__8805\,
            I => \N__8802\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__8802\,
            I => \N__8795\
        );

    \I__1466\ : InMux
    port map (
            O => \N__8801\,
            I => \N__8792\
        );

    \I__1465\ : InMux
    port map (
            O => \N__8800\,
            I => \N__8789\
        );

    \I__1464\ : InMux
    port map (
            O => \N__8799\,
            I => \N__8780\
        );

    \I__1463\ : InMux
    port map (
            O => \N__8798\,
            I => \N__8777\
        );

    \I__1462\ : Span4Mux_h
    port map (
            O => \N__8795\,
            I => \N__8770\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__8792\,
            I => \N__8770\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__8789\,
            I => \N__8770\
        );

    \I__1459\ : InMux
    port map (
            O => \N__8788\,
            I => \N__8765\
        );

    \I__1458\ : InMux
    port map (
            O => \N__8787\,
            I => \N__8765\
        );

    \I__1457\ : InMux
    port map (
            O => \N__8786\,
            I => \N__8762\
        );

    \I__1456\ : InMux
    port map (
            O => \N__8785\,
            I => \N__8755\
        );

    \I__1455\ : InMux
    port map (
            O => \N__8784\,
            I => \N__8755\
        );

    \I__1454\ : InMux
    port map (
            O => \N__8783\,
            I => \N__8755\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__8780\,
            I => \DUT_uart_inst0_recv_state_2\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__8777\,
            I => \DUT_uart_inst0_recv_state_2\
        );

    \I__1451\ : Odrv4
    port map (
            O => \N__8770\,
            I => \DUT_uart_inst0_recv_state_2\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__8765\,
            I => \DUT_uart_inst0_recv_state_2\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__8762\,
            I => \DUT_uart_inst0_recv_state_2\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__8755\,
            I => \DUT_uart_inst0_recv_state_2\
        );

    \I__1447\ : InMux
    port map (
            O => \N__8742\,
            I => \N__8732\
        );

    \I__1446\ : InMux
    port map (
            O => \N__8741\,
            I => \N__8732\
        );

    \I__1445\ : InMux
    port map (
            O => \N__8740\,
            I => \N__8732\
        );

    \I__1444\ : CascadeMux
    port map (
            O => \N__8739\,
            I => \N__8726\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__8732\,
            I => \N__8723\
        );

    \I__1442\ : InMux
    port map (
            O => \N__8731\,
            I => \N__8714\
        );

    \I__1441\ : InMux
    port map (
            O => \N__8730\,
            I => \N__8714\
        );

    \I__1440\ : InMux
    port map (
            O => \N__8729\,
            I => \N__8714\
        );

    \I__1439\ : InMux
    port map (
            O => \N__8726\,
            I => \N__8714\
        );

    \I__1438\ : Odrv12
    port map (
            O => \N__8723\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_2\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__8714\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_2\
        );

    \I__1436\ : InMux
    port map (
            O => \N__8709\,
            I => \N__8704\
        );

    \I__1435\ : InMux
    port map (
            O => \N__8708\,
            I => \N__8699\
        );

    \I__1434\ : InMux
    port map (
            O => \N__8707\,
            I => \N__8699\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__8704\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_3\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__8699\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_3\
        );

    \I__1431\ : CascadeMux
    port map (
            O => \N__8694\,
            I => \N__8689\
        );

    \I__1430\ : InMux
    port map (
            O => \N__8693\,
            I => \N__8683\
        );

    \I__1429\ : InMux
    port map (
            O => \N__8692\,
            I => \N__8683\
        );

    \I__1428\ : InMux
    port map (
            O => \N__8689\,
            I => \N__8680\
        );

    \I__1427\ : CascadeMux
    port map (
            O => \N__8688\,
            I => \N__8673\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__8683\,
            I => \N__8668\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__8680\,
            I => \N__8668\
        );

    \I__1424\ : InMux
    port map (
            O => \N__8679\,
            I => \N__8663\
        );

    \I__1423\ : InMux
    port map (
            O => \N__8678\,
            I => \N__8663\
        );

    \I__1422\ : InMux
    port map (
            O => \N__8677\,
            I => \N__8656\
        );

    \I__1421\ : InMux
    port map (
            O => \N__8676\,
            I => \N__8656\
        );

    \I__1420\ : InMux
    port map (
            O => \N__8673\,
            I => \N__8656\
        );

    \I__1419\ : Odrv4
    port map (
            O => \N__8668\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_1\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__8663\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_1\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__8656\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_1\
        );

    \I__1416\ : InMux
    port map (
            O => \N__8649\,
            I => \N__8640\
        );

    \I__1415\ : InMux
    port map (
            O => \N__8648\,
            I => \N__8640\
        );

    \I__1414\ : InMux
    port map (
            O => \N__8647\,
            I => \N__8640\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__8640\,
            I => \N__8634\
        );

    \I__1412\ : InMux
    port map (
            O => \N__8639\,
            I => \N__8631\
        );

    \I__1411\ : InMux
    port map (
            O => \N__8638\,
            I => \N__8626\
        );

    \I__1410\ : InMux
    port map (
            O => \N__8637\,
            I => \N__8626\
        );

    \I__1409\ : Odrv4
    port map (
            O => \N__8634\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_0\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__8631\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_0\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__8626\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_0\
        );

    \I__1406\ : InMux
    port map (
            O => \N__8619\,
            I => \N__8616\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__8616\,
            I => \N__8613\
        );

    \I__1404\ : Span4Mux_v
    port map (
            O => \N__8613\,
            I => \N__8610\
        );

    \I__1403\ : Odrv4
    port map (
            O => \N__8610\,
            I => \DUT.uart_inst0.recv_state_RNO_4Z0Z_2\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__8607\,
            I => \DUT.uart_inst0.N_21_cascade_\
        );

    \I__1401\ : CascadeMux
    port map (
            O => \N__8604\,
            I => \DUT.uart_inst0.N_21_mux_cascade_\
        );

    \I__1400\ : InMux
    port map (
            O => \N__8601\,
            I => \N__8598\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__8598\,
            I => \DUT.uart_inst0.N_19_mux\
        );

    \I__1398\ : CascadeMux
    port map (
            O => \N__8595\,
            I => \DUT.uart_inst0.N_13_cascade_\
        );

    \I__1397\ : InMux
    port map (
            O => \N__8592\,
            I => \N__8589\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__8589\,
            I => \DUT.uart_inst0.N_13_0\
        );

    \I__1395\ : CascadeMux
    port map (
            O => \N__8586\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_2_0_2_cascade_\
        );

    \I__1394\ : InMux
    port map (
            O => \N__8583\,
            I => \N__8580\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__8580\,
            I => \DUT.fifo_tx_inst.un1_i11_i\
        );

    \I__1392\ : InMux
    port map (
            O => \N__8577\,
            I => \N__8574\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__8574\,
            I => \N__8571\
        );

    \I__1390\ : Odrv4
    port map (
            O => \N__8571\,
            I => \DUT.uart_inst0.g0_0\
        );

    \I__1389\ : InMux
    port map (
            O => \N__8568\,
            I => \N__8565\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__8565\,
            I => \DUT.uart_inst0.N_49\
        );

    \I__1387\ : InMux
    port map (
            O => \N__8562\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_0_s1\
        );

    \I__1386\ : InMux
    port map (
            O => \N__8559\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_1_s1\
        );

    \I__1385\ : InMux
    port map (
            O => \N__8556\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_2_s1\
        );

    \I__1384\ : InMux
    port map (
            O => \N__8553\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_3_s1\
        );

    \I__1383\ : InMux
    port map (
            O => \N__8550\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_4_s1\
        );

    \I__1382\ : InMux
    port map (
            O => \N__8547\,
            I => \N__8544\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__8544\,
            I => \N__8540\
        );

    \I__1380\ : InMux
    port map (
            O => \N__8543\,
            I => \N__8537\
        );

    \I__1379\ : Span4Mux_s1_v
    port map (
            O => \N__8540\,
            I => \N__8533\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__8537\,
            I => \N__8530\
        );

    \I__1377\ : InMux
    port map (
            O => \N__8536\,
            I => \N__8527\
        );

    \I__1376\ : Span4Mux_v
    port map (
            O => \N__8533\,
            I => \N__8524\
        );

    \I__1375\ : Span12Mux_s8_v
    port map (
            O => \N__8530\,
            I => \N__8521\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__8527\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_0\
        );

    \I__1373\ : Odrv4
    port map (
            O => \N__8524\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_0\
        );

    \I__1372\ : Odrv12
    port map (
            O => \N__8521\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_0\
        );

    \I__1371\ : SRMux
    port map (
            O => \N__8514\,
            I => \N__8510\
        );

    \I__1370\ : SRMux
    port map (
            O => \N__8513\,
            I => \N__8506\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__8510\,
            I => \N__8503\
        );

    \I__1368\ : SRMux
    port map (
            O => \N__8509\,
            I => \N__8500\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__8506\,
            I => \N__8497\
        );

    \I__1366\ : Span4Mux_s1_v
    port map (
            O => \N__8503\,
            I => \N__8492\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__8500\,
            I => \N__8492\
        );

    \I__1364\ : Span4Mux_h
    port map (
            O => \N__8497\,
            I => \N__8489\
        );

    \I__1363\ : Span4Mux_v
    port map (
            O => \N__8492\,
            I => \N__8486\
        );

    \I__1362\ : Span4Mux_v
    port map (
            O => \N__8489\,
            I => \N__8483\
        );

    \I__1361\ : Span4Mux_s1_v
    port map (
            O => \N__8486\,
            I => \N__8480\
        );

    \I__1360\ : Odrv4
    port map (
            O => \N__8483\,
            I => \DUT.uart_inst0.N_20\
        );

    \I__1359\ : Odrv4
    port map (
            O => \N__8480\,
            I => \DUT.uart_inst0.N_20\
        );

    \I__1358\ : InMux
    port map (
            O => \N__8475\,
            I => \N__8472\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__8472\,
            I => \N__8469\
        );

    \I__1356\ : Span4Mux_h
    port map (
            O => \N__8469\,
            I => \N__8466\
        );

    \I__1355\ : Odrv4
    port map (
            O => \N__8466\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO\
        );

    \I__1354\ : InMux
    port map (
            O => \N__8463\,
            I => \N__8459\
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__8462\,
            I => \N__8455\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__8459\,
            I => \N__8452\
        );

    \I__1351\ : InMux
    port map (
            O => \N__8458\,
            I => \N__8447\
        );

    \I__1350\ : InMux
    port map (
            O => \N__8455\,
            I => \N__8447\
        );

    \I__1349\ : Odrv4
    port map (
            O => \N__8452\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_4\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__8447\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_4\
        );

    \I__1347\ : CascadeMux
    port map (
            O => \N__8442\,
            I => \DUT.uart_inst0.m6_3_cascade_\
        );

    \I__1346\ : CascadeMux
    port map (
            O => \N__8439\,
            I => \top_pll_inst.m12_1_1_cascade_\
        );

    \I__1345\ : InMux
    port map (
            O => \N__8436\,
            I => \N__8433\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__8433\,
            I => \DUT.uart_inst0.G_30_1\
        );

    \I__1343\ : CascadeMux
    port map (
            O => \N__8430\,
            I => \P18_mux_cascade_\
        );

    \I__1342\ : InMux
    port map (
            O => \N__8427\,
            I => \N__8424\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__8424\,
            I => \N__8421\
        );

    \I__1340\ : Odrv4
    port map (
            O => \N__8421\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_11\
        );

    \I__1339\ : InMux
    port map (
            O => \N__8418\,
            I => \N__8415\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__8415\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_10\
        );

    \I__1337\ : CascadeMux
    port map (
            O => \N__8412\,
            I => \N__8409\
        );

    \I__1336\ : InMux
    port map (
            O => \N__8409\,
            I => \N__8406\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__8406\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_12\
        );

    \I__1334\ : InMux
    port map (
            O => \N__8403\,
            I => \N__8400\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__8400\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_13\
        );

    \I__1332\ : CascadeMux
    port map (
            O => \N__8397\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0_cascade_\
        );

    \I__1331\ : InMux
    port map (
            O => \N__8394\,
            I => \N__8387\
        );

    \I__1330\ : CascadeMux
    port map (
            O => \N__8393\,
            I => \N__8383\
        );

    \I__1329\ : CascadeMux
    port map (
            O => \N__8392\,
            I => \N__8379\
        );

    \I__1328\ : CascadeMux
    port map (
            O => \N__8391\,
            I => \N__8376\
        );

    \I__1327\ : InMux
    port map (
            O => \N__8390\,
            I => \N__8373\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__8387\,
            I => \N__8370\
        );

    \I__1325\ : CascadeMux
    port map (
            O => \N__8386\,
            I => \N__8366\
        );

    \I__1324\ : InMux
    port map (
            O => \N__8383\,
            I => \N__8358\
        );

    \I__1323\ : InMux
    port map (
            O => \N__8382\,
            I => \N__8355\
        );

    \I__1322\ : InMux
    port map (
            O => \N__8379\,
            I => \N__8352\
        );

    \I__1321\ : InMux
    port map (
            O => \N__8376\,
            I => \N__8349\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__8373\,
            I => \N__8344\
        );

    \I__1319\ : Span4Mux_s2_v
    port map (
            O => \N__8370\,
            I => \N__8344\
        );

    \I__1318\ : InMux
    port map (
            O => \N__8369\,
            I => \N__8341\
        );

    \I__1317\ : InMux
    port map (
            O => \N__8366\,
            I => \N__8334\
        );

    \I__1316\ : InMux
    port map (
            O => \N__8365\,
            I => \N__8334\
        );

    \I__1315\ : InMux
    port map (
            O => \N__8364\,
            I => \N__8334\
        );

    \I__1314\ : InMux
    port map (
            O => \N__8363\,
            I => \N__8327\
        );

    \I__1313\ : InMux
    port map (
            O => \N__8362\,
            I => \N__8327\
        );

    \I__1312\ : InMux
    port map (
            O => \N__8361\,
            I => \N__8327\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__8358\,
            I => \DUT.tx_state_1\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__8355\,
            I => \DUT.tx_state_1\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__8352\,
            I => \DUT.tx_state_1\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__8349\,
            I => \DUT.tx_state_1\
        );

    \I__1307\ : Odrv4
    port map (
            O => \N__8344\,
            I => \DUT.tx_state_1\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__8341\,
            I => \DUT.tx_state_1\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__8334\,
            I => \DUT.tx_state_1\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__8327\,
            I => \DUT.tx_state_1\
        );

    \I__1303\ : CascadeMux
    port map (
            O => \N__8310\,
            I => \DUT.N_114_cascade_\
        );

    \I__1302\ : CascadeMux
    port map (
            O => \N__8307\,
            I => \N__8304\
        );

    \I__1301\ : InMux
    port map (
            O => \N__8304\,
            I => \N__8294\
        );

    \I__1300\ : InMux
    port map (
            O => \N__8303\,
            I => \N__8289\
        );

    \I__1299\ : InMux
    port map (
            O => \N__8302\,
            I => \N__8289\
        );

    \I__1298\ : CascadeMux
    port map (
            O => \N__8301\,
            I => \N__8286\
        );

    \I__1297\ : InMux
    port map (
            O => \N__8300\,
            I => \N__8283\
        );

    \I__1296\ : CascadeMux
    port map (
            O => \N__8299\,
            I => \N__8280\
        );

    \I__1295\ : CascadeMux
    port map (
            O => \N__8298\,
            I => \N__8274\
        );

    \I__1294\ : CascadeMux
    port map (
            O => \N__8297\,
            I => \N__8269\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__8294\,
            I => \N__8256\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__8289\,
            I => \N__8253\
        );

    \I__1291\ : InMux
    port map (
            O => \N__8286\,
            I => \N__8247\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__8283\,
            I => \N__8244\
        );

    \I__1289\ : InMux
    port map (
            O => \N__8280\,
            I => \N__8239\
        );

    \I__1288\ : InMux
    port map (
            O => \N__8279\,
            I => \N__8239\
        );

    \I__1287\ : InMux
    port map (
            O => \N__8278\,
            I => \N__8236\
        );

    \I__1286\ : InMux
    port map (
            O => \N__8277\,
            I => \N__8233\
        );

    \I__1285\ : InMux
    port map (
            O => \N__8274\,
            I => \N__8228\
        );

    \I__1284\ : InMux
    port map (
            O => \N__8273\,
            I => \N__8228\
        );

    \I__1283\ : InMux
    port map (
            O => \N__8272\,
            I => \N__8223\
        );

    \I__1282\ : InMux
    port map (
            O => \N__8269\,
            I => \N__8223\
        );

    \I__1281\ : InMux
    port map (
            O => \N__8268\,
            I => \N__8218\
        );

    \I__1280\ : InMux
    port map (
            O => \N__8267\,
            I => \N__8218\
        );

    \I__1279\ : InMux
    port map (
            O => \N__8266\,
            I => \N__8201\
        );

    \I__1278\ : InMux
    port map (
            O => \N__8265\,
            I => \N__8201\
        );

    \I__1277\ : InMux
    port map (
            O => \N__8264\,
            I => \N__8201\
        );

    \I__1276\ : InMux
    port map (
            O => \N__8263\,
            I => \N__8201\
        );

    \I__1275\ : InMux
    port map (
            O => \N__8262\,
            I => \N__8201\
        );

    \I__1274\ : InMux
    port map (
            O => \N__8261\,
            I => \N__8201\
        );

    \I__1273\ : InMux
    port map (
            O => \N__8260\,
            I => \N__8201\
        );

    \I__1272\ : InMux
    port map (
            O => \N__8259\,
            I => \N__8201\
        );

    \I__1271\ : Span4Mux_s3_v
    port map (
            O => \N__8256\,
            I => \N__8196\
        );

    \I__1270\ : Span4Mux_h
    port map (
            O => \N__8253\,
            I => \N__8196\
        );

    \I__1269\ : InMux
    port map (
            O => \N__8252\,
            I => \N__8189\
        );

    \I__1268\ : InMux
    port map (
            O => \N__8251\,
            I => \N__8189\
        );

    \I__1267\ : InMux
    port map (
            O => \N__8250\,
            I => \N__8189\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__8247\,
            I => \N__8182\
        );

    \I__1265\ : Span4Mux_s2_v
    port map (
            O => \N__8244\,
            I => \N__8182\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__8239\,
            I => \N__8182\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__8236\,
            I => \DUT.tx_state_0\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__8233\,
            I => \DUT.tx_state_0\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__8228\,
            I => \DUT.tx_state_0\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__8223\,
            I => \DUT.tx_state_0\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__8218\,
            I => \DUT.tx_state_0\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__8201\,
            I => \DUT.tx_state_0\
        );

    \I__1257\ : Odrv4
    port map (
            O => \N__8196\,
            I => \DUT.tx_state_0\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__8189\,
            I => \DUT.tx_state_0\
        );

    \I__1255\ : Odrv4
    port map (
            O => \N__8182\,
            I => \DUT.tx_state_0\
        );

    \I__1254\ : CascadeMux
    port map (
            O => \N__8163\,
            I => \N__8160\
        );

    \I__1253\ : InMux
    port map (
            O => \N__8160\,
            I => \N__8157\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__8157\,
            I => \N__8152\
        );

    \I__1251\ : InMux
    port map (
            O => \N__8156\,
            I => \N__8149\
        );

    \I__1250\ : InMux
    port map (
            O => \N__8155\,
            I => \N__8146\
        );

    \I__1249\ : Odrv4
    port map (
            O => \N__8152\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_16\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__8149\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_16\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__8146\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_16\
        );

    \I__1246\ : CascadeMux
    port map (
            O => \N__8139\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_9_cascade_\
        );

    \I__1245\ : CascadeMux
    port map (
            O => \N__8136\,
            I => \N__8133\
        );

    \I__1244\ : InMux
    port map (
            O => \N__8133\,
            I => \N__8130\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__8130\,
            I => \N__8125\
        );

    \I__1242\ : InMux
    port map (
            O => \N__8129\,
            I => \N__8120\
        );

    \I__1241\ : InMux
    port map (
            O => \N__8128\,
            I => \N__8120\
        );

    \I__1240\ : Odrv4
    port map (
            O => \N__8125\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_1\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__8120\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_1\
        );

    \I__1238\ : InMux
    port map (
            O => \N__8115\,
            I => \N__8112\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__8112\,
            I => \N__8109\
        );

    \I__1236\ : Odrv4
    port map (
            O => \N__8109\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO\
        );

    \I__1235\ : InMux
    port map (
            O => \N__8106\,
            I => \N__8103\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__8103\,
            I => \N__8098\
        );

    \I__1233\ : InMux
    port map (
            O => \N__8102\,
            I => \N__8093\
        );

    \I__1232\ : InMux
    port map (
            O => \N__8101\,
            I => \N__8093\
        );

    \I__1231\ : Odrv4
    port map (
            O => \N__8098\,
            I => \DUT.uart_inst0.rx_clk_dividerZ1Z_1\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__8093\,
            I => \DUT.uart_inst0.rx_clk_dividerZ1Z_1\
        );

    \I__1229\ : InMux
    port map (
            O => \N__8088\,
            I => \N__8085\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__8085\,
            I => \N__8082\
        );

    \I__1227\ : Odrv4
    port map (
            O => \N__8082\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO\
        );

    \I__1226\ : InMux
    port map (
            O => \N__8079\,
            I => \N__8076\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__8076\,
            I => \N__8071\
        );

    \I__1224\ : InMux
    port map (
            O => \N__8075\,
            I => \N__8066\
        );

    \I__1223\ : InMux
    port map (
            O => \N__8074\,
            I => \N__8066\
        );

    \I__1222\ : Odrv4
    port map (
            O => \N__8071\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_2\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__8066\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_2\
        );

    \I__1220\ : InMux
    port map (
            O => \N__8061\,
            I => \N__8058\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__8058\,
            I => \N__8055\
        );

    \I__1218\ : Odrv12
    port map (
            O => \N__8055\,
            I => \DUT.uart_inst0.rx_clk_divider_1_3\
        );

    \I__1217\ : InMux
    port map (
            O => \N__8052\,
            I => \N__8049\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__8049\,
            I => \N__8045\
        );

    \I__1215\ : InMux
    port map (
            O => \N__8048\,
            I => \N__8042\
        );

    \I__1214\ : Odrv4
    port map (
            O => \N__8045\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_3\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__8042\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_3\
        );

    \I__1212\ : CascadeMux
    port map (
            O => \N__8037\,
            I => \N__8034\
        );

    \I__1211\ : InMux
    port map (
            O => \N__8034\,
            I => \N__8031\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__8031\,
            I => \DUT.uart_inst0.tx_dataZ0Z_1\
        );

    \I__1209\ : CascadeMux
    port map (
            O => \N__8028\,
            I => \N__8025\
        );

    \I__1208\ : InMux
    port map (
            O => \N__8025\,
            I => \N__8022\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__8022\,
            I => \DUT.uart_inst0.tx_dataZ0Z_2\
        );

    \I__1206\ : CascadeMux
    port map (
            O => \N__8019\,
            I => \N__8016\
        );

    \I__1205\ : InMux
    port map (
            O => \N__8016\,
            I => \N__8013\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__8013\,
            I => \N__8010\
        );

    \I__1203\ : Odrv4
    port map (
            O => \N__8010\,
            I => \DUT.uart_inst0.tx_dataZ0Z_3\
        );

    \I__1202\ : CascadeMux
    port map (
            O => \N__8007\,
            I => \N__8004\
        );

    \I__1201\ : InMux
    port map (
            O => \N__8004\,
            I => \N__8001\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__8001\,
            I => \DUT.uart_inst0.tx_dataZ0Z_4\
        );

    \I__1199\ : CascadeMux
    port map (
            O => \N__7998\,
            I => \N__7995\
        );

    \I__1198\ : InMux
    port map (
            O => \N__7995\,
            I => \N__7992\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__7992\,
            I => \DUT.uart_inst0.tx_dataZ0Z_5\
        );

    \I__1196\ : CascadeMux
    port map (
            O => \N__7989\,
            I => \N__7986\
        );

    \I__1195\ : InMux
    port map (
            O => \N__7986\,
            I => \N__7983\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__7983\,
            I => \DUT.uart_inst0.tx_dataZ0Z_7\
        );

    \I__1193\ : CascadeMux
    port map (
            O => \N__7980\,
            I => \N__7977\
        );

    \I__1192\ : InMux
    port map (
            O => \N__7977\,
            I => \N__7974\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__7974\,
            I => \DUT.uart_inst0.tx_dataZ0Z_6\
        );

    \I__1190\ : CEMux
    port map (
            O => \N__7971\,
            I => \N__7967\
        );

    \I__1189\ : CEMux
    port map (
            O => \N__7970\,
            I => \N__7964\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__7967\,
            I => \DUT.uart_inst0.N_22_i\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__7964\,
            I => \DUT.uart_inst0.N_22_i\
        );

    \I__1186\ : InMux
    port map (
            O => \N__7959\,
            I => \N__7950\
        );

    \I__1185\ : InMux
    port map (
            O => \N__7958\,
            I => \N__7950\
        );

    \I__1184\ : InMux
    port map (
            O => \N__7957\,
            I => \N__7950\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__7950\,
            I => \DUT.uart_inst0.N_102\
        );

    \I__1182\ : InMux
    port map (
            O => \N__7947\,
            I => \N__7944\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__7944\,
            I => \N__7941\
        );

    \I__1180\ : Span4Mux_h
    port map (
            O => \N__7941\,
            I => \N__7938\
        );

    \I__1179\ : Odrv4
    port map (
            O => \N__7938\,
            I => \DUT.uart_inst0.tx_state_0_sqmuxa_i_i_a3_0_1\
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__7935\,
            I => \G_110_cascade_\
        );

    \I__1177\ : InMux
    port map (
            O => \N__7932\,
            I => \N__7929\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__7929\,
            I => \fifo_inst_ftdi_input_inst_oTxFull_0\
        );

    \I__1175\ : InMux
    port map (
            O => \N__7926\,
            I => \N__7918\
        );

    \I__1174\ : InMux
    port map (
            O => \N__7925\,
            I => \N__7918\
        );

    \I__1173\ : InMux
    port map (
            O => \N__7924\,
            I => \N__7913\
        );

    \I__1172\ : InMux
    port map (
            O => \N__7923\,
            I => \N__7913\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__7918\,
            I => \G_108\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__7913\,
            I => \G_108\
        );

    \I__1169\ : InMux
    port map (
            O => \N__7908\,
            I => \N__7905\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__7905\,
            I => \fifo_inst.ftdi_input_inst.SUMZ0Z_3\
        );

    \I__1167\ : InMux
    port map (
            O => \N__7902\,
            I => \N__7893\
        );

    \I__1166\ : InMux
    port map (
            O => \N__7901\,
            I => \N__7893\
        );

    \I__1165\ : InMux
    port map (
            O => \N__7900\,
            I => \N__7886\
        );

    \I__1164\ : InMux
    port map (
            O => \N__7899\,
            I => \N__7886\
        );

    \I__1163\ : InMux
    port map (
            O => \N__7898\,
            I => \N__7886\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__7893\,
            I => \G_109\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__7886\,
            I => \G_109\
        );

    \I__1160\ : CascadeMux
    port map (
            O => \N__7881\,
            I => \N__7875\
        );

    \I__1159\ : CascadeMux
    port map (
            O => \N__7880\,
            I => \N__7872\
        );

    \I__1158\ : CascadeMux
    port map (
            O => \N__7879\,
            I => \N__7869\
        );

    \I__1157\ : InMux
    port map (
            O => \N__7878\,
            I => \N__7863\
        );

    \I__1156\ : InMux
    port map (
            O => \N__7875\,
            I => \N__7863\
        );

    \I__1155\ : InMux
    port map (
            O => \N__7872\,
            I => \N__7856\
        );

    \I__1154\ : InMux
    port map (
            O => \N__7869\,
            I => \N__7856\
        );

    \I__1153\ : InMux
    port map (
            O => \N__7868\,
            I => \N__7856\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__7863\,
            I => \G_110\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__7856\,
            I => \G_110\
        );

    \I__1150\ : CascadeMux
    port map (
            O => \N__7851\,
            I => \N__7848\
        );

    \I__1149\ : InMux
    port map (
            O => \N__7848\,
            I => \N__7840\
        );

    \I__1148\ : InMux
    port map (
            O => \N__7847\,
            I => \N__7840\
        );

    \I__1147\ : InMux
    port map (
            O => \N__7846\,
            I => \N__7835\
        );

    \I__1146\ : InMux
    port map (
            O => \N__7845\,
            I => \N__7835\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__7840\,
            I => \G_111\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__7835\,
            I => \G_111\
        );

    \I__1143\ : InMux
    port map (
            O => \N__7830\,
            I => \N__7821\
        );

    \I__1142\ : InMux
    port map (
            O => \N__7829\,
            I => \N__7821\
        );

    \I__1141\ : InMux
    port map (
            O => \N__7828\,
            I => \N__7814\
        );

    \I__1140\ : InMux
    port map (
            O => \N__7827\,
            I => \N__7814\
        );

    \I__1139\ : InMux
    port map (
            O => \N__7826\,
            I => \N__7814\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__7821\,
            I => \G_112\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__7814\,
            I => \G_112\
        );

    \I__1136\ : InMux
    port map (
            O => \N__7809\,
            I => \N__7806\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__7806\,
            I => \N__7803\
        );

    \I__1134\ : Span4Mux_h
    port map (
            O => \N__7803\,
            I => \N__7800\
        );

    \I__1133\ : Odrv4
    port map (
            O => \N__7800\,
            I => \fifo_inst.ftdi_input_inst.un2_oPacketAvail_iZ0\
        );

    \I__1132\ : InMux
    port map (
            O => \N__7797\,
            I => \N__7794\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__7794\,
            I => \N__7791\
        );

    \I__1130\ : Span4Mux_h
    port map (
            O => \N__7791\,
            I => \N__7787\
        );

    \I__1129\ : InMux
    port map (
            O => \N__7790\,
            I => \N__7784\
        );

    \I__1128\ : Odrv4
    port map (
            O => \N__7787\,
            I => \DUT.uart_inst0.tx_dataZ0Z_0\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__7784\,
            I => \DUT.uart_inst0.tx_dataZ0Z_0\
        );

    \I__1126\ : IoInMux
    port map (
            O => \N__7779\,
            I => \N__7775\
        );

    \I__1125\ : CascadeMux
    port map (
            O => \N__7778\,
            I => \N__7772\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__7775\,
            I => \N__7769\
        );

    \I__1123\ : InMux
    port map (
            O => \N__7772\,
            I => \N__7765\
        );

    \I__1122\ : Span4Mux_s3_v
    port map (
            O => \N__7769\,
            I => \N__7762\
        );

    \I__1121\ : InMux
    port map (
            O => \N__7768\,
            I => \N__7759\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__7765\,
            I => \N__7755\
        );

    \I__1119\ : Span4Mux_h
    port map (
            O => \N__7762\,
            I => \N__7752\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__7759\,
            I => \N__7749\
        );

    \I__1117\ : InMux
    port map (
            O => \N__7758\,
            I => \N__7746\
        );

    \I__1116\ : Span4Mux_v
    port map (
            O => \N__7755\,
            I => \N__7743\
        );

    \I__1115\ : Odrv4
    port map (
            O => \N__7752\,
            I => \P1A7_c\
        );

    \I__1114\ : Odrv4
    port map (
            O => \N__7749\,
            I => \P1A7_c\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__7746\,
            I => \P1A7_c\
        );

    \I__1112\ : Odrv4
    port map (
            O => \N__7743\,
            I => \P1A7_c\
        );

    \I__1111\ : InMux
    port map (
            O => \N__7734\,
            I => \N__7731\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__7731\,
            I => \N__7728\
        );

    \I__1109\ : Odrv12
    port map (
            O => \N__7728\,
            I => \DUT.uart_inst0.N_116\
        );

    \I__1108\ : CascadeMux
    port map (
            O => \N__7725\,
            I => \DUT.uart_inst0.m13_2_cascade_\
        );

    \I__1107\ : InMux
    port map (
            O => \N__7722\,
            I => \N__7719\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__7719\,
            I => \DUT.uart_inst0.m13_3\
        );

    \I__1105\ : CascadeMux
    port map (
            O => \N__7716\,
            I => \DUT.uart_inst0.P19_mux_cascade_\
        );

    \I__1104\ : InMux
    port map (
            O => \N__7713\,
            I => \N__7710\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__7710\,
            I => \N__7707\
        );

    \I__1102\ : Odrv4
    port map (
            O => \N__7707\,
            I => \DUT.uart_inst0.g0_0_1\
        );

    \I__1101\ : IoInMux
    port map (
            O => \N__7704\,
            I => \N__7701\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__7701\,
            I => \N__7698\
        );

    \I__1099\ : Span4Mux_s1_v
    port map (
            O => \N__7698\,
            I => \N__7695\
        );

    \I__1098\ : Odrv4
    port map (
            O => \N__7695\,
            I => \N_1257_i\
        );

    \I__1097\ : CascadeMux
    port map (
            O => \N__7692\,
            I => \G_111_cascade_\
        );

    \I__1096\ : CascadeMux
    port map (
            O => \N__7689\,
            I => \fifo_inst.ftdi_input_inst.SUMZ0Z_2_cascade_\
        );

    \I__1095\ : InMux
    port map (
            O => \N__7686\,
            I => \N__7683\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__7683\,
            I => \DUT.uart_inst0.g0_0_0_a3_0_4\
        );

    \I__1093\ : CascadeMux
    port map (
            O => \N__7680\,
            I => \DUT.uart_inst0.g0_0_0_a3_4_cascade_\
        );

    \I__1092\ : InMux
    port map (
            O => \N__7677\,
            I => \N__7674\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__7674\,
            I => \DUT.uart_inst0.g0_0_0_a3_3\
        );

    \I__1090\ : CascadeMux
    port map (
            O => \N__7671\,
            I => \DUT.fifo_tx_inst.un1_i11_i_cascade_\
        );

    \I__1089\ : CascadeMux
    port map (
            O => \N__7668\,
            I => \DUT.fifo_rx_inst.N_57_cascade_\
        );

    \I__1088\ : InMux
    port map (
            O => \N__7665\,
            I => \N__7659\
        );

    \I__1087\ : InMux
    port map (
            O => \N__7664\,
            I => \N__7659\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__7659\,
            I => \DUT.fifo_rx_inst.un1_i11_i\
        );

    \I__1085\ : CascadeMux
    port map (
            O => \N__7656\,
            I => \DUT.uart_inst0.N_21_0_cascade_\
        );

    \I__1084\ : InMux
    port map (
            O => \N__7653\,
            I => \N__7650\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__7650\,
            I => \DUT.uart_inst0.N_21_mux_0\
        );

    \I__1082\ : InMux
    port map (
            O => \N__7647\,
            I => \N__7644\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__7644\,
            I => \DUT.uart_inst0.m5_1\
        );

    \I__1080\ : InMux
    port map (
            O => \N__7641\,
            I => \N__7638\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__7638\,
            I => \DUT.uart_inst0.N_6\
        );

    \I__1078\ : CascadeMux
    port map (
            O => \N__7635\,
            I => \DUT.uart_inst0.N_6_cascade_\
        );

    \I__1077\ : InMux
    port map (
            O => \N__7632\,
            I => \N__7629\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__7629\,
            I => \N__7626\
        );

    \I__1075\ : Odrv4
    port map (
            O => \N__7626\,
            I => \DUT.uart_inst0.N_18\
        );

    \I__1074\ : InMux
    port map (
            O => \N__7623\,
            I => \N__7620\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__7620\,
            I => \DUT.uart_inst0.N_18_mux_0\
        );

    \I__1072\ : InMux
    port map (
            O => \N__7617\,
            I => \N__7614\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__7614\,
            I => \N__7611\
        );

    \I__1070\ : Span4Mux_h
    port map (
            O => \N__7611\,
            I => \N__7608\
        );

    \I__1069\ : Odrv4
    port map (
            O => \N__7608\,
            I => \DUT.uart_inst0.N_30\
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__7605\,
            I => \N__7602\
        );

    \I__1067\ : InMux
    port map (
            O => \N__7602\,
            I => \N__7599\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__7599\,
            I => \N__7596\
        );

    \I__1065\ : Odrv4
    port map (
            O => \N__7596\,
            I => \DUT.uart_inst0.g1_i_a4_0_4\
        );

    \I__1064\ : CascadeMux
    port map (
            O => \N__7593\,
            I => \DUT.uart_inst0.g1_i_a4_0_5_cascade_\
        );

    \I__1063\ : CascadeMux
    port map (
            O => \N__7590\,
            I => \DUT.uart_inst0.m7_e_1_cascade_\
        );

    \I__1062\ : CascadeMux
    port map (
            O => \N__7587\,
            I => \DUT.uart_inst0.m7_e_3_cascade_\
        );

    \I__1061\ : CascadeMux
    port map (
            O => \N__7584\,
            I => \DUT.uart_inst0.m9_1_cascade_\
        );

    \I__1060\ : InMux
    port map (
            O => \N__7581\,
            I => \N__7578\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__7578\,
            I => \DUT.uart_inst0.N_11_mux\
        );

    \I__1058\ : InMux
    port map (
            O => \N__7575\,
            I => \N__7572\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__7572\,
            I => \DUT.uart_inst0.N_66\
        );

    \I__1056\ : CascadeMux
    port map (
            O => \N__7569\,
            I => \N__7566\
        );

    \I__1055\ : InMux
    port map (
            O => \N__7566\,
            I => \N__7563\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__7563\,
            I => \N__7560\
        );

    \I__1053\ : Span4Mux_h
    port map (
            O => \N__7560\,
            I => \N__7557\
        );

    \I__1052\ : Odrv4
    port map (
            O => \N__7557\,
            I => \DUT.uart_inst0.m4_e_0\
        );

    \I__1051\ : InMux
    port map (
            O => \N__7554\,
            I => \N__7551\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__7551\,
            I => \DUT.uart_inst0.m4_e_3\
        );

    \I__1049\ : CascadeMux
    port map (
            O => \N__7548\,
            I => \N__7545\
        );

    \I__1048\ : InMux
    port map (
            O => \N__7545\,
            I => \N__7542\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__7542\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO\
        );

    \I__1046\ : InMux
    port map (
            O => \N__7539\,
            I => \N__7534\
        );

    \I__1045\ : InMux
    port map (
            O => \N__7538\,
            I => \N__7531\
        );

    \I__1044\ : InMux
    port map (
            O => \N__7537\,
            I => \N__7528\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__7534\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_11\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__7531\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_11\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__7528\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_11\
        );

    \I__1040\ : InMux
    port map (
            O => \N__7521\,
            I => \N__7518\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__7518\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO\
        );

    \I__1038\ : CascadeMux
    port map (
            O => \N__7515\,
            I => \N__7512\
        );

    \I__1037\ : InMux
    port map (
            O => \N__7512\,
            I => \N__7507\
        );

    \I__1036\ : InMux
    port map (
            O => \N__7511\,
            I => \N__7504\
        );

    \I__1035\ : InMux
    port map (
            O => \N__7510\,
            I => \N__7501\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__7507\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_7\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__7504\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_7\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__7501\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_7\
        );

    \I__1031\ : InMux
    port map (
            O => \N__7494\,
            I => \N__7491\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__7491\,
            I => \DUT.uart_inst0.rx_clk_divider_1_5\
        );

    \I__1029\ : InMux
    port map (
            O => \N__7488\,
            I => \N__7484\
        );

    \I__1028\ : InMux
    port map (
            O => \N__7487\,
            I => \N__7481\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__7484\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_5\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__7481\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_5\
        );

    \I__1025\ : InMux
    port map (
            O => \N__7476\,
            I => \N__7473\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__7473\,
            I => \DUT.uart_inst0.rx_clk_divider_1_6\
        );

    \I__1023\ : InMux
    port map (
            O => \N__7470\,
            I => \N__7466\
        );

    \I__1022\ : InMux
    port map (
            O => \N__7469\,
            I => \N__7463\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__7466\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_6\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__7463\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_6\
        );

    \I__1019\ : InMux
    port map (
            O => \N__7458\,
            I => \N__7455\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__7455\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO\
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__7452\,
            I => \N__7447\
        );

    \I__1016\ : InMux
    port map (
            O => \N__7451\,
            I => \N__7444\
        );

    \I__1015\ : InMux
    port map (
            O => \N__7450\,
            I => \N__7439\
        );

    \I__1014\ : InMux
    port map (
            O => \N__7447\,
            I => \N__7439\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__7444\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_8\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__7439\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_8\
        );

    \I__1011\ : InMux
    port map (
            O => \N__7434\,
            I => \N__7431\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__7431\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO\
        );

    \I__1009\ : CascadeMux
    port map (
            O => \N__7428\,
            I => \N__7423\
        );

    \I__1008\ : InMux
    port map (
            O => \N__7427\,
            I => \N__7420\
        );

    \I__1007\ : InMux
    port map (
            O => \N__7426\,
            I => \N__7417\
        );

    \I__1006\ : InMux
    port map (
            O => \N__7423\,
            I => \N__7414\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__7420\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_12\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__7417\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_12\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__7414\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_12\
        );

    \I__1002\ : InMux
    port map (
            O => \N__7407\,
            I => \N__7404\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__7404\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO\
        );

    \I__1000\ : CascadeMux
    port map (
            O => \N__7401\,
            I => \N__7398\
        );

    \I__999\ : InMux
    port map (
            O => \N__7398\,
            I => \N__7394\
        );

    \I__998\ : InMux
    port map (
            O => \N__7397\,
            I => \N__7391\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__7394\,
            I => \DUT.uart_inst0.tx_countdown_30_5\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__7391\,
            I => \DUT.uart_inst0.tx_countdown_30_5\
        );

    \I__995\ : InMux
    port map (
            O => \N__7386\,
            I => \N__7383\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__7383\,
            I => \N__7380\
        );

    \I__993\ : Odrv4
    port map (
            O => \N__7380\,
            I => \DUT.uart_inst0.tx_countdown_7_m1_0_a3_0_2\
        );

    \I__992\ : CascadeMux
    port map (
            O => \N__7377\,
            I => \N__7374\
        );

    \I__991\ : InMux
    port map (
            O => \N__7374\,
            I => \N__7371\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__7371\,
            I => \DUT.uart_inst0.N_113\
        );

    \I__989\ : InMux
    port map (
            O => \N__7368\,
            I => \N__7358\
        );

    \I__988\ : InMux
    port map (
            O => \N__7367\,
            I => \N__7358\
        );

    \I__987\ : InMux
    port map (
            O => \N__7366\,
            I => \N__7351\
        );

    \I__986\ : InMux
    port map (
            O => \N__7365\,
            I => \N__7351\
        );

    \I__985\ : InMux
    port map (
            O => \N__7364\,
            I => \N__7351\
        );

    \I__984\ : InMux
    port map (
            O => \N__7363\,
            I => \N__7348\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__7358\,
            I => \N__7345\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__7351\,
            I => \N__7342\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__7348\,
            I => \DUT.uart_inst0.tx_countdown_7_sm0_0\
        );

    \I__980\ : Odrv4
    port map (
            O => \N__7345\,
            I => \DUT.uart_inst0.tx_countdown_7_sm0_0\
        );

    \I__979\ : Odrv4
    port map (
            O => \N__7342\,
            I => \DUT.uart_inst0.tx_countdown_7_sm0_0\
        );

    \I__978\ : CascadeMux
    port map (
            O => \N__7335\,
            I => \N__7332\
        );

    \I__977\ : InMux
    port map (
            O => \N__7332\,
            I => \N__7328\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__7331\,
            I => \N__7325\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__7328\,
            I => \N__7322\
        );

    \I__974\ : InMux
    port map (
            O => \N__7325\,
            I => \N__7314\
        );

    \I__973\ : Span4Mux_s2_v
    port map (
            O => \N__7322\,
            I => \N__7311\
        );

    \I__972\ : InMux
    port map (
            O => \N__7321\,
            I => \N__7308\
        );

    \I__971\ : InMux
    port map (
            O => \N__7320\,
            I => \N__7303\
        );

    \I__970\ : InMux
    port map (
            O => \N__7319\,
            I => \N__7303\
        );

    \I__969\ : InMux
    port map (
            O => \N__7318\,
            I => \N__7298\
        );

    \I__968\ : InMux
    port map (
            O => \N__7317\,
            I => \N__7298\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__7314\,
            I => \DUT.uart_inst0.N_84\
        );

    \I__966\ : Odrv4
    port map (
            O => \N__7311\,
            I => \DUT.uart_inst0.N_84\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__7308\,
            I => \DUT.uart_inst0.N_84\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__7303\,
            I => \DUT.uart_inst0.N_84\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__7298\,
            I => \DUT.uart_inst0.N_84\
        );

    \I__962\ : CascadeMux
    port map (
            O => \N__7287\,
            I => \N__7283\
        );

    \I__961\ : CascadeMux
    port map (
            O => \N__7286\,
            I => \N__7280\
        );

    \I__960\ : InMux
    port map (
            O => \N__7283\,
            I => \N__7277\
        );

    \I__959\ : InMux
    port map (
            O => \N__7280\,
            I => \N__7274\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__7277\,
            I => \N__7271\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__7274\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_17\
        );

    \I__956\ : Odrv4
    port map (
            O => \N__7271\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_17\
        );

    \I__955\ : InMux
    port map (
            O => \N__7266\,
            I => \N__7263\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__7263\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO\
        );

    \I__953\ : InMux
    port map (
            O => \N__7260\,
            I => \N__7255\
        );

    \I__952\ : InMux
    port map (
            O => \N__7259\,
            I => \N__7252\
        );

    \I__951\ : InMux
    port map (
            O => \N__7258\,
            I => \N__7249\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__7255\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_13\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__7252\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_13\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__7249\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_13\
        );

    \I__947\ : InMux
    port map (
            O => \N__7242\,
            I => \N__7239\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__7239\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO\
        );

    \I__945\ : CascadeMux
    port map (
            O => \N__7236\,
            I => \N__7233\
        );

    \I__944\ : InMux
    port map (
            O => \N__7233\,
            I => \N__7228\
        );

    \I__943\ : InMux
    port map (
            O => \N__7232\,
            I => \N__7225\
        );

    \I__942\ : InMux
    port map (
            O => \N__7231\,
            I => \N__7222\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__7228\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_14\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__7225\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_14\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__7222\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_14\
        );

    \I__938\ : InMux
    port map (
            O => \N__7215\,
            I => \N__7212\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__7212\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO\
        );

    \I__936\ : InMux
    port map (
            O => \N__7209\,
            I => \N__7204\
        );

    \I__935\ : InMux
    port map (
            O => \N__7208\,
            I => \N__7199\
        );

    \I__934\ : InMux
    port map (
            O => \N__7207\,
            I => \N__7199\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__7204\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_15\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__7199\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_15\
        );

    \I__931\ : CascadeMux
    port map (
            O => \N__7194\,
            I => \N__7191\
        );

    \I__930\ : InMux
    port map (
            O => \N__7191\,
            I => \N__7188\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__7188\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO\
        );

    \I__928\ : InMux
    port map (
            O => \N__7185\,
            I => \N__7180\
        );

    \I__927\ : InMux
    port map (
            O => \N__7184\,
            I => \N__7175\
        );

    \I__926\ : InMux
    port map (
            O => \N__7183\,
            I => \N__7175\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__7180\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_10\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__7175\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_10\
        );

    \I__923\ : CascadeMux
    port map (
            O => \N__7170\,
            I => \N__7167\
        );

    \I__922\ : InMux
    port map (
            O => \N__7167\,
            I => \N__7164\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__7164\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO\
        );

    \I__920\ : InMux
    port map (
            O => \N__7161\,
            I => \N__7156\
        );

    \I__919\ : InMux
    port map (
            O => \N__7160\,
            I => \N__7151\
        );

    \I__918\ : InMux
    port map (
            O => \N__7159\,
            I => \N__7151\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__7156\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_9\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__7151\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_9\
        );

    \I__915\ : CascadeMux
    port map (
            O => \N__7146\,
            I => \DUT.uart_inst0.N_218_cascade_\
        );

    \I__914\ : InMux
    port map (
            O => \N__7143\,
            I => \N__7138\
        );

    \I__913\ : InMux
    port map (
            O => \N__7142\,
            I => \N__7133\
        );

    \I__912\ : InMux
    port map (
            O => \N__7141\,
            I => \N__7133\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__7138\,
            I => \DUT.uart_inst0.N_109\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__7133\,
            I => \DUT.uart_inst0.N_109\
        );

    \I__909\ : InMux
    port map (
            O => \N__7128\,
            I => \N__7115\
        );

    \I__908\ : InMux
    port map (
            O => \N__7127\,
            I => \N__7115\
        );

    \I__907\ : InMux
    port map (
            O => \N__7126\,
            I => \N__7110\
        );

    \I__906\ : InMux
    port map (
            O => \N__7125\,
            I => \N__7110\
        );

    \I__905\ : InMux
    port map (
            O => \N__7124\,
            I => \N__7105\
        );

    \I__904\ : InMux
    port map (
            O => \N__7123\,
            I => \N__7105\
        );

    \I__903\ : InMux
    port map (
            O => \N__7122\,
            I => \N__7098\
        );

    \I__902\ : InMux
    port map (
            O => \N__7121\,
            I => \N__7098\
        );

    \I__901\ : InMux
    port map (
            O => \N__7120\,
            I => \N__7098\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__7115\,
            I => \N__7095\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__7110\,
            I => \N__7088\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__7105\,
            I => \N__7088\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__7098\,
            I => \N__7088\
        );

    \I__896\ : Odrv4
    port map (
            O => \N__7095\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__895\ : Odrv4
    port map (
            O => \N__7088\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__894\ : CascadeMux
    port map (
            O => \N__7083\,
            I => \N__7077\
        );

    \I__893\ : InMux
    port map (
            O => \N__7082\,
            I => \N__7073\
        );

    \I__892\ : CascadeMux
    port map (
            O => \N__7081\,
            I => \N__7066\
        );

    \I__891\ : InMux
    port map (
            O => \N__7080\,
            I => \N__7061\
        );

    \I__890\ : InMux
    port map (
            O => \N__7077\,
            I => \N__7061\
        );

    \I__889\ : InMux
    port map (
            O => \N__7076\,
            I => \N__7058\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__7073\,
            I => \N__7055\
        );

    \I__887\ : InMux
    port map (
            O => \N__7072\,
            I => \N__7048\
        );

    \I__886\ : InMux
    port map (
            O => \N__7071\,
            I => \N__7048\
        );

    \I__885\ : InMux
    port map (
            O => \N__7070\,
            I => \N__7048\
        );

    \I__884\ : InMux
    port map (
            O => \N__7069\,
            I => \N__7043\
        );

    \I__883\ : InMux
    port map (
            O => \N__7066\,
            I => \N__7043\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__7061\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__7058\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__880\ : Odrv4
    port map (
            O => \N__7055\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__7048\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__7043\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__877\ : InMux
    port map (
            O => \N__7032\,
            I => \N__7029\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__7029\,
            I => \N__7025\
        );

    \I__875\ : InMux
    port map (
            O => \N__7028\,
            I => \N__7022\
        );

    \I__874\ : Odrv4
    port map (
            O => \N__7025\,
            I => \DUT.uart_inst0.N_120\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__7022\,
            I => \DUT.uart_inst0.N_120\
        );

    \I__872\ : CascadeMux
    port map (
            O => \N__7017\,
            I => \DUT.uart_inst0.tx_countdown_RNO_1Z0Z_3_cascade_\
        );

    \I__871\ : InMux
    port map (
            O => \N__7014\,
            I => \N__7005\
        );

    \I__870\ : InMux
    port map (
            O => \N__7013\,
            I => \N__7002\
        );

    \I__869\ : InMux
    port map (
            O => \N__7012\,
            I => \N__6989\
        );

    \I__868\ : InMux
    port map (
            O => \N__7011\,
            I => \N__6989\
        );

    \I__867\ : InMux
    port map (
            O => \N__7010\,
            I => \N__6989\
        );

    \I__866\ : InMux
    port map (
            O => \N__7009\,
            I => \N__6989\
        );

    \I__865\ : InMux
    port map (
            O => \N__7008\,
            I => \N__6986\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__7005\,
            I => \N__6983\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__7002\,
            I => \N__6980\
        );

    \I__862\ : InMux
    port map (
            O => \N__7001\,
            I => \N__6971\
        );

    \I__861\ : InMux
    port map (
            O => \N__7000\,
            I => \N__6971\
        );

    \I__860\ : InMux
    port map (
            O => \N__6999\,
            I => \N__6971\
        );

    \I__859\ : InMux
    port map (
            O => \N__6998\,
            I => \N__6971\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__6989\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__6986\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0\
        );

    \I__856\ : Odrv4
    port map (
            O => \N__6983\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0\
        );

    \I__855\ : Odrv4
    port map (
            O => \N__6980\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__6971\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0\
        );

    \I__853\ : InMux
    port map (
            O => \N__6960\,
            I => \N__6951\
        );

    \I__852\ : InMux
    port map (
            O => \N__6959\,
            I => \N__6951\
        );

    \I__851\ : InMux
    port map (
            O => \N__6958\,
            I => \N__6951\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__6951\,
            I => \DUT.uart_inst0.N_164\
        );

    \I__849\ : CascadeMux
    port map (
            O => \N__6948\,
            I => \DUT.uart_inst0.N_164_cascade_\
        );

    \I__848\ : InMux
    port map (
            O => \N__6945\,
            I => \N__6942\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__6942\,
            I => \DUT.uart_inst0.tx_countdown_RNO_0Z0Z_3\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__6939\,
            I => \N__6935\
        );

    \I__845\ : InMux
    port map (
            O => \N__6938\,
            I => \N__6928\
        );

    \I__844\ : InMux
    port map (
            O => \N__6935\,
            I => \N__6928\
        );

    \I__843\ : InMux
    port map (
            O => \N__6934\,
            I => \N__6923\
        );

    \I__842\ : InMux
    port map (
            O => \N__6933\,
            I => \N__6923\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__6928\,
            I => \N__6918\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__6923\,
            I => \N__6918\
        );

    \I__839\ : Odrv4
    port map (
            O => \N__6918\,
            I => \DUT.uart_inst0.tx_state_ns_i_i_o2_a0_2_0\
        );

    \I__838\ : InMux
    port map (
            O => \N__6915\,
            I => \N__6912\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__6912\,
            I => \N__6905\
        );

    \I__836\ : InMux
    port map (
            O => \N__6911\,
            I => \N__6900\
        );

    \I__835\ : InMux
    port map (
            O => \N__6910\,
            I => \N__6900\
        );

    \I__834\ : InMux
    port map (
            O => \N__6909\,
            I => \N__6895\
        );

    \I__833\ : InMux
    port map (
            O => \N__6908\,
            I => \N__6895\
        );

    \I__832\ : Span4Mux_v
    port map (
            O => \N__6905\,
            I => \N__6888\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__6900\,
            I => \N__6888\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__6895\,
            I => \N__6888\
        );

    \I__829\ : Odrv4
    port map (
            O => \N__6888\,
            I => \DUT.uart_inst0.N_159\
        );

    \I__828\ : InMux
    port map (
            O => \N__6885\,
            I => \N__6882\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__6882\,
            I => \N__6875\
        );

    \I__826\ : InMux
    port map (
            O => \N__6881\,
            I => \N__6870\
        );

    \I__825\ : InMux
    port map (
            O => \N__6880\,
            I => \N__6870\
        );

    \I__824\ : InMux
    port map (
            O => \N__6879\,
            I => \N__6867\
        );

    \I__823\ : InMux
    port map (
            O => \N__6878\,
            I => \N__6864\
        );

    \I__822\ : Span4Mux_s1_v
    port map (
            O => \N__6875\,
            I => \N__6859\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__6870\,
            I => \N__6859\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__6867\,
            I => \DUT.uart_inst0.N_100\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__6864\,
            I => \DUT.uart_inst0.N_100\
        );

    \I__818\ : Odrv4
    port map (
            O => \N__6859\,
            I => \DUT.uart_inst0.N_100\
        );

    \I__817\ : InMux
    port map (
            O => \N__6852\,
            I => \N__6849\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__6849\,
            I => \DUT.uart_inst0.N_163\
        );

    \I__815\ : InMux
    port map (
            O => \N__6846\,
            I => \N__6843\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__6843\,
            I => \N__6839\
        );

    \I__813\ : InMux
    port map (
            O => \N__6842\,
            I => \N__6832\
        );

    \I__812\ : Span4Mux_s2_v
    port map (
            O => \N__6839\,
            I => \N__6829\
        );

    \I__811\ : InMux
    port map (
            O => \N__6838\,
            I => \N__6824\
        );

    \I__810\ : InMux
    port map (
            O => \N__6837\,
            I => \N__6824\
        );

    \I__809\ : InMux
    port map (
            O => \N__6836\,
            I => \N__6819\
        );

    \I__808\ : InMux
    port map (
            O => \N__6835\,
            I => \N__6819\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__6832\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_5\
        );

    \I__806\ : Odrv4
    port map (
            O => \N__6829\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_5\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__6824\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_5\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__6819\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_5\
        );

    \I__803\ : CascadeMux
    port map (
            O => \N__6810\,
            I => \N__6807\
        );

    \I__802\ : InMux
    port map (
            O => \N__6807\,
            I => \N__6802\
        );

    \I__801\ : InMux
    port map (
            O => \N__6806\,
            I => \N__6797\
        );

    \I__800\ : InMux
    port map (
            O => \N__6805\,
            I => \N__6797\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__6802\,
            I => \DUT.uart_inst0.tx_countdown_0_c3\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__6797\,
            I => \DUT.uart_inst0.tx_countdown_0_c3\
        );

    \I__797\ : InMux
    port map (
            O => \N__6792\,
            I => \N__6785\
        );

    \I__796\ : CascadeMux
    port map (
            O => \N__6791\,
            I => \N__6781\
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__6790\,
            I => \N__6775\
        );

    \I__794\ : CascadeMux
    port map (
            O => \N__6789\,
            I => \N__6772\
        );

    \I__793\ : InMux
    port map (
            O => \N__6788\,
            I => \N__6769\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__6785\,
            I => \N__6766\
        );

    \I__791\ : InMux
    port map (
            O => \N__6784\,
            I => \N__6759\
        );

    \I__790\ : InMux
    port map (
            O => \N__6781\,
            I => \N__6759\
        );

    \I__789\ : InMux
    port map (
            O => \N__6780\,
            I => \N__6759\
        );

    \I__788\ : InMux
    port map (
            O => \N__6779\,
            I => \N__6750\
        );

    \I__787\ : InMux
    port map (
            O => \N__6778\,
            I => \N__6750\
        );

    \I__786\ : InMux
    port map (
            O => \N__6775\,
            I => \N__6750\
        );

    \I__785\ : InMux
    port map (
            O => \N__6772\,
            I => \N__6750\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__6769\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__783\ : Odrv4
    port map (
            O => \N__6766\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__6759\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__6750\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__780\ : CascadeMux
    port map (
            O => \N__6741\,
            I => \N__6737\
        );

    \I__779\ : InMux
    port map (
            O => \N__6740\,
            I => \N__6734\
        );

    \I__778\ : InMux
    port map (
            O => \N__6737\,
            I => \N__6725\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__6734\,
            I => \N__6722\
        );

    \I__776\ : InMux
    port map (
            O => \N__6733\,
            I => \N__6713\
        );

    \I__775\ : InMux
    port map (
            O => \N__6732\,
            I => \N__6713\
        );

    \I__774\ : InMux
    port map (
            O => \N__6731\,
            I => \N__6713\
        );

    \I__773\ : InMux
    port map (
            O => \N__6730\,
            I => \N__6713\
        );

    \I__772\ : InMux
    port map (
            O => \N__6729\,
            I => \N__6708\
        );

    \I__771\ : InMux
    port map (
            O => \N__6728\,
            I => \N__6708\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__6725\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_4\
        );

    \I__769\ : Odrv4
    port map (
            O => \N__6722\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_4\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__6713\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_4\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__6708\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_4\
        );

    \I__766\ : CascadeMux
    port map (
            O => \N__6699\,
            I => \DUT.uart_inst0.N_160_cascade_\
        );

    \I__765\ : InMux
    port map (
            O => \N__6696\,
            I => \N__6688\
        );

    \I__764\ : InMux
    port map (
            O => \N__6695\,
            I => \N__6688\
        );

    \I__763\ : InMux
    port map (
            O => \N__6694\,
            I => \N__6683\
        );

    \I__762\ : InMux
    port map (
            O => \N__6693\,
            I => \N__6683\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__6688\,
            I => \DUT.uart_inst0.tx_countdown_0_ac0_1\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__6683\,
            I => \DUT.uart_inst0.tx_countdown_0_ac0_1\
        );

    \I__759\ : InMux
    port map (
            O => \N__6678\,
            I => \N__6675\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__6675\,
            I => \DUT.uart_inst0.N_154\
        );

    \I__757\ : CascadeMux
    port map (
            O => \N__6672\,
            I => \N__6666\
        );

    \I__756\ : InMux
    port map (
            O => \N__6671\,
            I => \N__6662\
        );

    \I__755\ : InMux
    port map (
            O => \N__6670\,
            I => \N__6657\
        );

    \I__754\ : InMux
    port map (
            O => \N__6669\,
            I => \N__6657\
        );

    \I__753\ : InMux
    port map (
            O => \N__6666\,
            I => \N__6654\
        );

    \I__752\ : InMux
    port map (
            O => \N__6665\,
            I => \N__6651\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__6662\,
            I => \N__6648\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__6657\,
            I => \N__6645\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__6654\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_3\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__6651\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_3\
        );

    \I__747\ : Odrv4
    port map (
            O => \N__6648\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_3\
        );

    \I__746\ : Odrv4
    port map (
            O => \N__6645\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_3\
        );

    \I__745\ : InMux
    port map (
            O => \N__6636\,
            I => \N__6633\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__6633\,
            I => \DUT.uart_inst0.N_72\
        );

    \I__743\ : InMux
    port map (
            O => \N__6630\,
            I => \N__6626\
        );

    \I__742\ : InMux
    port map (
            O => \N__6629\,
            I => \N__6623\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__6626\,
            I => \DUT.uart_inst0.N_99\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__6623\,
            I => \DUT.uart_inst0.N_99\
        );

    \I__739\ : InMux
    port map (
            O => \N__6618\,
            I => \N__6615\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__6615\,
            I => \N__6612\
        );

    \I__737\ : Span4Mux_s3_v
    port map (
            O => \N__6612\,
            I => \N__6609\
        );

    \I__736\ : Odrv4
    port map (
            O => \N__6609\,
            I => \DUT.uart_inst0.tx_countdown_RNO_0Z0Z_1\
        );

    \I__735\ : SRMux
    port map (
            O => \N__6606\,
            I => \N__6602\
        );

    \I__734\ : SRMux
    port map (
            O => \N__6605\,
            I => \N__6599\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__6602\,
            I => \N__6594\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__6599\,
            I => \N__6594\
        );

    \I__731\ : Span4Mux_v
    port map (
            O => \N__6594\,
            I => \N__6591\
        );

    \I__730\ : Span4Mux_h
    port map (
            O => \N__6591\,
            I => \N__6588\
        );

    \I__729\ : Odrv4
    port map (
            O => \N__6588\,
            I => \DUT.uart_inst0.N_88_i\
        );

    \I__728\ : CascadeMux
    port map (
            O => \N__6585\,
            I => \N__6581\
        );

    \I__727\ : InMux
    port map (
            O => \N__6584\,
            I => \N__6577\
        );

    \I__726\ : InMux
    port map (
            O => \N__6581\,
            I => \N__6574\
        );

    \I__725\ : InMux
    port map (
            O => \N__6580\,
            I => \N__6571\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__6577\,
            I => \DUT.uart_inst0.N_160\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__6574\,
            I => \DUT.uart_inst0.N_160\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__6571\,
            I => \DUT.uart_inst0.N_160\
        );

    \I__721\ : InMux
    port map (
            O => \N__6564\,
            I => \N__6561\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__6561\,
            I => \DUT.uart_inst0.N_218\
        );

    \I__719\ : InMux
    port map (
            O => \N__6558\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_8\
        );

    \I__718\ : InMux
    port map (
            O => \N__6555\,
            I => \N__6551\
        );

    \I__717\ : InMux
    port map (
            O => \N__6554\,
            I => \N__6548\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__6551\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_10\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__6548\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_10\
        );

    \I__714\ : InMux
    port map (
            O => \N__6543\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_9\
        );

    \I__713\ : CascadeMux
    port map (
            O => \N__6540\,
            I => \N__6536\
        );

    \I__712\ : InMux
    port map (
            O => \N__6539\,
            I => \N__6533\
        );

    \I__711\ : InMux
    port map (
            O => \N__6536\,
            I => \N__6530\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__6533\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_11\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__6530\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_11\
        );

    \I__708\ : InMux
    port map (
            O => \N__6525\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_10\
        );

    \I__707\ : InMux
    port map (
            O => \N__6522\,
            I => \N__6518\
        );

    \I__706\ : InMux
    port map (
            O => \N__6521\,
            I => \N__6515\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__6518\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_12\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__6515\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_12\
        );

    \I__703\ : InMux
    port map (
            O => \N__6510\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_11\
        );

    \I__702\ : InMux
    port map (
            O => \N__6507\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_12\
        );

    \I__701\ : CascadeMux
    port map (
            O => \N__6504\,
            I => \N__6500\
        );

    \I__700\ : InMux
    port map (
            O => \N__6503\,
            I => \N__6497\
        );

    \I__699\ : InMux
    port map (
            O => \N__6500\,
            I => \N__6494\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__6497\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_13\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__6494\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_13\
        );

    \I__696\ : InMux
    port map (
            O => \N__6489\,
            I => \N__6486\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__6486\,
            I => \N__6480\
        );

    \I__694\ : InMux
    port map (
            O => \N__6485\,
            I => \N__6473\
        );

    \I__693\ : InMux
    port map (
            O => \N__6484\,
            I => \N__6473\
        );

    \I__692\ : InMux
    port map (
            O => \N__6483\,
            I => \N__6473\
        );

    \I__691\ : Odrv4
    port map (
            O => \N__6480\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_2\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__6473\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_2\
        );

    \I__689\ : InMux
    port map (
            O => \N__6468\,
            I => \N__6465\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__6465\,
            I => \N__6461\
        );

    \I__687\ : InMux
    port map (
            O => \N__6464\,
            I => \N__6455\
        );

    \I__686\ : Span4Mux_v
    port map (
            O => \N__6461\,
            I => \N__6452\
        );

    \I__685\ : InMux
    port map (
            O => \N__6460\,
            I => \N__6445\
        );

    \I__684\ : InMux
    port map (
            O => \N__6459\,
            I => \N__6445\
        );

    \I__683\ : InMux
    port map (
            O => \N__6458\,
            I => \N__6445\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__6455\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_1\
        );

    \I__681\ : Odrv4
    port map (
            O => \N__6452\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_1\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__6445\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_1\
        );

    \I__679\ : InMux
    port map (
            O => \N__6438\,
            I => \N__6435\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__6435\,
            I => \N__6432\
        );

    \I__677\ : Odrv4
    port map (
            O => \N__6432\,
            I => \DUT.uart_inst0.m9_e_0_3\
        );

    \I__676\ : InMux
    port map (
            O => \N__6429\,
            I => \N__6423\
        );

    \I__675\ : CascadeMux
    port map (
            O => \N__6428\,
            I => \N__6418\
        );

    \I__674\ : CascadeMux
    port map (
            O => \N__6427\,
            I => \N__6415\
        );

    \I__673\ : InMux
    port map (
            O => \N__6426\,
            I => \N__6412\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__6423\,
            I => \N__6409\
        );

    \I__671\ : InMux
    port map (
            O => \N__6422\,
            I => \N__6400\
        );

    \I__670\ : InMux
    port map (
            O => \N__6421\,
            I => \N__6400\
        );

    \I__669\ : InMux
    port map (
            O => \N__6418\,
            I => \N__6400\
        );

    \I__668\ : InMux
    port map (
            O => \N__6415\,
            I => \N__6400\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__6412\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_0\
        );

    \I__666\ : Odrv4
    port map (
            O => \N__6409\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_0\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__6400\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_0\
        );

    \I__664\ : InMux
    port map (
            O => \N__6393\,
            I => \N__6390\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__6390\,
            I => \DUT.uart_inst0.m9_e_0_0\
        );

    \I__662\ : InMux
    port map (
            O => \N__6387\,
            I => \N__6383\
        );

    \I__661\ : InMux
    port map (
            O => \N__6386\,
            I => \N__6380\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__6383\,
            I => \DUT.uart_inst0.N_152\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__6380\,
            I => \DUT.uart_inst0.N_152\
        );

    \I__658\ : CascadeMux
    port map (
            O => \N__6375\,
            I => \DUT.uart_inst0.tx_state_0_sqmuxa_i_i_a3_c_cascade_\
        );

    \I__657\ : InMux
    port map (
            O => \N__6372\,
            I => \N__6368\
        );

    \I__656\ : InMux
    port map (
            O => \N__6371\,
            I => \N__6365\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__6368\,
            I => \N__6362\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__6365\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_1\
        );

    \I__653\ : Odrv4
    port map (
            O => \N__6362\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_1\
        );

    \I__652\ : InMux
    port map (
            O => \N__6357\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_0\
        );

    \I__651\ : CascadeMux
    port map (
            O => \N__6354\,
            I => \N__6350\
        );

    \I__650\ : InMux
    port map (
            O => \N__6353\,
            I => \N__6347\
        );

    \I__649\ : InMux
    port map (
            O => \N__6350\,
            I => \N__6344\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__6347\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_2\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__6344\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_2\
        );

    \I__646\ : InMux
    port map (
            O => \N__6339\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_1\
        );

    \I__645\ : InMux
    port map (
            O => \N__6336\,
            I => \N__6332\
        );

    \I__644\ : InMux
    port map (
            O => \N__6335\,
            I => \N__6329\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__6332\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_3\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__6329\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_3\
        );

    \I__641\ : InMux
    port map (
            O => \N__6324\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_2\
        );

    \I__640\ : InMux
    port map (
            O => \N__6321\,
            I => \N__6317\
        );

    \I__639\ : InMux
    port map (
            O => \N__6320\,
            I => \N__6314\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__6317\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_4\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__6314\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_4\
        );

    \I__636\ : InMux
    port map (
            O => \N__6309\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_3\
        );

    \I__635\ : InMux
    port map (
            O => \N__6306\,
            I => \N__6302\
        );

    \I__634\ : InMux
    port map (
            O => \N__6305\,
            I => \N__6299\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__6302\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_5\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__6299\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_5\
        );

    \I__631\ : InMux
    port map (
            O => \N__6294\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_4\
        );

    \I__630\ : InMux
    port map (
            O => \N__6291\,
            I => \N__6287\
        );

    \I__629\ : InMux
    port map (
            O => \N__6290\,
            I => \N__6284\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__6287\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_6\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__6284\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_6\
        );

    \I__626\ : InMux
    port map (
            O => \N__6279\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_5\
        );

    \I__625\ : InMux
    port map (
            O => \N__6276\,
            I => \N__6272\
        );

    \I__624\ : InMux
    port map (
            O => \N__6275\,
            I => \N__6269\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__6272\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_7\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__6269\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_7\
        );

    \I__621\ : InMux
    port map (
            O => \N__6264\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_6\
        );

    \I__620\ : InMux
    port map (
            O => \N__6261\,
            I => \N__6257\
        );

    \I__619\ : InMux
    port map (
            O => \N__6260\,
            I => \N__6254\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__6257\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_8\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__6254\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_8\
        );

    \I__616\ : InMux
    port map (
            O => \N__6249\,
            I => \bfn_14_3_0_\
        );

    \I__615\ : InMux
    port map (
            O => \N__6246\,
            I => \N__6242\
        );

    \I__614\ : InMux
    port map (
            O => \N__6245\,
            I => \N__6239\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__6242\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_9\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__6239\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_9\
        );

    \I__611\ : CascadeMux
    port map (
            O => \N__6234\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_1_2_cascade_\
        );

    \I__610\ : InMux
    port map (
            O => \N__6231\,
            I => \N__6228\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__6228\,
            I => \DUT.uart_inst0.N_67\
        );

    \I__608\ : CascadeMux
    port map (
            O => \N__6225\,
            I => \DUT.uart_inst0.g0_0_0_a3_0_3_cascade_\
        );

    \I__607\ : InMux
    port map (
            O => \N__6222\,
            I => \N__6219\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__6219\,
            I => \DUT.uart_inst0.N_159_0\
        );

    \I__605\ : InMux
    port map (
            O => \N__6216\,
            I => \N__6213\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__6213\,
            I => \DUT.uart_inst0.N_4\
        );

    \I__603\ : InMux
    port map (
            O => \N__6210\,
            I => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0\
        );

    \I__602\ : InMux
    port map (
            O => \N__6207\,
            I => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1\
        );

    \I__601\ : InMux
    port map (
            O => \N__6204\,
            I => \N__6201\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__6201\,
            I => \DUT.fifo_tx_inst.rFifoCount_RNISSQ21Z0Z_1\
        );

    \I__599\ : CascadeMux
    port map (
            O => \N__6198\,
            I => \DUT.fifo_tx_inst.N_108_cascade_\
        );

    \I__598\ : InMux
    port map (
            O => \N__6195\,
            I => \N__6192\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__6192\,
            I => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0\
        );

    \I__596\ : InMux
    port map (
            O => \N__6189\,
            I => \N__6184\
        );

    \I__595\ : InMux
    port map (
            O => \N__6188\,
            I => \N__6179\
        );

    \I__594\ : InMux
    port map (
            O => \N__6187\,
            I => \N__6179\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__6184\,
            I => \DUT.fifo_tx_inst.N_108\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__6179\,
            I => \DUT.fifo_tx_inst.N_108\
        );

    \I__591\ : CascadeMux
    port map (
            O => \N__6174\,
            I => \N__6170\
        );

    \I__590\ : CascadeMux
    port map (
            O => \N__6173\,
            I => \N__6167\
        );

    \I__589\ : InMux
    port map (
            O => \N__6170\,
            I => \N__6159\
        );

    \I__588\ : InMux
    port map (
            O => \N__6167\,
            I => \N__6159\
        );

    \I__587\ : InMux
    port map (
            O => \N__6166\,
            I => \N__6159\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__6159\,
            I => \rTxWriteZ0\
        );

    \I__585\ : CascadeMux
    port map (
            O => \N__6156\,
            I => \DUT.fifo_tx_inst.N_104_cascade_\
        );

    \I__584\ : InMux
    port map (
            O => \N__6153\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_9\
        );

    \I__583\ : InMux
    port map (
            O => \N__6150\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_10\
        );

    \I__582\ : InMux
    port map (
            O => \N__6147\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_11\
        );

    \I__581\ : InMux
    port map (
            O => \N__6144\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_12\
        );

    \I__580\ : InMux
    port map (
            O => \N__6141\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_13\
        );

    \I__579\ : InMux
    port map (
            O => \N__6138\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_14\
        );

    \I__578\ : InMux
    port map (
            O => \N__6135\,
            I => \bfn_13_9_0_\
        );

    \I__577\ : InMux
    port map (
            O => \N__6132\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_16\
        );

    \I__576\ : InMux
    port map (
            O => \N__6129\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_0\
        );

    \I__575\ : InMux
    port map (
            O => \N__6126\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_1\
        );

    \I__574\ : InMux
    port map (
            O => \N__6123\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_2\
        );

    \I__573\ : InMux
    port map (
            O => \N__6120\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_3\
        );

    \I__572\ : InMux
    port map (
            O => \N__6117\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_4\
        );

    \I__571\ : InMux
    port map (
            O => \N__6114\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_5\
        );

    \I__570\ : InMux
    port map (
            O => \N__6111\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_6\
        );

    \I__569\ : InMux
    port map (
            O => \N__6108\,
            I => \bfn_13_8_0_\
        );

    \I__568\ : InMux
    port map (
            O => \N__6105\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_8\
        );

    \I__567\ : CascadeMux
    port map (
            O => \N__6102\,
            I => \DUT.uart_inst0.tx_countdown_RNO_0Z0Z_4_cascade_\
        );

    \I__566\ : CascadeMux
    port map (
            O => \N__6099\,
            I => \DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0_cascade_\
        );

    \I__565\ : CascadeMux
    port map (
            O => \N__6096\,
            I => \DUT.uart_inst0.m25_e_3_cascade_\
        );

    \I__564\ : CascadeMux
    port map (
            O => \N__6093\,
            I => \N__6090\
        );

    \I__563\ : InMux
    port map (
            O => \N__6090\,
            I => \N__6087\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__6087\,
            I => \N__6084\
        );

    \I__561\ : Odrv4
    port map (
            O => \N__6084\,
            I => \DUT.uart_inst0.m3_0\
        );

    \I__560\ : InMux
    port map (
            O => \N__6081\,
            I => \N__6078\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__6078\,
            I => \DUT.uart_inst0.N_5\
        );

    \I__558\ : CascadeMux
    port map (
            O => \N__6075\,
            I => \DUT.uart_inst0.tx_countdown_7_m1_0_o2_2_2_cascade_\
        );

    \I__557\ : CascadeMux
    port map (
            O => \N__6072\,
            I => \DUT.uart_inst0.tx_out_6_iv_0_a3_0_1_cascade_\
        );

    \I__556\ : CascadeMux
    port map (
            O => \N__6069\,
            I => \DUT.uart_inst0.tx_out_6_iv_0_1_cascade_\
        );

    \I__555\ : InMux
    port map (
            O => \N__6066\,
            I => \N__6063\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__6063\,
            I => \DUT.uart_inst0.N_119\
        );

    \I__553\ : CascadeMux
    port map (
            O => \N__6060\,
            I => \DUT.uart_inst0.g2_3_cascade_\
        );

    \I__552\ : InMux
    port map (
            O => \N__6057\,
            I => \N__6054\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__6054\,
            I => \DUT.uart_inst0.g2\
        );

    \I__550\ : InMux
    port map (
            O => \N__6051\,
            I => \N__6048\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__6048\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_9\
        );

    \I__548\ : InMux
    port map (
            O => \N__6045\,
            I => \N__6042\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__6042\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_8\
        );

    \I__546\ : CascadeMux
    port map (
            O => \N__6039\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_6_cascade_\
        );

    \I__545\ : InMux
    port map (
            O => \N__6036\,
            I => \N__6033\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__6033\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_7\
        );

    \I__543\ : CascadeMux
    port map (
            O => \N__6030\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0_cascade_\
        );

    \I__542\ : CascadeMux
    port map (
            O => \N__6027\,
            I => \DUT.uart_inst0.N_152_cascade_\
        );

    \I__541\ : CascadeMux
    port map (
            O => \N__6024\,
            I => \DUT.uart_inst0.N_6_0_cascade_\
        );

    \I__540\ : CascadeMux
    port map (
            O => \N__6021\,
            I => \DUT.uart_inst0.N_22_cascade_\
        );

    \I__539\ : CascadeMux
    port map (
            O => \N__6018\,
            I => \N__6015\
        );

    \I__538\ : InMux
    port map (
            O => \N__6015\,
            I => \N__6009\
        );

    \I__537\ : InMux
    port map (
            O => \N__6014\,
            I => \N__6009\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__6009\,
            I => \DUT.uart_inst0.N_22\
        );

    \I__535\ : IoInMux
    port map (
            O => \N__6006\,
            I => \N__6003\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__6003\,
            I => \N__6000\
        );

    \I__533\ : IoSpan4Mux
    port map (
            O => \N__6000\,
            I => \N__5997\
        );

    \I__532\ : Sp12to4
    port map (
            O => \N__5997\,
            I => \N__5994\
        );

    \I__531\ : Span12Mux_s7_v
    port map (
            O => \N__5994\,
            I => \N__5991\
        );

    \I__530\ : Odrv12
    port map (
            O => \N__5991\,
            I => \wRamRdData_0\
        );

    \I__529\ : IoInMux
    port map (
            O => \N__5988\,
            I => \N__5985\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__5985\,
            I => \N__5982\
        );

    \I__527\ : Span4Mux_s3_v
    port map (
            O => \N__5982\,
            I => \N__5979\
        );

    \I__526\ : Span4Mux_v
    port map (
            O => \N__5979\,
            I => \N__5976\
        );

    \I__525\ : Odrv4
    port map (
            O => \N__5976\,
            I => \wRamRdData_3\
        );

    \I__524\ : InMux
    port map (
            O => \N__5973\,
            I => \N__5970\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__5970\,
            I => \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO\
        );

    \I__522\ : IoInMux
    port map (
            O => \N__5967\,
            I => \N__5964\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__5964\,
            I => \top_pll_inst.wPllLocked_iso_i\
        );

    \I__520\ : IoInMux
    port map (
            O => \N__5961\,
            I => \N__5958\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__5958\,
            I => \N__5955\
        );

    \I__518\ : Span12Mux_s1_v
    port map (
            O => \N__5955\,
            I => \N__5952\
        );

    \I__517\ : Odrv12
    port map (
            O => \N__5952\,
            I => \wRamRdData_4\
        );

    \I__516\ : IoInMux
    port map (
            O => \N__5949\,
            I => \N__5946\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__5946\,
            I => \N__5943\
        );

    \I__514\ : Span12Mux_s9_v
    port map (
            O => \N__5943\,
            I => \N__5940\
        );

    \I__513\ : Span12Mux_v
    port map (
            O => \N__5940\,
            I => \N__5937\
        );

    \I__512\ : Odrv12
    port map (
            O => \N__5937\,
            I => \BTN_N_c\
        );

    \I__511\ : IoInMux
    port map (
            O => \N__5934\,
            I => \N__5931\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__5931\,
            I => \N__5928\
        );

    \I__509\ : Span12Mux_s2_v
    port map (
            O => \N__5928\,
            I => \N__5925\
        );

    \I__508\ : Span12Mux_v
    port map (
            O => \N__5925\,
            I => \N__5922\
        );

    \I__507\ : Odrv12
    port map (
            O => \N__5922\,
            I => \wRamRdData_7\
        );

    \I__506\ : IoInMux
    port map (
            O => \N__5919\,
            I => \N__5916\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__5916\,
            I => \N__5913\
        );

    \I__504\ : IoSpan4Mux
    port map (
            O => \N__5913\,
            I => \N__5910\
        );

    \I__503\ : Sp12to4
    port map (
            O => \N__5910\,
            I => \N__5907\
        );

    \I__502\ : Span12Mux_s7_v
    port map (
            O => \N__5907\,
            I => \N__5904\
        );

    \I__501\ : Odrv12
    port map (
            O => \N__5904\,
            I => \wRamRdData_1\
        );

    \I__500\ : IoInMux
    port map (
            O => \N__5901\,
            I => \N__5898\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__5898\,
            I => \N__5895\
        );

    \I__498\ : Sp12to4
    port map (
            O => \N__5895\,
            I => \N__5892\
        );

    \I__497\ : Span12Mux_v
    port map (
            O => \N__5892\,
            I => \N__5889\
        );

    \I__496\ : Odrv12
    port map (
            O => \N__5889\,
            I => \wRamRdData_6\
        );

    \I__495\ : IoInMux
    port map (
            O => \N__5886\,
            I => \N__5883\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__5883\,
            I => \N__5880\
        );

    \I__493\ : Span4Mux_s3_v
    port map (
            O => \N__5880\,
            I => \N__5877\
        );

    \I__492\ : Span4Mux_v
    port map (
            O => \N__5877\,
            I => \N__5874\
        );

    \I__491\ : Odrv4
    port map (
            O => \N__5874\,
            I => \wRamRdData_2\
        );

    \I__490\ : IoInMux
    port map (
            O => \N__5871\,
            I => \N__5868\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__5868\,
            I => \N__5865\
        );

    \I__488\ : Span12Mux_s6_v
    port map (
            O => \N__5865\,
            I => \N__5862\
        );

    \I__487\ : Odrv12
    port map (
            O => \N__5862\,
            I => \wRamRdData_5\
        );

    \IN_MUX_bfv_14_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_2_0_\
        );

    \IN_MUX_bfv_14_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DUT.uart_inst0.tx_clk_divider_cry_7\,
            carryinitout => \bfn_14_3_0_\
        );

    \IN_MUX_bfv_13_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_7_0_\
        );

    \IN_MUX_bfv_13_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DUT.uart_inst0.rx_clk_divider_1_cry_7\,
            carryinitout => \bfn_13_8_0_\
        );

    \IN_MUX_bfv_13_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DUT.uart_inst0.rx_clk_divider_1_cry_15\,
            carryinitout => \bfn_13_9_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_18_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_12_0_\
        );

    \IN_MUX_bfv_15_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_9_0_\
        );

    \top_pll_inst.top_pll_inst_RNISDA2_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5967\,
            GLOBALBUFFEROUTPUT => \wPllLocked_iso_i_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \top_pll_inst.top_pll_inst_RNISDA2\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__10822\,
            GLOBALBUFFEROUTPUT => \wPllLocked_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5973\,
            lcout => \wPllLocked\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.oPacketAvail_latch_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__14548\,
            in1 => \N__14588\,
            in2 => \_gnd_net_\,
            in3 => \N__7809\,
            lcout => \G_120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \top_pll_inst.top_pll_inst_RNISDA2_0_LC_12_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__14574\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \top_pll_inst.wPllLocked_iso_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_0_2_LC_13_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6484\,
            in1 => \N__6459\,
            in2 => \N__6428\,
            in3 => \N__6670\,
            lcout => \DUT.uart_inst0.N_159_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNI92K37_0_LC_13_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__6885\,
            in1 => \N__6057\,
            in2 => \N__8307\,
            in3 => \N__7014\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNINQKO8_1_LC_13_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__10787\,
            in1 => \N__8394\,
            in2 => \N__6024\,
            in3 => \N__6216\,
            lcout => \DUT.uart_inst0.N_22\,
            ltout => \DUT.uart_inst0.N_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_1_LC_13_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6422\,
            in2 => \N__6021\,
            in3 => \N__6464\,
            lcout => \DUT.uart_inst0.tx_bits_remainingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15035\,
            ce => 'H',
            sr => \N__6606\
        );

    \DUT.uart_inst0.tx_bits_remaining_2_LC_13_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101001"
        )
    port map (
            in0 => \N__6485\,
            in1 => \N__6460\,
            in2 => \N__6018\,
            in3 => \N__6426\,
            lcout => \DUT.uart_inst0.tx_bits_remainingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15035\,
            ce => 'H',
            sr => \N__6606\
        );

    \DUT.uart_inst0.tx_bits_remaining_0_LC_13_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6421\,
            in2 => \_gnd_net_\,
            in3 => \N__6014\,
            lcout => \DUT.uart_inst0.tx_bits_remainingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15035\,
            ce => 'H',
            sr => \N__6606\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_2_LC_13_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6483\,
            in1 => \N__6458\,
            in2 => \N__6427\,
            in3 => \N__6669\,
            lcout => \DUT.uart_inst0.N_159\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_RNI2V95_2_LC_13_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6320\,
            in1 => \N__6335\,
            in2 => \N__6354\,
            in3 => \N__6305\,
            lcout => \DUT.uart_inst0.un1_tx_clk_divider_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_13_LC_13_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6521\,
            in1 => \N__6275\,
            in2 => \N__6504\,
            in3 => \N__6290\,
            lcout => \DUT.uart_inst0.un1_tx_clk_divider_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_8_LC_13_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6554\,
            in1 => \N__6245\,
            in2 => \N__6540\,
            in3 => \N__6260\,
            lcout => \DUT.uart_inst0.un1_tx_clk_divider_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNI01HK1_5_LC_13_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__7127\,
            in1 => \N__6846\,
            in2 => \N__7335\,
            in3 => \N__7082\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNIJKPE2_4_LC_13_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__6740\,
            in1 => \_gnd_net_\,
            in2 => \N__6060\,
            in3 => \N__6792\,
            lcout => \DUT.uart_inst0.g2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_1_LC_13_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7128\,
            in1 => \N__6618\,
            in2 => \_gnd_net_\,
            in3 => \N__7363\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15029\,
            ce => \N__14421\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_RNIBPK2_0_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__6372\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8543\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.un1_tx_clk_divider_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_RNITC2S1_0_LC_13_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6051\,
            in1 => \N__6045\,
            in2 => \N__6039\,
            in3 => \N__6036\,
            lcout => \DUT.uart_inst0.un1_tx_clk_divider_0\,
            ltout => \DUT.uart_inst0.un1_tx_clk_divider_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNI3MLP6_0_LC_13_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101110000"
        )
    port map (
            in0 => \N__6695\,
            in1 => \N__6938\,
            in2 => \N__6030\,
            in3 => \N__6881\,
            lcout => \DUT.uart_inst0.N_109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_13_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__7001\,
            in1 => \N__6636\,
            in2 => \N__6093\,
            in3 => \N__8303\,
            lcout => \DUT.uart_inst0.N_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNIMDQK4_0_0_LC_13_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__8302\,
            in1 => \N__6880\,
            in2 => \_gnd_net_\,
            in3 => \N__6998\,
            lcout => \DUT.uart_inst0.N_152\,
            ltout => \DUT.uart_inst0.N_152_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNIBVOQB_1_LC_13_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__7000\,
            in1 => \N__6629\,
            in2 => \N__6027\,
            in3 => \N__6678\,
            lcout => \DUT.uart_inst0.tx_countdown_7_sm0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_3_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__6081\,
            in1 => \N__6438\,
            in2 => \N__6672\,
            in3 => \N__6387\,
            lcout => \DUT.uart_inst0.tx_bits_remainingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15023\,
            ce => 'H',
            sr => \N__6605\
        );

    \DUT.uart_inst0.tx_state_RNISP995_0_LC_13_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6999\,
            in1 => \N__6696\,
            in2 => \N__6939\,
            in3 => \N__6580\,
            lcout => \DUT.uart_inst0.N_120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNIDD8Q_0_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7121\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7071\,
            lcout => \DUT.uart_inst0.tx_countdown_0_ac0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_2_2_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__7072\,
            in1 => \N__6788\,
            in2 => \N__6741\,
            in3 => \N__7122\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_countdown_7_m1_0_o2_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_1_2_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__8273\,
            in1 => \N__7397\,
            in2 => \N__6075\,
            in3 => \N__6630\,
            lcout => \DUT.uart_inst0.N_113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNILLC71_2_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__7070\,
            in1 => \N__7120\,
            in2 => \_gnd_net_\,
            in3 => \N__7321\,
            lcout => \DUT.uart_inst0.tx_countdown_0_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_RNO_1_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__6911\,
            in1 => \N__7797\,
            in2 => \N__8298\,
            in3 => \N__8390\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_out_6_iv_0_a3_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_RNO_0_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111110"
        )
    port map (
            in0 => \N__7734\,
            in1 => \N__6066\,
            in2 => \N__6072\,
            in3 => \N__7141\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_out_6_iv_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__7142\,
            in1 => \N__7768\,
            in2 => \N__6069\,
            in3 => \N__8272\,
            lcout => \P1A7_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15017\,
            ce => \N__14428\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_RNO_3_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010000000100"
        )
    port map (
            in0 => \N__9425\,
            in1 => \N__7758\,
            in2 => \N__8297\,
            in3 => \N__6910\,
            lcout => \DUT.uart_inst0.N_119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_0_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000100010"
        )
    port map (
            in0 => \N__6959\,
            in1 => \N__7069\,
            in2 => \_gnd_net_\,
            in3 => \N__7364\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15012\,
            ce => \N__14435\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_0_4_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100100000000"
        )
    port map (
            in0 => \N__6784\,
            in1 => \N__6732\,
            in2 => \N__6810\,
            in3 => \N__6958\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_countdown_RNO_0Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_4_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__6733\,
            in1 => \_gnd_net_\,
            in2 => \N__6102\,
            in3 => \N__7365\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15012\,
            ce => \N__14435\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNI34HK1_5_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6837\,
            in1 => \N__6730\,
            in2 => \N__7081\,
            in3 => \N__7319\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNIJKPE2_1_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6780\,
            in2 => \N__6099\,
            in3 => \N__7123\,
            lcout => \DUT.uart_inst0.N_100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNO_5_3_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6838\,
            in1 => \N__7320\,
            in2 => \N__6791\,
            in3 => \N__6731\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.m25_e_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNO_3_3_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001001100"
        )
    port map (
            in0 => \N__7076\,
            in1 => \N__6671\,
            in2 => \N__6096\,
            in3 => \N__7124\,
            lcout => \DUT.uart_inst0.m3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_5_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101001000000"
        )
    port map (
            in0 => \N__7366\,
            in1 => \N__6960\,
            in2 => \N__7401\,
            in3 => \N__6842\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15012\,
            ce => \N__14435\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8136\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_7_0_\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8106\,
            in2 => \N__9180\,
            in3 => \N__6129\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_0\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8079\,
            in2 => \N__9188\,
            in3 => \N__6126\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_1\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNO_0_3_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8052\,
            in2 => \N__9182\,
            in3 => \N__6123\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_3\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_2\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8463\,
            in2 => \N__9189\,
            in3 => \N__6120\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_3\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNO_0_5_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7488\,
            in2 => \N__9183\,
            in3 => \N__6117\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_5\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_4\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNO_0_6_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7470\,
            in2 => \N__9190\,
            in3 => \N__6114\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_6\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_5\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7511\,
            in2 => \N__9181\,
            in3 => \N__6111\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_6\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7451\,
            in2 => \N__9186\,
            in3 => \N__6108\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_13_8_0_\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7161\,
            in2 => \N__9194\,
            in3 => \N__6105\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_8\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_LUT4_0_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7185\,
            in2 => \N__9187\,
            in3 => \N__6153\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_9\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_LUT4_0_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7538\,
            in2 => \N__9191\,
            in3 => \N__6150\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_10\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_LUT4_0_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7426\,
            in2 => \N__9184\,
            in3 => \N__6147\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_11\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_LUT4_0_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7259\,
            in2 => \N__9192\,
            in3 => \N__6144\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_12\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_LUT4_0_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7232\,
            in2 => \N__9185\,
            in3 => \N__6141\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_13\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_LUT4_0_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7209\,
            in2 => \N__9193\,
            in3 => \N__6138\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_14\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_LUT4_0_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8156\,
            in2 => \N__9195\,
            in3 => \N__6135\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_13_9_0_\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_17_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000000001011"
        )
    port map (
            in0 => \N__10518\,
            in1 => \N__11013\,
            in2 => \N__7286\,
            in3 => \N__6132\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15000\,
            ce => \N__14450\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6195\,
            in2 => \N__9469\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_10_0_\,
            carryout => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_1_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6204\,
            in2 => \N__9511\,
            in3 => \N__6210\,
            lcout => \DUT.fifo_tx_inst.rFifoCountZ0Z_1\,
            ltout => OPEN,
            carryin => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0\,
            carryout => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1\,
            clk => \N__14997\,
            ce => 'H',
            sr => \N__15219\
        );

    \DUT.fifo_tx_inst.rFifoCount_2_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110001110011100"
        )
    port map (
            in0 => \N__6189\,
            in1 => \N__9325\,
            in2 => \N__9434\,
            in3 => \N__6207\,
            lcout => \DUT.fifo_tx_inst.rFifoCountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14997\,
            ce => 'H',
            sr => \N__15219\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNISSQ21_1_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \N__9496\,
            in1 => \N__9430\,
            in2 => \_gnd_net_\,
            in3 => \N__6187\,
            lcout => \DUT.fifo_tx_inst.rFifoCount_RNISSQ21Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNI0AJL_0_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__9318\,
            in1 => \N__9495\,
            in2 => \N__6173\,
            in3 => \N__9455\,
            lcout => \DUT.fifo_tx_inst.N_108\,
            ltout => \DUT.fifo_tx_inst.N_108_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000111111"
        )
    port map (
            in0 => \N__9457\,
            in1 => \N__9429\,
            in2 => \N__6198\,
            in3 => \N__12238\,
            lcout => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_2_1_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__9319\,
            in1 => \N__12311\,
            in2 => \N__6174\,
            in3 => \N__12263\,
            lcout => \DUT.fifo_tx_inst.rFifoData_awe3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_0_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001101010010101"
        )
    port map (
            in0 => \N__9456\,
            in1 => \N__6188\,
            in2 => \N__9435\,
            in3 => \N__12239\,
            lcout => \DUT.fifo_tx_inst.rFifoCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14995\,
            ce => 'H',
            sr => \N__15218\
        );

    \rTxWrite_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14824\,
            in2 => \_gnd_net_\,
            in3 => \N__12549\,
            lcout => \rTxWriteZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14995\,
            ce => 'H',
            sr => \N__15218\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNI7FOF_2_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6166\,
            in2 => \_gnd_net_\,
            in3 => \N__9317\,
            lcout => \DUT.fifo_tx_inst.N_104\,
            ltout => \DUT.fifo_tx_inst.N_104_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_0_1_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12312\,
            in2 => \N__6156\,
            in3 => \N__12264\,
            lcout => \DUT.fifo_tx_inst.rFifoData_awe1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110001101"
        )
    port map (
            in0 => \N__10708\,
            in1 => \N__10170\,
            in2 => \N__9210\,
            in3 => \N__10296\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.rx_countdown_8_i_o2_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_2_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001110"
        )
    port map (
            in0 => \N__7617\,
            in1 => \N__6231\,
            in2 => \N__6234\,
            in3 => \N__8907\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14994\,
            ce => \N__14460\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_5_2_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__11568\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11117\,
            lcout => \DUT.uart_inst0.m4_e_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_2_2_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000100000"
        )
    port map (
            in0 => \N__11119\,
            in1 => \N__10707\,
            in2 => \N__10851\,
            in3 => \N__10001\,
            lcout => \DUT.uart_inst0.N_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNIUMLT1_5_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11489\,
            in1 => \N__11245\,
            in2 => \N__11574\,
            in3 => \N__11118\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g0_0_0_a3_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNI7CGS2_1_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11400\,
            in2 => \N__6225\,
            in3 => \N__10101\,
            lcout => \DUT.uart_inst0.g0_0_0_a3_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_3_1_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11488\,
            in1 => \N__11244\,
            in2 => \N__11573\,
            in3 => \N__11116\,
            lcout => \DUT.uart_inst0.N_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNIBTN81_0_LC_14_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100010001"
        )
    port map (
            in0 => \N__9416\,
            in1 => \N__8300\,
            in2 => \_gnd_net_\,
            in3 => \N__6222\,
            lcout => \DUT.uart_inst0.N_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_14_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8547\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_2_0_\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_1_LC_14_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6371\,
            in2 => \N__9054\,
            in3 => \N__6357\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_1\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_0\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_1\,
            clk => \N__15043\,
            ce => 'H',
            sr => \N__8514\
        );

    \DUT.uart_inst0.tx_clk_divider_2_LC_14_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6353\,
            in2 => \N__9058\,
            in3 => \N__6339\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_2\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_1\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_2\,
            clk => \N__15043\,
            ce => 'H',
            sr => \N__8514\
        );

    \DUT.uart_inst0.tx_clk_divider_3_LC_14_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6336\,
            in2 => \N__9055\,
            in3 => \N__6324\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_3\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_2\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_3\,
            clk => \N__15043\,
            ce => 'H',
            sr => \N__8514\
        );

    \DUT.uart_inst0.tx_clk_divider_4_LC_14_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6321\,
            in2 => \N__9059\,
            in3 => \N__6309\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_4\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_3\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_4\,
            clk => \N__15043\,
            ce => 'H',
            sr => \N__8514\
        );

    \DUT.uart_inst0.tx_clk_divider_5_LC_14_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6306\,
            in2 => \N__9056\,
            in3 => \N__6294\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_5\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_4\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_5\,
            clk => \N__15043\,
            ce => 'H',
            sr => \N__8514\
        );

    \DUT.uart_inst0.tx_clk_divider_6_LC_14_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6291\,
            in2 => \N__9060\,
            in3 => \N__6279\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_6\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_5\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_6\,
            clk => \N__15043\,
            ce => 'H',
            sr => \N__8514\
        );

    \DUT.uart_inst0.tx_clk_divider_7_LC_14_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6276\,
            in2 => \N__9057\,
            in3 => \N__6264\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_7\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_6\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_7\,
            clk => \N__15043\,
            ce => 'H',
            sr => \N__8514\
        );

    \DUT.uart_inst0.tx_clk_divider_8_LC_14_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6261\,
            in2 => \N__9126\,
            in3 => \N__6249\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_14_3_0_\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_8\,
            clk => \N__15036\,
            ce => 'H',
            sr => \N__8509\
        );

    \DUT.uart_inst0.tx_clk_divider_9_LC_14_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6246\,
            in2 => \N__9128\,
            in3 => \N__6558\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_9\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_8\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_9\,
            clk => \N__15036\,
            ce => 'H',
            sr => \N__8509\
        );

    \DUT.uart_inst0.tx_clk_divider_10_LC_14_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6555\,
            in2 => \N__9124\,
            in3 => \N__6543\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_10\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_9\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_10\,
            clk => \N__15036\,
            ce => 'H',
            sr => \N__8509\
        );

    \DUT.uart_inst0.tx_clk_divider_11_LC_14_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6539\,
            in2 => \N__9127\,
            in3 => \N__6525\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_11\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_10\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_11\,
            clk => \N__15036\,
            ce => 'H',
            sr => \N__8509\
        );

    \DUT.uart_inst0.tx_clk_divider_12_LC_14_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6522\,
            in2 => \N__9125\,
            in3 => \N__6510\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_12\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_11\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_12\,
            clk => \N__15036\,
            ce => 'H',
            sr => \N__8509\
        );

    \DUT.uart_inst0.tx_clk_divider_13_LC_14_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6503\,
            in2 => \_gnd_net_\,
            in3 => \N__6507\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15036\,
            ce => 'H',
            sr => \N__8509\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNO_1_3_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__6489\,
            in1 => \N__6393\,
            in2 => \N__8386\,
            in3 => \N__6468\,
            lcout => \DUT.uart_inst0.m9_e_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNO_4_3_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__14547\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6429\,
            lcout => \DUT.uart_inst0.m9_e_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNIMDQK4_0_LC_14_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__6694\,
            in1 => \N__7008\,
            in2 => \N__8301\,
            in3 => \N__6934\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_state_0_sqmuxa_i_i_a3_c_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNI00K8B_0_LC_14_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6386\,
            in1 => \N__7947\,
            in2 => \N__6375\,
            in3 => \N__6584\,
            lcout => \DUT.uart_inst0.N_22_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNICODU_0_LC_14_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8279\,
            in2 => \_gnd_net_\,
            in3 => \N__6908\,
            lcout => \DUT.uart_inst0.N_160\,
            ltout => \DUT.uart_inst0.N_160_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNI6Q5N3_1_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__6933\,
            in1 => \N__8365\,
            in2 => \N__6699\,
            in3 => \N__6693\,
            lcout => \DUT.uart_inst0.N_154\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNO_2_3_LC_14_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__9398\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6665\,
            lcout => \DUT.uart_inst0.N_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNIIAMI1_1_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011101111"
        )
    port map (
            in0 => \N__6909\,
            in1 => \N__8364\,
            in2 => \N__8299\,
            in3 => \N__9399\,
            lcout => \DUT.uart_inst0.N_99\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNI5PJS2_1_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__7959\,
            in1 => \N__14549\,
            in2 => \_gnd_net_\,
            in3 => \N__7012\,
            lcout => \DUT.uart_inst0.N_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_0_1_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000001000"
        )
    port map (
            in0 => \N__7010\,
            in1 => \N__7957\,
            in2 => \N__7083\,
            in3 => \N__7125\,
            lcout => \DUT.uart_inst0.tx_countdown_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNI8CH01_0_1_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7958\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14550\,
            lcout => \DUT.uart_inst0.N_88_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_0_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001110"
        )
    port map (
            in0 => \N__8277\,
            in1 => \N__9397\,
            in2 => \N__8393\,
            in3 => \N__6564\,
            lcout => \DUT.tx_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15024\,
            ce => 'H',
            sr => \N__15229\
        );

    \DUT.uart_inst0.tx_state_RNIOJJIA_0_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__6879\,
            in1 => \N__7028\,
            in2 => \N__6585\,
            in3 => \N__7011\,
            lcout => \DUT.uart_inst0.N_218\,
            ltout => \DUT.uart_inst0.N_218_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_1_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8382\,
            in2 => \N__7146\,
            in3 => \N__7143\,
            lcout => \DUT.tx_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15024\,
            ce => 'H',
            sr => \N__15229\
        );

    \DUT.uart_inst0.tx_countdown_RNO_0_2_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111000000000"
        )
    port map (
            in0 => \N__7126\,
            in1 => \N__7080\,
            in2 => \N__7331\,
            in3 => \N__7009\,
            lcout => \DUT.uart_inst0.tx_countdown_7_m1_0_a3_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__6779\,
            in1 => \N__6852\,
            in2 => \_gnd_net_\,
            in3 => \N__7032\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_countdown_RNO_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_3_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6945\,
            in2 => \N__7017\,
            in3 => \N__7367\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15018\,
            ce => \N__14436\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNI9B9Q2_1_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110100000000"
        )
    port map (
            in0 => \N__9408\,
            in1 => \N__8267\,
            in2 => \N__8391\,
            in3 => \N__7013\,
            lcout => \DUT.uart_inst0.N_164\,
            ltout => \DUT.uart_inst0.N_164_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000001010000"
        )
    port map (
            in0 => \N__6806\,
            in1 => \_gnd_net_\,
            in2 => \N__6948\,
            in3 => \N__6778\,
            lcout => \DUT.uart_inst0.tx_countdown_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNI67HK1_5_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6835\,
            in1 => \N__7317\,
            in2 => \N__6789\,
            in3 => \N__6728\,
            lcout => \DUT.uart_inst0.tx_state_ns_i_i_o2_a0_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_2_3_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__8268\,
            in1 => \N__6915\,
            in2 => \N__8392\,
            in3 => \N__6878\,
            lcout => \DUT.uart_inst0.N_163\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNIJKPE2_5_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101001"
        )
    port map (
            in0 => \N__6836\,
            in1 => \N__6805\,
            in2 => \N__6790\,
            in3 => \N__6729\,
            lcout => \DUT.uart_inst0.tx_countdown_30_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_2_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000111111"
        )
    port map (
            in0 => \N__7318\,
            in1 => \N__7386\,
            in2 => \N__7377\,
            in3 => \N__7368\,
            lcout => \DUT.uart_inst0.N_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15018\,
            ce => \N__14436\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNI3ALC_17_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7207\,
            in1 => \N__7231\,
            in2 => \N__7287\,
            in3 => \N__7258\,
            lcout => \DUT.uart_inst0.un2_rx_clk_divider_a_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_13_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110000100011"
        )
    port map (
            in0 => \N__10504\,
            in1 => \N__7260\,
            in2 => \N__11016\,
            in3 => \N__7266\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15013\,
            ce => \N__14443\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_14_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001101000001"
        )
    port map (
            in0 => \N__11012\,
            in1 => \N__7242\,
            in2 => \N__7236\,
            in3 => \N__10505\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15013\,
            ce => \N__14443\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_15_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010000110001"
        )
    port map (
            in0 => \N__11005\,
            in1 => \N__7215\,
            in2 => \N__10557\,
            in3 => \N__7208\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15013\,
            ce => \N__14443\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_10_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000010010100101"
        )
    port map (
            in0 => \N__7184\,
            in1 => \N__10502\,
            in2 => \N__7194\,
            in3 => \N__11009\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15013\,
            ce => \N__14443\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIB99J_10_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7537\,
            in1 => \N__7183\,
            in2 => \N__7428\,
            in3 => \N__7159\,
            lcout => \DUT.uart_inst0.un2_rx_clk_divider_a_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_9_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000010010100101"
        )
    port map (
            in0 => \N__7160\,
            in1 => \N__10509\,
            in2 => \N__7170\,
            in3 => \N__11010\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15013\,
            ce => \N__14443\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_11_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000001011000011"
        )
    port map (
            in0 => \N__10503\,
            in1 => \N__7539\,
            in2 => \N__7548\,
            in3 => \N__11011\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15013\,
            ce => \N__14443\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNI6B671_5_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7510\,
            in1 => \N__7469\,
            in2 => \N__7452\,
            in3 => \N__7487\,
            lcout => \DUT.uart_inst0.un2_rx_clk_divider_a_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_7_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001101000001"
        )
    port map (
            in0 => \N__10995\,
            in1 => \N__7521\,
            in2 => \N__7515\,
            in3 => \N__10535\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15007\,
            ce => \N__14451\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_5_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__7494\,
            in1 => \N__10996\,
            in2 => \N__10562\,
            in3 => \N__10683\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15007\,
            ce => \N__14451\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_6_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__10682\,
            in1 => \N__10531\,
            in2 => \N__11014\,
            in3 => \N__7476\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15007\,
            ce => \N__14451\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_8_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001001010001"
        )
    port map (
            in0 => \N__7450\,
            in1 => \N__10997\,
            in2 => \N__10563\,
            in3 => \N__7458\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15007\,
            ce => \N__14451\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_12_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101001000101"
        )
    port map (
            in0 => \N__7434\,
            in1 => \N__10526\,
            in2 => \N__11015\,
            in3 => \N__7427\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15007\,
            ce => \N__14451\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_16_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000001011000011"
        )
    port map (
            in0 => \N__10527\,
            in1 => \N__7407\,
            in2 => \N__8163\,
            in3 => \N__11004\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15007\,
            ce => \N__14451\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011101"
        )
    port map (
            in0 => \N__10994\,
            in1 => \N__10536\,
            in2 => \_gnd_net_\,
            in3 => \N__7575\,
            lcout => \DUT.uart_inst0.rx_countdownZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15007\,
            ce => \N__14451\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_6_2_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10276\,
            in2 => \_gnd_net_\,
            in3 => \N__10157\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.m7_e_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_3_2_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__9909\,
            in1 => \N__9984\,
            in2 => \N__7590\,
            in3 => \N__10218\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.m7_e_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_2_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111011101"
        )
    port map (
            in0 => \N__7554\,
            in1 => \N__10677\,
            in2 => \N__7587\,
            in3 => \N__10099\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.m9_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_2_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000010001010"
        )
    port map (
            in0 => \N__10812\,
            in1 => \N__8799\,
            in2 => \N__7584\,
            in3 => \N__7581\,
            lcout => \DUT_uart_inst0_recv_state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15003\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_1_2_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011110011"
        )
    port map (
            in0 => \N__8619\,
            in1 => \N__8874\,
            in2 => \N__10482\,
            in3 => \N__8798\,
            lcout => \DUT.uart_inst0.N_11_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_3_1_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10275\,
            in1 => \N__9983\,
            in2 => \N__10168\,
            in3 => \N__10217\,
            lcout => \DUT.uart_inst0.g1_i_a4_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_0_3_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001101"
        )
    port map (
            in0 => \N__11220\,
            in1 => \N__10676\,
            in2 => \N__10890\,
            in3 => \N__10158\,
            lcout => \DUT.uart_inst0.N_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_2_2_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__11498\,
            in1 => \N__11219\,
            in2 => \N__7569\,
            in3 => \N__11399\,
            lcout => \DUT.uart_inst0.m4_e_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_0_1_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__7623\,
            in1 => \N__10695\,
            in2 => \_gnd_net_\,
            in3 => \N__7653\,
            lcout => \DUT.uart_inst0.N_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNI9JOT_0_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8637\,
            in2 => \N__8688\,
            in3 => \N__8783\,
            lcout => \DUT.uart_inst0.m5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_4_1_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10271\,
            in1 => \N__10142\,
            in2 => \N__9995\,
            in3 => \N__10216\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_21_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_2_1_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111110101"
        )
    port map (
            in0 => \N__8677\,
            in1 => \_gnd_net_\,
            in2 => \N__7656\,
            in3 => \N__7641\,
            lcout => \DUT.uart_inst0.N_21_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNIO2V22_1_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110011"
        )
    port map (
            in0 => \N__8784\,
            in1 => \N__8863\,
            in2 => \N__10567\,
            in3 => \N__7647\,
            lcout => \DUT.uart_inst0.N_6\,
            ltout => \DUT.uart_inst0.N_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_1_1_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__8676\,
            in1 => \_gnd_net_\,
            in2 => \N__7635\,
            in3 => \N__7632\,
            lcout => \DUT.uart_inst0.N_18_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_0_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__8638\,
            in1 => \N__8865\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.uart_inst0.rx_bits_remainingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15001\,
            ce => \N__8826\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__8864\,
            in1 => \N__10547\,
            in2 => \_gnd_net_\,
            in3 => \N__8785\,
            lcout => \DUT.uart_inst0.N_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_1_1_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__11040\,
            in1 => \N__10093\,
            in2 => \N__7605\,
            in3 => \N__9926\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g1_i_a4_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_1_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001000100"
        )
    port map (
            in0 => \N__9819\,
            in1 => \N__8577\,
            in2 => \N__7593\,
            in3 => \N__10702\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14998\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNIS6O94_0_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__7677\,
            in1 => \N__10291\,
            in2 => \_gnd_net_\,
            in3 => \N__10229\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g0_0_0_a3_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNIL139C_1_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__7686\,
            in1 => \N__7713\,
            in2 => \N__7680\,
            in3 => \N__10701\,
            lcout => \DUT.uart_inst0.recv_state_RNIL139CZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_3_6_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10164\,
            in1 => \N__9925\,
            in2 => \N__10002\,
            in3 => \N__10290\,
            lcout => \DUT.uart_inst0.m13_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNI69LM2_0_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__9997\,
            in1 => \N__9913\,
            in2 => \N__10100\,
            in3 => \N__10163\,
            lcout => \DUT.uart_inst0.g0_0_0_a3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_RNI4PUO_1_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__14561\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12659\,
            lcout => \DUT.fifo_tx_inst.un1_i11_i\,
            ltout => \DUT.fifo_tx_inst.un1_i11_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_1_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000000110"
        )
    port map (
            in0 => \N__12315\,
            in1 => \N__12271\,
            in2 => \N__7671\,
            in3 => \N__12240\,
            lcout => \DUT.fifo_tx_inst.rWritePtrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14998\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_0_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__12369\,
            in1 => \N__12179\,
            in2 => \_gnd_net_\,
            in3 => \N__7664\,
            lcout => \DUT.fifo_rx_inst.rWritePtrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14996\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_1_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101000000"
        )
    port map (
            in0 => \N__7665\,
            in1 => \N__12370\,
            in2 => \N__12183\,
            in3 => \N__12329\,
            lcout => \DUT.fifo_rx_inst.rWritePtrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14996\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNI96D91_2_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__12328\,
            in1 => \N__12592\,
            in2 => \N__12374\,
            in3 => \N__13902\,
            lcout => \DUT.fifo_rx_inst.N_57\,
            ltout => \DUT.fifo_rx_inst.N_57_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNI5KNB1_2_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7668\,
            in3 => \N__14562\,
            lcout => \DUT.fifo_rx_inst.un1_i11_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_2_6_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__10230\,
            in1 => \N__10791\,
            in2 => \N__10568\,
            in3 => \N__11337\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.m13_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_6_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__10578\,
            in1 => \N__10097\,
            in2 => \N__7725\,
            in3 => \N__7722\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.P19_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_6_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010010000"
        )
    port map (
            in0 => \N__10098\,
            in1 => \N__10710\,
            in2 => \N__7716\,
            in3 => \N__9927\,
            lcout => \DUT.wRcvd\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14996\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNIBTG71_1_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010000000000"
        )
    port map (
            in0 => \N__10548\,
            in1 => \N__8869\,
            in2 => \N__8808\,
            in3 => \N__14563\,
            lcout => \DUT.uart_inst0.g0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ioFifoData_iobuf_RNO_0_LC_15_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13836\,
            lcout => \N_1257_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.oTxFull_0_LC_15_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7845\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7898\,
            lcout => \fifo_inst_ftdi_input_inst_oTxFull_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.rPacketCount_latch_1_LC_15_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100100000"
        )
    port map (
            in0 => \N__7925\,
            in1 => \N__15285\,
            in2 => \N__7880\,
            in3 => \N__7846\,
            lcout => \G_111\,
            ltout => \G_111_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.SUM_2_LC_15_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__7827\,
            in1 => \_gnd_net_\,
            in2 => \N__7692\,
            in3 => \N__7868\,
            lcout => OPEN,
            ltout => \fifo_inst.ftdi_input_inst.SUMZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.rPacketCount_latch_2_LC_15_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__7926\,
            in1 => \N__7828\,
            in2 => \N__7689\,
            in3 => \N__15286\,
            lcout => \G_112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.rPacketCount_latch_3_LC_15_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__7924\,
            in1 => \N__7908\,
            in2 => \N__15291\,
            in3 => \N__7900\,
            lcout => \G_109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.rPacketCount_latch_0_LC_15_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15284\,
            in2 => \N__7879\,
            in3 => \N__7923\,
            lcout => \G_110\,
            ltout => \G_110_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.wTxEn_1_LC_15_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011001100"
        )
    port map (
            in0 => \N__7826\,
            in1 => \N__14546\,
            in2 => \N__7935\,
            in3 => \N__7932\,
            lcout => \G_114\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.rPacketCount15_LC_15_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7899\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9570\,
            lcout => \G_108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.SUM_3_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__7829\,
            in1 => \N__7847\,
            in2 => \N__7881\,
            in3 => \N__7901\,
            lcout => \fifo_inst.ftdi_input_inst.SUMZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.un2_oPacketAvail_i_LC_15_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__7902\,
            in1 => \N__7878\,
            in2 => \N__7851\,
            in3 => \N__7830\,
            lcout => \fifo_inst.ftdi_input_inst.un2_oPacketAvail_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_7_LC_15_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000101010"
        )
    port map (
            in0 => \N__8940\,
            in1 => \N__9609\,
            in2 => \N__9624\,
            in3 => \N__8278\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15037\,
            ce => \N__7970\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_0_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__8260\,
            in1 => \N__9273\,
            in2 => \N__8037\,
            in3 => \N__9588\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15030\,
            ce => \N__7971\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_RNO_2_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011000000"
        )
    port map (
            in0 => \N__7790\,
            in1 => \N__8369\,
            in2 => \N__7778\,
            in3 => \N__8259\,
            lcout => \DUT.uart_inst0.N_116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_1_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__8261\,
            in1 => \N__9249\,
            in2 => \N__8028\,
            in3 => \N__9589\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15030\,
            ce => \N__7971\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_2_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__9590\,
            in1 => \N__11760\,
            in2 => \N__8019\,
            in3 => \N__8264\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15030\,
            ce => \N__7971\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_3_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__8262\,
            in1 => \N__11589\,
            in2 => \N__8007\,
            in3 => \N__9591\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15030\,
            ce => \N__7971\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_4_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__9592\,
            in1 => \N__9240\,
            in2 => \N__7998\,
            in3 => \N__8265\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15030\,
            ce => \N__7971\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_5_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__8263\,
            in1 => \N__9543\,
            in2 => \N__7980\,
            in3 => \N__9593\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15030\,
            ce => \N__7971\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_6_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__9594\,
            in1 => \N__9519\,
            in2 => \N__7989\,
            in3 => \N__8266\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15030\,
            ce => \N__7971\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNICU6U_1_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__8361\,
            in1 => \N__9372\,
            in2 => \_gnd_net_\,
            in3 => \N__8250\,
            lcout => \DUT.uart_inst0.N_102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.rWrState_latch_1_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9754\,
            in1 => \N__14552\,
            in2 => \_gnd_net_\,
            in3 => \N__9730\,
            lcout => \G_113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNI8CH01_1_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110111111"
        )
    port map (
            in0 => \N__8362\,
            in1 => \N__9373\,
            in2 => \N__14575\,
            in3 => \N__8251\,
            lcout => \DUT.uart_inst0.tx_state_0_sqmuxa_i_i_a3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNIN9O8_0_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__9513\,
            in1 => \N__9477\,
            in2 => \_gnd_net_\,
            in3 => \N__9333\,
            lcout => OPEN,
            ltout => \DUT.N_114_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.rTransmit_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8363\,
            in1 => \N__14551\,
            in2 => \N__8310\,
            in3 => \N__8252\,
            lcout => \DUT.rTransmitZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15025\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_0_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110110011"
        )
    port map (
            in0 => \N__10953\,
            in1 => \N__14557\,
            in2 => \N__10558\,
            in3 => \N__12608\,
            lcout => \DUT.uart_inst0.G_19_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIMQ571_1_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8048\,
            in1 => \N__8074\,
            in2 => \N__8462\,
            in3 => \N__8101\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.un2_rx_clk_divider_a_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIJI4K1_16_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8155\,
            in2 => \N__8139\,
            in3 => \N__8128\,
            lcout => \DUT.uart_inst0.un2_rx_clk_divider_a_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_0_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__8129\,
            in1 => \N__10513\,
            in2 => \_gnd_net_\,
            in3 => \N__10959\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15019\,
            ce => \N__14452\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101001000101"
        )
    port map (
            in0 => \N__8102\,
            in1 => \N__10519\,
            in2 => \N__10993\,
            in3 => \N__8115\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15019\,
            ce => \N__14452\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_2_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001001010001"
        )
    port map (
            in0 => \N__8088\,
            in1 => \N__10955\,
            in2 => \N__10560\,
            in3 => \N__8075\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15019\,
            ce => \N__14452\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_3_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__10954\,
            in1 => \N__8061\,
            in2 => \N__10559\,
            in3 => \N__10686\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15019\,
            ce => \N__14452\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_4_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001000010011001"
        )
    port map (
            in0 => \N__8458\,
            in1 => \N__8475\,
            in2 => \N__10561\,
            in3 => \N__10960\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15019\,
            ce => \N__14452\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNINK4E1_2_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__8787\,
            in1 => \N__11455\,
            in2 => \N__14576\,
            in3 => \N__11218\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.m6_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNI3V794_0_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010110111111"
        )
    port map (
            in0 => \N__10057\,
            in1 => \N__9771\,
            in2 => \N__8442\,
            in3 => \N__9903\,
            lcout => \DUT.uart_inst0.G_30_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \top_pll_inst.top_pll_inst_RNIIIF42_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__8788\,
            in1 => \N__10824\,
            in2 => \N__9921\,
            in3 => \N__9982\,
            lcout => OPEN,
            ltout => \top_pll_inst.m12_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \top_pll_inst.top_pll_inst_RNI0MK94_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__10159\,
            in1 => \N__10277\,
            in2 => \N__8439\,
            in3 => \N__10219\,
            lcout => OPEN,
            ltout => \P18_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNIEGJTC_0_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000110001"
        )
    port map (
            in0 => \N__10065\,
            in1 => \N__8436\,
            in2 => \N__8430\,
            in3 => \N__10675\,
            lcout => \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNI7H9R3_10_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8427\,
            in1 => \N__8418\,
            in2 => \N__8412\,
            in3 => \N__8403\,
            lcout => \DUT.uart_inst0.un2_rx_clk_divider_0\,
            ltout => \DUT.uart_inst0.un2_rx_clk_divider_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNI15HA8_0_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001101111011"
        )
    port map (
            in0 => \N__10064\,
            in1 => \N__9792\,
            in2 => \N__8397\,
            in3 => \N__9919\,
            lcout => \DUT.uart_inst0.rx_countdown_8_i_o2_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_4_3_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__11149\,
            in1 => \N__10049\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.uart_inst0.m6_e_2\,
            ltout => OPEN,
            carryin => \bfn_15_9_0_\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_0_s1_c_RNIKPDT_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9113\,
            in2 => \N__11393\,
            in3 => \N__8562\,
            lcout => \DUT_uart_inst0_rx_countdown_3_s1_1\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_countdown_3_cry_0_s1\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNIMVNN_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9177\,
            in2 => \N__11156\,
            in3 => \N__8559\,
            lcout => \DUT_uart_inst0_rx_countdown_3_s1_2\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_countdown_3_cry_1_s1\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_2_s1_c_RNIO52I_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9114\,
            in2 => \N__11224\,
            in3 => \N__8556\,
            lcout => \DUT_uart_inst0_rx_countdown_3_s1_3\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_countdown_3_cry_2_s1\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_3_s1_c_RNIQBCS_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9178\,
            in2 => \N__11467\,
            in3 => \N__8553\,
            lcout => \DUT_uart_inst0_rx_countdown_3_s1_4\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_countdown_3_cry_3_s1\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_4_s1_c_RNISHMM_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11544\,
            in2 => \_gnd_net_\,
            in3 => \N__8550\,
            lcout => \DUT_uart_inst0_rx_countdown_3_s1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_0_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__9115\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8536\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15008\,
            ce => 'H',
            sr => \N__8513\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNIP8561_0_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111000001111"
        )
    port map (
            in0 => \N__8678\,
            in1 => \N__8639\,
            in2 => \N__8739\,
            in3 => \N__8786\,
            lcout => \DUT.uart_inst0.m6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_1_2_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__9225\,
            in1 => \N__8729\,
            in2 => \_gnd_net_\,
            in3 => \N__8921\,
            lcout => \DUT.uart_inst0.N_19_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_4_2_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10292\,
            in1 => \N__10228\,
            in2 => \N__10169\,
            in3 => \N__9985\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_2_2_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8730\,
            in2 => \N__8607\,
            in3 => \N__8922\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_21_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_0_2_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__10699\,
            in1 => \_gnd_net_\,
            in2 => \N__8604\,
            in3 => \N__8601\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_2_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001001110"
        )
    port map (
            in0 => \N__10814\,
            in1 => \N__8731\,
            in2 => \N__8595\,
            in3 => \N__10314\,
            lcout => \DUT.uart_inst0.rx_bits_remainingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15004\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNI40IN5_1_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111111100"
        )
    port map (
            in0 => \N__9908\,
            in1 => \N__11392\,
            in2 => \N__10709\,
            in3 => \N__10081\,
            lcout => \DUT.uart_inst0.rx_countdown_8_i_o2_2_0_2\,
            ltout => \DUT.uart_inst0.rx_countdown_8_i_o2_2_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_1_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100000010"
        )
    port map (
            in0 => \N__10813\,
            in1 => \N__8592\,
            in2 => \N__8586\,
            in3 => \N__8679\,
            lcout => \DUT.uart_inst0.rx_bits_remainingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15004\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_5_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__8568\,
            in1 => \N__8905\,
            in2 => \N__10823\,
            in3 => \N__8913\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15002\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_0_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__12314\,
            in1 => \N__12243\,
            in2 => \_gnd_net_\,
            in3 => \N__8583\,
            lcout => \DUT.fifo_tx_inst.rWritePtrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15002\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_1_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__8867\,
            in1 => \N__14564\,
            in2 => \_gnd_net_\,
            in3 => \N__11035\,
            lcout => \DUT.uart_inst0.g0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_5_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11332\,
            in1 => \N__10555\,
            in2 => \_gnd_net_\,
            in3 => \N__8868\,
            lcout => \DUT.uart_inst0.N_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNI8OBB2_1_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110001"
        )
    port map (
            in0 => \N__8866\,
            in1 => \N__8928\,
            in2 => \N__10569\,
            in3 => \N__8800\,
            lcout => \DUT.uart_inst0.N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNI4AOF7_3_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111110101"
        )
    port map (
            in0 => \N__9216\,
            in1 => \N__10302\,
            in2 => \N__11265\,
            in3 => \N__10700\,
            lcout => \DUT.uart_inst0.recv_state_srsts_1_5\,
            ltout => \DUT.uart_inst0.recv_state_srsts_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_4_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__10879\,
            in1 => \N__8906\,
            in2 => \N__8883\,
            in3 => \N__8880\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15002\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_4_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__14565\,
            in1 => \N__11175\,
            in2 => \_gnd_net_\,
            in3 => \N__10878\,
            lcout => \DUT.uart_inst0.recv_state_srsts_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_0_3_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8693\,
            in2 => \_gnd_net_\,
            in3 => \N__8649\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_43_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_3_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011101011"
        )
    port map (
            in0 => \N__8873\,
            in1 => \N__8709\,
            in2 => \N__8829\,
            in3 => \N__8742\,
            lcout => \DUT.uart_inst0.rx_bits_remainingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__14999\,
            ce => \N__8825\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNIV9PG_3_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8707\,
            in2 => \_gnd_net_\,
            in3 => \N__8647\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.m3_e_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNIAVHE1_2_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__8692\,
            in1 => \N__8741\,
            in2 => \N__8811\,
            in3 => \N__8801\,
            lcout => \DUT.uart_inst0.N_15_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_4_2_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__8740\,
            in1 => \N__8708\,
            in2 => \N__8694\,
            in3 => \N__8648\,
            lcout => \DUT.uart_inst0.recv_state_RNO_4Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_3_2_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11490\,
            in1 => \N__11261\,
            in2 => \N__11572\,
            in3 => \N__11139\,
            lcout => \DUT.uart_inst0.N_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNIEQQU_2_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__11140\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11491\,
            lcout => \DUT.uart_inst0.G_8_i_a3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_3_2_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__11492\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11262\,
            lcout => \DUT.uart_inst0.rx_countdown_8_i_o2_1_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_16_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_16_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12903\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15049\,
            ce => \N__11853\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_16_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13116\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15049\,
            ce => \N__11853\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_16_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__11744\,
            in1 => \N__11781\,
            in2 => \N__11678\,
            in3 => \N__8934\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_16_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__12690\,
            in1 => \N__11865\,
            in2 => \N__8943\,
            in3 => \N__11674\,
            lcout => \DUT.rFifoDatarx_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_16_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12963\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15044\,
            ce => \N__11834\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_16_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__9264\,
            in1 => \N__11666\,
            in2 => \N__11073\,
            in3 => \N__11743\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_16_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__11673\,
            in1 => \N__12474\,
            in2 => \N__9276\,
            in3 => \N__11925\,
            lcout => \DUT.rFifoDatarx_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_16_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13011\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15044\,
            ce => \N__11834\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_16_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__11745\,
            in1 => \N__11064\,
            in2 => \N__11679\,
            in3 => \N__9258\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_16_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__12462\,
            in1 => \N__11913\,
            in2 => \N__9252\,
            in3 => \N__11675\,
            lcout => \DUT.rFifoDatarx_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__9234\,
            in1 => \N__11657\,
            in2 => \N__11058\,
            in3 => \N__11740\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__11662\,
            in1 => \N__12723\,
            in2 => \N__9243\,
            in3 => \N__11886\,
            lcout => \DUT.rFifoDatarx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13292\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15038\,
            ce => \N__11848\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_16_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__11739\,
            in1 => \N__11799\,
            in2 => \N__11677\,
            in3 => \N__9537\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__12711\,
            in1 => \N__11880\,
            in2 => \N__9228\,
            in3 => \N__11664\,
            lcout => \DUT.rFifoDatarx_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_16_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13058\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15038\,
            ce => \N__11848\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_16_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__9531\,
            in1 => \N__11658\,
            in2 => \N__11790\,
            in3 => \N__11741\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_16_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__11663\,
            in1 => \N__12699\,
            in2 => \N__9522\,
            in3 => \N__11874\,
            lcout => \DUT.rFifoDatarx_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNIME2J_0_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__9512\,
            in1 => \N__9476\,
            in2 => \N__9412\,
            in3 => \N__9332\,
            lcout => \DUT.fifo_tx_inst.rReadPtr11\,
            ltout => \DUT.fifo_tx_inst.rReadPtr11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rReadPtr_RNILV421_0_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010101010101"
        )
    port map (
            in0 => \N__14556\,
            in1 => \N__11636\,
            in2 => \N__9297\,
            in3 => \N__11728\,
            lcout => \DUT.fifo_tx_inst.un1_i11_2_i\,
            ltout => \DUT.fifo_tx_inst.un1_i11_2_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rReadPtr_1_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001010"
        )
    port map (
            in0 => \N__11637\,
            in1 => \N__11742\,
            in2 => \N__9294\,
            in3 => \N__9291\,
            lcout => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15031\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rReadPtr_0_LC_16_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__9290\,
            in1 => \N__9282\,
            in2 => \_gnd_net_\,
            in3 => \N__11729\,
            lcout => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15031\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111101111111"
        )
    port map (
            in0 => \N__11726\,
            in1 => \N__11936\,
            in2 => \N__11665\,
            in3 => \N__11948\,
            lcout => \DUT.rFifoDataror_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_0_RNI86BE_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111011101"
        )
    port map (
            in0 => \N__12012\,
            in1 => \N__11635\,
            in2 => \N__11964\,
            in3 => \N__11727\,
            lcout => \DUT.rFifoDataror_1\,
            ltout => \DUT.rFifoDataror_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_0_RNIKCMS_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9612\,
            in3 => \N__9605\,
            lcout => \DUT.rFifoDataror_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.rRamWrEn_latch_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__9731\,
            in1 => \N__15282\,
            in2 => \N__9765\,
            in3 => \N__9556\,
            lcout => \G_115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_0_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13569\,
            lcout => \DUT.wRxByte_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15026\,
            ce => \N__9783\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_1_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15146\,
            lcout => \DUT.wRxByte_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15026\,
            ce => \N__9783\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_2_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13515\,
            lcout => \DUT.wRxByte_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15026\,
            ce => \N__9783\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_3_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13467\,
            lcout => \DUT.wRxByte_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15026\,
            ce => \N__9783\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_4_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15081\,
            lcout => \DUT.wRxByte_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15026\,
            ce => \N__9783\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_5_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13415\,
            lcout => \DUT.wRxByte_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15026\,
            ce => \N__9783\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_6_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14066\,
            lcout => \DUT.wRxByte_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15026\,
            ce => \N__9783\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_7_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10517\,
            lcout => \DUT.wRxByte_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15026\,
            ce => \N__9783\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNIK68E1_1_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__11545\,
            in1 => \N__11157\,
            in2 => \_gnd_net_\,
            in3 => \N__11377\,
            lcout => \DUT.uart_inst0.m6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.un1_rWrState_1_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__9764\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9735\,
            lcout => \fifo_inst.ftdi_input_inst.un1_rWrStateZ0Z_1\,
            ltout => \fifo_inst.ftdi_input_inst.un1_rWrStateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_2_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__15281\,
            in1 => \N__9690\,
            in2 => \N__9714\,
            in3 => \N__9704\,
            lcout => \G_118\,
            ltout => \G_118_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.SUM_0_2_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__9640\,
            in1 => \_gnd_net_\,
            in2 => \N__9693\,
            in3 => \N__9676\,
            lcout => \G_119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_0_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__9839\,
            in1 => \N__10685\,
            in2 => \_gnd_net_\,
            in3 => \N__10071\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15020\,
            ce => \N__14456\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_4_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__10684\,
            in1 => \N__9840\,
            in2 => \N__11487\,
            in3 => \N__10289\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15020\,
            ce => \N__14456\,
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_0_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__15279\,
            in1 => \N__9659\,
            in2 => \_gnd_net_\,
            in3 => \N__9677\,
            lcout => \G_116\,
            ltout => \G_116_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_1_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__9660\,
            in1 => \N__9641\,
            in2 => \N__9651\,
            in3 => \N__15280\,
            lcout => \G_117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_2_1_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__11547\,
            in1 => \N__11039\,
            in2 => \N__9807\,
            in3 => \N__11153\,
            lcout => \DUT.uart_inst0.g1_i_a4_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_4_1_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10050\,
            in1 => \N__11256\,
            in2 => \N__11497\,
            in3 => \N__11379\,
            lcout => \DUT.uart_inst0.g1_i_a4_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_0_1_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__11380\,
            in1 => \N__10889\,
            in2 => \N__9920\,
            in3 => \N__10678\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_78_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_1_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111110000"
        )
    port map (
            in0 => \N__10424\,
            in1 => \_gnd_net_\,
            in2 => \N__9798\,
            in3 => \N__10952\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15014\,
            ce => \N__14461\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNIEQQU_1_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11546\,
            in2 => \_gnd_net_\,
            in3 => \N__11378\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_10_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNI2GC23_0_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001110100"
        )
    port map (
            in0 => \N__9899\,
            in1 => \N__10051\,
            in2 => \N__9795\,
            in3 => \N__10214\,
            lcout => \DUT.uart_inst0.P6_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_5_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__10215\,
            in1 => \N__9838\,
            in2 => \N__10706\,
            in3 => \N__11548\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15014\,
            ce => \N__14461\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_3_0_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__10221\,
            in1 => \N__11174\,
            in2 => \_gnd_net_\,
            in3 => \N__9981\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.G_19_0_a5_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_1_0_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__10153\,
            in1 => \N__10694\,
            in2 => \N__9786\,
            in3 => \N__10274\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.G_19_0_a5_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_0_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011111110"
        )
    port map (
            in0 => \N__10329\,
            in1 => \N__9846\,
            in2 => \N__10317\,
            in3 => \N__10313\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15009\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rReadPtr_0_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11048\,
            in1 => \N__13817\,
            in2 => \_gnd_net_\,
            in3 => \N__12573\,
            lcout => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15009\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNI8H662_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__10272\,
            in1 => \N__9977\,
            in2 => \_gnd_net_\,
            in3 => \N__10151\,
            lcout => \DUT.uart_inst0.G_8_i_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_2_3_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10273\,
            in2 => \_gnd_net_\,
            in3 => \N__10220\,
            lcout => \DUT.uart_inst0.m10_e_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rReadPtr_1_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__12572\,
            in1 => \N__13733\,
            in2 => \N__13821\,
            in3 => \N__11049\,
            lcout => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15009\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_3_3_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__10152\,
            in1 => \N__10080\,
            in2 => \N__9996\,
            in3 => \N__9907\,
            lcout => \DUT.uart_inst0.m10_e_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_2_0_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__10692\,
            in1 => \N__11564\,
            in2 => \N__11085\,
            in3 => \N__11480\,
            lcout => \DUT.uart_inst0.G_19_0_a5_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNIHH651_5_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__10927\,
            in1 => \N__10877\,
            in2 => \_gnd_net_\,
            in3 => \N__10565\,
            lcout => \DUT.uart_inst0.N_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_1_1_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__12301\,
            in1 => \N__12272\,
            in2 => \_gnd_net_\,
            in3 => \N__12241\,
            lcout => \DUT.fifo_tx_inst.rFifoData_awe0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rReadPtr_RNI4NC92_0_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011111111"
        )
    port map (
            in0 => \N__13736\,
            in1 => \N__13813\,
            in2 => \N__12566\,
            in3 => \N__14566\,
            lcout => \DUT.fifo_rx_inst.N_77_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNI237O_0_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__10564\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10925\,
            lcout => \DUT.uart_inst0.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_4_2_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__10926\,
            in1 => \N__10876\,
            in2 => \_gnd_net_\,
            in3 => \N__10566\,
            lcout => \DUT.uart_inst0.rx_countdown_8_i_a2_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_3_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100001111"
        )
    port map (
            in0 => \N__10836\,
            in1 => \N__11285\,
            in2 => \N__11336\,
            in3 => \N__10830\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_20_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_3_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110001000100"
        )
    port map (
            in0 => \N__11271\,
            in1 => \N__10821\,
            in2 => \N__10713\,
            in3 => \N__10693\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15005\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_4_6_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__11321\,
            in1 => \N__11493\,
            in2 => \N__10338\,
            in3 => \N__11264\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.m7_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_1_6_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__11562\,
            in1 => \N__11155\,
            in2 => \N__10581\,
            in3 => \N__11397\,
            lcout => \DUT.uart_inst0.N_28_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_5_6_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10556\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14572\,
            lcout => \DUT.uart_inst0.m2_e_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.oRxFlag_RNIHCKH1_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__15278\,
            in1 => \N__14812\,
            in2 => \_gnd_net_\,
            in3 => \N__12539\,
            lcout => \rTxByte_1_sqmuxa_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_5_3_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11563\,
            in1 => \N__11257\,
            in2 => \N__11499\,
            in3 => \N__11398\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.m6_e_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_1_3_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010111010101"
        )
    port map (
            in0 => \N__11322\,
            in1 => \N__11301\,
            in2 => \N__11289\,
            in3 => \N__11286\,
            lcout => \DUT.uart_inst0.N_18_mux_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_4_0_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__11263\,
            in1 => \N__11173\,
            in2 => \_gnd_net_\,
            in3 => \N__11154\,
            lcout => \DUT.uart_inst0.G_19_0_a5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_17_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13007\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15050\,
            ce => \N__11997\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_17_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12902\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15050\,
            ce => \N__11997\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_17_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12843\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15050\,
            ce => \N__11997\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_17_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13371\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15050\,
            ce => \N__11997\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_17_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13293\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15050\,
            ce => \N__11997\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_17_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13059\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15050\,
            ce => \N__11997\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_17_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13115\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15050\,
            ce => \N__11997\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_17_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12959\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15050\,
            ce => \N__11997\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_17_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__11751\,
            in1 => \N__11654\,
            in2 => \N__11775\,
            in3 => \N__11731\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_17_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__11656\,
            in1 => \N__12738\,
            in2 => \N__11763\,
            in3 => \N__11901\,
            lcout => \DUT.rFifoDatarx_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_17_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12839\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15045\,
            ce => \N__11852\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_17_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__11730\,
            in1 => \N__11688\,
            in2 => \N__11676\,
            in3 => \N__11580\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_17_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__12732\,
            in1 => \N__11892\,
            in2 => \N__11682\,
            in3 => \N__11655\,
            lcout => \DUT.rFifoDatarx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_17_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13367\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15045\,
            ce => \N__11852\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13000\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15039\,
            ce => \N__12207\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_17_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12895\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15039\,
            ce => \N__12207\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_17_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12838\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15039\,
            ce => \N__12207\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_17_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13366\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15039\,
            ce => \N__12207\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_17_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13285\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15039\,
            ce => \N__12207\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_17_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13051\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15039\,
            ce => \N__12207\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_17_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13108\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15039\,
            ce => \N__12207\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_17_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12958\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15039\,
            ce => \N__12207\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_3_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12083\,
            in2 => \_gnd_net_\,
            in3 => \N__12026\,
            lcout => \DUT.fifo_rx_inst.rFifoDataro_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15032\,
            ce => 'H',
            sr => \N__15231\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_0_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12011\,
            in2 => \_gnd_net_\,
            in3 => \N__11838\,
            lcout => \DUT.fifo_tx_inst.rFifoDataro_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15032\,
            ce => 'H',
            sr => \N__15231\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_1_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11963\,
            in2 => \_gnd_net_\,
            in3 => \N__11993\,
            lcout => \DUT.fifo_tx_inst.rFifoDataro_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15032\,
            ce => 'H',
            sr => \N__15231\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_2_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12203\,
            in2 => \_gnd_net_\,
            in3 => \N__11949\,
            lcout => \DUT.fifo_tx_inst.rFifoDataro_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15032\,
            ce => 'H',
            sr => \N__15231\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_3_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11937\,
            in2 => \_gnd_net_\,
            in3 => \N__12671\,
            lcout => \DUT.fifo_tx_inst.rFifoDataro_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15032\,
            ce => 'H',
            sr => \N__15231\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13612\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15027\,
            ce => \N__12084\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13570\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15027\,
            ce => \N__12084\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15147\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15027\,
            ce => \N__12084\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13516\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15027\,
            ce => \N__12084\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13468\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15027\,
            ce => \N__12084\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15082\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15027\,
            ce => \N__12084\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13416\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15027\,
            ce => \N__12084\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14067\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15027\,
            ce => \N__12084\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__13808\,
            in1 => \N__13700\,
            in2 => \N__14100\,
            in3 => \N__12048\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIT6K22_6_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__12057\,
            in1 => \N__13155\,
            in2 => \N__12051\,
            in3 => \N__13709\,
            lcout => \DUT.fifo_rx_inst.rFifoDatarx_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13426\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15021\,
            ce => \N__14859\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111110011"
        )
    port map (
            in0 => \N__14040\,
            in1 => \N__12033\,
            in2 => \N__13734\,
            in3 => \N__13809\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI1BK22_7_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__12042\,
            in1 => \N__13149\,
            in2 => \N__12036\,
            in3 => \N__13704\,
            lcout => \DUT.fifo_rx_inst.rFifoDatarx_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14086\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15021\,
            ce => \N__14859\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010101110101"
        )
    port map (
            in0 => \N__13807\,
            in1 => \N__12027\,
            in2 => \N__13735\,
            in3 => \N__12417\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoDataror_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_0_RNI5NR43_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110101"
        )
    port map (
            in0 => \N__12434\,
            in1 => \N__12450\,
            in2 => \N__12138\,
            in3 => \N__13708\,
            lcout => \DUT.fifo_rx_inst.rFifoDataror_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111110011"
        )
    port map (
            in0 => \N__13494\,
            in1 => \N__12123\,
            in2 => \N__13739\,
            in3 => \N__13810\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIHQJ22_3_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__12135\,
            in1 => \N__12759\,
            in2 => \N__12126\,
            in3 => \N__13731\,
            lcout => \DUT.fifo_rx_inst.rFifoDatarx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13536\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15015\,
            ce => \N__14866\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__13811\,
            in1 => \N__13446\,
            in2 => \N__12105\,
            in3 => \N__13729\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNILUJ22_4_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__13730\,
            in1 => \N__12117\,
            in2 => \N__12108\,
            in3 => \N__12747\,
            lcout => \DUT.fifo_rx_inst.rFifoDatarx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13480\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15015\,
            ce => \N__14866\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111110011"
        )
    port map (
            in0 => \N__13440\,
            in1 => \N__15063\,
            in2 => \N__13740\,
            in3 => \N__13812\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIP2K22_5_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__12096\,
            in1 => \N__13167\,
            in2 => \N__12087\,
            in3 => \N__13732\,
            lcout => \DUT.fifo_rx_inst.rFifoDatarx_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_0_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110111001100"
        )
    port map (
            in0 => \N__12349\,
            in1 => \N__12449\,
            in2 => \N__12401\,
            in3 => \N__12167\,
            lcout => \DUT.fifo_rx_inst.rFifoDataro_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15010\,
            ce => 'H',
            sr => \N__15224\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_1_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__12168\,
            in1 => \N__12396\,
            in2 => \N__12435\,
            in3 => \N__12350\,
            lcout => \DUT.fifo_rx_inst.rFifoDataro_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15010\,
            ce => 'H',
            sr => \N__15224\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_2_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__12351\,
            in1 => \N__12169\,
            in2 => \N__12402\,
            in3 => \N__12416\,
            lcout => \DUT.fifo_rx_inst.rFifoDataro_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15010\,
            ce => 'H',
            sr => \N__15224\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__12164\,
            in1 => \N__12388\,
            in2 => \_gnd_net_\,
            in3 => \N__12346\,
            lcout => \DUT.fifo_rx_inst.rFifoData_awe1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__12348\,
            in1 => \_gnd_net_\,
            in2 => \N__12400\,
            in3 => \N__12166\,
            lcout => \DUT.fifo_rx_inst.rFifoData_awe2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__12165\,
            in1 => \N__12389\,
            in2 => \_gnd_net_\,
            in3 => \N__12347\,
            lcout => \DUT.fifo_rx_inst.rFifoData_awe0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_1_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__12313\,
            in1 => \N__12276\,
            in2 => \_gnd_net_\,
            in3 => \N__12242\,
            lcout => \DUT.fifo_tx_inst.rFifoData_awe2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12604\,
            in2 => \_gnd_net_\,
            in3 => \N__13895\,
            lcout => \DUT.fifo_rx_inst.rWritePtr16\,
            ltout => \DUT.fifo_rx_inst.rWritePtr16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__13925\,
            in1 => \N__14011\,
            in2 => \N__12186\,
            in3 => \N__13947\,
            lcout => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_0_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101000111100"
        )
    port map (
            in0 => \N__13949\,
            in1 => \N__12170\,
            in2 => \N__14015\,
            in3 => \N__13928\,
            lcout => \DUT.fifo_rx_inst.rFifoCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15006\,
            ce => 'H',
            sr => \N__15223\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNI110Q1_1_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__13894\,
            in1 => \N__13968\,
            in2 => \N__12609\,
            in3 => \N__14005\,
            lcout => \DUT.fifo_rx_inst.N_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNI9EGD1_1_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__14006\,
            in1 => \N__13924\,
            in2 => \N__13976\,
            in3 => \N__13896\,
            lcout => \DUT.fifo_rx_inst.N_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNIPTFQ1_1_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13926\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13948\,
            lcout => \DUT.fifo_rx_inst.rFifoCount_RNIPTFQ1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_1_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__14007\,
            in1 => \_gnd_net_\,
            in2 => \N__13977\,
            in3 => \N__13897\,
            lcout => \N_69_mux\,
            ltout => \N_69_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rRxRead_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__13927\,
            in1 => \_gnd_net_\,
            in2 => \N__12528\,
            in3 => \N__14813\,
            lcout => \rRxReadZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15006\,
            ce => 'H',
            sr => \N__15223\
        );

    \ioFifoData_iobuf_RNO_1_LC_18_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13851\,
            lcout => \N_1258_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.oTx_n_RNIPDL9_LC_18_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14215\,
            lcout => \P1A4_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_18_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12999\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15051\,
            ce => \N__12678\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_18_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12894\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15051\,
            ce => \N__12678\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_18_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12837\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15051\,
            ce => \N__12678\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_18_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13365\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15051\,
            ce => \N__12678\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_18_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13275\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15051\,
            ce => \N__12678\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_18_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13050\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15051\,
            ce => \N__12678\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_18_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13104\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15051\,
            ce => \N__12678\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_18_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12948\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15051\,
            ce => \N__12678\,
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rRxData_esr_3_LC_18_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12648\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \wRxFifoData_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15046\,
            ce => \N__14267\,
            sr => \N__15240\
        );

    \fifo_inst.ftdi_output_inst.rRxData_esr_1_LC_18_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12633\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \wRxFifoData_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15040\,
            ce => \N__14268\,
            sr => \N__15236\
        );

    \fifo_inst.ftdi_output_inst.rRxData_esr_5_LC_18_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12618\,
            lcout => \wRxFifoData_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15040\,
            ce => \N__14268\,
            sr => \N__15236\
        );

    \fifo_inst.ftdi_output_inst.rRxData_esr_2_LC_18_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12810\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \wRxFifoData_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15040\,
            ce => \N__14268\,
            sr => \N__15236\
        );

    \fifo_inst.ftdi_output_inst.rRxData_esr_0_LC_18_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12798\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \wRxFifoData_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15040\,
            ce => \N__14268\,
            sr => \N__15236\
        );

    \fifo_inst.ftdi_output_inst.rRxData_esr_6_LC_18_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12786\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \wRxFifoData_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15040\,
            ce => \N__14268\,
            sr => \N__15236\
        );

    \fifo_inst.ftdi_output_inst.rRxData_esr_4_LC_18_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12771\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \wRxFifoData_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15040\,
            ce => \N__14268\,
            sr => \N__15236\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13630\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15033\,
            ce => \N__13143\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13588\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15033\,
            ce => \N__13143\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15166\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15033\,
            ce => \N__13143\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13534\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15033\,
            ce => \N__13143\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13487\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15033\,
            ce => \N__13143\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15106\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15033\,
            ce => \N__13143\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13433\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15033\,
            ce => \N__13143\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14087\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15033\,
            ce => \N__13143\,
            sr => \_gnd_net_\
        );

    \rTxByte_esr_6_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011001010"
        )
    port map (
            in0 => \N__13131\,
            in1 => \N__13125\,
            in2 => \N__14826\,
            in3 => \N__13337\,
            lcout => \rTxByteZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15028\,
            ce => \N__13257\,
            sr => \N__15230\
        );

    \rTxByte_esr_5_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__13336\,
            in1 => \N__14819\,
            in2 => \N__13077\,
            in3 => \N__13065\,
            lcout => \rTxByteZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15028\,
            ce => \N__13257\,
            sr => \N__15230\
        );

    \rTxByte_esr_0_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__14814\,
            in1 => \N__13221\,
            in2 => \N__13023\,
            in3 => \N__13331\,
            lcout => \rTxByteZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15028\,
            ce => \N__13257\,
            sr => \N__15230\
        );

    \rTxByte_esr_7_LC_18_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__13338\,
            in1 => \N__14823\,
            in2 => \N__14286\,
            in3 => \N__12969\,
            lcout => \rTxByteZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15028\,
            ce => \N__13257\,
            sr => \N__15230\
        );

    \rTxByte_esr_1_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__14815\,
            in1 => \N__13185\,
            in2 => \N__12915\,
            in3 => \N__13332\,
            lcout => \rTxByteZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15028\,
            ce => \N__13257\,
            sr => \N__15230\
        );

    \rTxByte_esr_2_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__13333\,
            in1 => \N__14816\,
            in2 => \N__12855\,
            in3 => \N__13638\,
            lcout => \rTxByteZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15028\,
            ce => \N__13257\,
            sr => \N__15230\
        );

    \rTxByte_esr_3_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__14817\,
            in1 => \N__13389\,
            in2 => \N__13383\,
            in3 => \N__13334\,
            lcout => \rTxByteZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15028\,
            ce => \N__13257\,
            sr => \N__15230\
        );

    \rTxByte_esr_4_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__13335\,
            in1 => \N__14818\,
            in2 => \N__13311\,
            in3 => \N__13299\,
            lcout => \rTxByteZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15028\,
            ce => \N__13257\,
            sr => \N__15230\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111110011"
        )
    port map (
            in0 => \N__13596\,
            in1 => \N__13215\,
            in2 => \N__13737\,
            in3 => \N__13815\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI5EJ22_0_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__13245\,
            in1 => \N__13236\,
            in2 => \N__13224\,
            in3 => \N__13721\,
            lcout => \DUT.fifo_rx_inst.rFifoDatarx_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13631\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15022\,
            ce => \N__14867\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__13814\,
            in1 => \N__13548\,
            in2 => \N__13179\,
            in3 => \N__13716\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI9IJ22_1_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__13720\,
            in1 => \N__13209\,
            in2 => \N__13197\,
            in3 => \N__13194\,
            lcout => \DUT.fifo_rx_inst.rFifoDatarx_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13589\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15022\,
            ce => \N__14867\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111110011"
        )
    port map (
            in0 => \N__13542\,
            in1 => \N__15120\,
            in2 => \N__13738\,
            in3 => \N__13816\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIDMJ22_2_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__13764\,
            in1 => \N__13752\,
            in2 => \N__13743\,
            in3 => \N__13722\,
            lcout => \DUT.fifo_rx_inst.rFifoDatarx_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13632\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15016\,
            ce => \N__14028\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13590\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15016\,
            ce => \N__14028\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15167\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15016\,
            ce => \N__14028\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13535\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15016\,
            ce => \N__14028\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13488\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15016\,
            ce => \N__14028\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15111\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15016\,
            ce => \N__14028\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13434\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15016\,
            ce => \N__14028\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14088\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15016\,
            ce => \N__14028\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14022\,
            in2 => \N__14016\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_12_0_\,
            carryout => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_1_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13975\,
            in2 => \N__13986\,
            in3 => \N__13953\,
            lcout => \DUT.fifo_rx_inst.rFifoCountZ0Z_1\,
            ltout => OPEN,
            carryin => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0\,
            carryout => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1\,
            clk => \N__15011\,
            ce => 'H',
            sr => \N__15225\
        );

    \DUT.fifo_rx_inst.rFifoCount_2_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001010101101010"
        )
    port map (
            in0 => \N__13901\,
            in1 => \N__13950\,
            in2 => \N__13932\,
            in3 => \N__13905\,
            lcout => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15011\,
            ce => 'H',
            sr => \N__15225\
        );

    \ioFifoData_iobuf_RNO_4_LC_20_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13860\,
            lcout => \N_1261_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.oTx_n_rep4_ess_LC_20_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__15358\,
            in1 => \_gnd_net_\,
            in2 => \N__15422\,
            in3 => \_gnd_net_\,
            lcout => \oTx_n_rep4_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15053\,
            ce => \N__15302\,
            sr => \N__15248\
        );

    \fifo_inst.ftdi_output_inst.oTx_n_rep1_ess_LC_20_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__15357\,
            in1 => \_gnd_net_\,
            in2 => \N__15421\,
            in3 => \_gnd_net_\,
            lcout => \oTx_n_rep1_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15053\,
            ce => \N__15302\,
            sr => \N__15248\
        );

    \fifo_inst.ftdi_output_inst.oTx_n_rep0_ess_LC_20_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15410\,
            in2 => \_gnd_net_\,
            in3 => \N__15356\,
            lcout => \oTx_n_rep0_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15053\,
            ce => \N__15302\,
            sr => \N__15248\
        );

    \fifo_inst.ftdi_output_inst.oRamRdAddr_0_LC_20_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__15341\,
            in1 => \N__14567\,
            in2 => \N__15408\,
            in3 => \N__14172\,
            lcout => \fifo_inst.wRamRdAddr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_RNIFFVH_4_LC_20_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15387\,
            in2 => \_gnd_net_\,
            in3 => \N__15339\,
            lcout => \fifo_inst.ftdi_output_inst.N_77_0\,
            ltout => \fifo_inst.ftdi_output_inst.N_77_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_RNIUEQM_3_LC_20_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15290\,
            in2 => \N__14235\,
            in3 => \N__14113\,
            lcout => \fifo_inst.ftdi_output_inst.N_88_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.oTx_n_LC_20_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101001111"
        )
    port map (
            in0 => \N__14114\,
            in1 => \N__14197\,
            in2 => \N__14577\,
            in3 => \N__14336\,
            lcout => \P1A4_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_RNIBT9K_4_LC_20_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__14571\,
            in1 => \N__15388\,
            in2 => \_gnd_net_\,
            in3 => \N__15340\,
            lcout => \fifo_inst.ftdi_output_inst.oPacketRead_1_sqmuxa_1\,
            ltout => \fifo_inst.ftdi_output_inst.oPacketRead_1_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.oRamRdAddr_1_LC_20_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14149\,
            in2 => \N__14181\,
            in3 => \N__14173\,
            lcout => \fifo_inst.wRamRdAddr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.oRamRdAddr_2_LC_20_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__14174\,
            in1 => \N__14126\,
            in2 => \N__14156\,
            in3 => \N__14136\,
            lcout => \fifo_inst.wRamRdAddr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_3_LC_20_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__14324\,
            in1 => \N__14648\,
            in2 => \N__14679\,
            in3 => \N__14603\,
            lcout => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15048\,
            ce => 'H',
            sr => \N__15241\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_4_LC_20_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100001010"
        )
    port map (
            in0 => \N__15343\,
            in1 => \_gnd_net_\,
            in2 => \N__15409\,
            in3 => \N__14115\,
            lcout => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15048\,
            ce => 'H',
            sr => \N__15241\
        );

    \fifo_inst.ftdi_output_inst.rWrDelay_LC_20_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15392\,
            in2 => \_gnd_net_\,
            in3 => \N__15342\,
            lcout => \fifo_inst.ftdi_output_inst.rWrDelayZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15048\,
            ce => 'H',
            sr => \N__15241\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_1_LC_20_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__14647\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14323\,
            lcout => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15048\,
            ce => 'H',
            sr => \N__15241\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_2_LC_20_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14694\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15048\,
            ce => 'H',
            sr => \N__15241\
        );

    \fifo_inst.ftdi_output_inst.oRxFlag_LC_20_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__14357\,
            in1 => \N__14773\,
            in2 => \_gnd_net_\,
            in3 => \N__14693\,
            lcout => \P1A2_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15048\,
            ce => 'H',
            sr => \N__15241\
        );

    \fifo_inst.ftdi_output_inst.oRx_n_LC_20_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110110011101110"
        )
    port map (
            in0 => \N__14710\,
            in1 => \N__14356\,
            in2 => \N__14649\,
            in3 => \N__14325\,
            lcout => \P1A3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15048\,
            ce => 'H',
            sr => \N__15241\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_RNIDTQ4_1_LC_20_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15283\,
            in2 => \_gnd_net_\,
            in3 => \N__14692\,
            lcout => \fifo_inst.ftdi_output_inst.rFifoState_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_RNO_0_0_LC_20_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110000000000"
        )
    port map (
            in0 => \N__14669\,
            in1 => \N__14636\,
            in2 => \N__14607\,
            in3 => \N__14322\,
            lcout => OPEN,
            ltout => \fifo_inst.ftdi_output_inst.N_87_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_0_LC_20_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__14573\,
            in1 => \N__14358\,
            in2 => \N__14343\,
            in3 => \N__14340\,
            lcout => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15041\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rRxData_esr_7_LC_20_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14307\,
            lcout => \wRxFifoData_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15034\,
            ce => \N__14266\,
            sr => \N__15232\
        );

    \ioFifoData_iobuf_RNO_3_LC_21_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15432\,
            lcout => \N_1260_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ioFifoData_iobuf_RNO_2_LC_21_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15312\,
            lcout => \N_1259_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.oTx_n_rep3_ess_LC_21_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__15360\,
            in1 => \_gnd_net_\,
            in2 => \N__15423\,
            in3 => \_gnd_net_\,
            lcout => \oTx_n_rep3_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15054\,
            ce => \N__15303\,
            sr => \N__15249\
        );

    \fifo_inst.ftdi_output_inst.oTx_n_rep2_ess_LC_21_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15417\,
            in2 => \_gnd_net_\,
            in3 => \N__15359\,
            lcout => \oTx_n_rep2_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15054\,
            ce => \N__15303\,
            sr => \N__15249\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_21_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15171\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15042\,
            ce => \N__14868\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_21_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15110\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__15042\,
            ce => \N__14868\,
            sr => \_gnd_net_\
        );
end \INTERFACE\;
