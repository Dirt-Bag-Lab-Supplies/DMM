-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Mar 29 2020 23:01:15

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    ioFifoData : out std_logic_vector(7 downto 0);
    P1A9 : out std_logic;
    P1A1 : in std_logic;
    P1A8 : out std_logic;
    oRx_n : out std_logic;
    P1A7 : out std_logic;
    P1A3 : out std_logic;
    iTxE_n : in std_logic;
    iRxF_n : in std_logic;
    iClk : in std_logic;
    P1A2 : out std_logic;
    BTN_N : in std_logic;
    BTN1 : in std_logic;
    oTx_n : out std_logic;
    P1A4 : out std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__13526\ : std_logic;
signal \N__13512\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13501\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13483\ : std_logic;
signal \N__13476\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13458\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13438\ : std_logic;
signal \N__13431\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13429\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13412\ : std_logic;
signal \N__13411\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13402\ : std_logic;
signal \N__13395\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13377\ : std_logic;
signal \N__13376\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13366\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13357\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13321\ : std_logic;
signal \N__13320\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13310\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13302\ : std_logic;
signal \N__13299\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13277\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13274\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13254\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13248\ : std_logic;
signal \N__13245\ : std_logic;
signal \N__13242\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13209\ : std_logic;
signal \N__13204\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13164\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13158\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13105\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13067\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13058\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13048\ : std_logic;
signal \N__13047\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13039\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13034\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13028\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13006\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13003\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12856\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12847\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12841\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12814\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12760\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12757\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12748\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12715\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12703\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12695\ : std_logic;
signal \N__12692\ : std_logic;
signal \N__12689\ : std_logic;
signal \N__12686\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12605\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12596\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12569\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12551\ : std_logic;
signal \N__12548\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12527\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12382\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12362\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12311\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12227\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12208\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12189\ : std_logic;
signal \N__12182\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12067\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12001\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11767\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11714\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11240\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10434\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10232\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7893\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7629\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6993\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6705\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5672\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5174\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5159\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \BTN_N_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remaining_RNO_1Z0Z_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.m5_1_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_6_0_0\ : std_logic;
signal \DUT.uart_inst0.N_6_0_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_15_mux_0\ : std_logic;
signal \DUT.uart_inst0.recv_state_ns_0_i_a2_0_2_3_cascade_\ : std_logic;
signal \DUT.uart_inst0.m16_N_3L3_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remaining_RNO_4Z0Z_1\ : std_logic;
signal \DUT.uart_inst0.g0_i_a3_5_cascade_\ : std_logic;
signal \DUT.uart_inst0.g0_0_i_a3_0_3\ : std_logic;
signal \DUT.uart_inst0.g0_0_i_a3_0_4_cascade_\ : std_logic;
signal \DUT.uart_inst0.g0_0\ : std_logic;
signal \DUT.uart_inst0.g0_i_a3_0_5_cascade_\ : std_logic;
signal \DUT.uart_inst0.g0_i_a3_8\ : std_logic;
signal \DUT.uart_inst0.g0_i_a3_0_6\ : std_logic;
signal \DUT.uart_inst0.g0_i_a3_0_7_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_6_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_40\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remainingZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remainingZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.recv_state_RNIL139CZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.N_35_0\ : std_logic;
signal \DUT.uart_inst0.g0_0_2_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remainingZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.m8_e_3\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remainingZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.g0_i_a3_6\ : std_logic;
signal \DUT.uart_inst0.recv_state_ns_0_i_a2_0_0_3\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.g0_0_0\ : std_logic;
signal \DUT.uart_inst0.g0_0_1\ : std_logic;
signal \DUT.uart_inst0.N_81_mux_i_i_a5_0_4_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_81_mux_i_i_a5_0_4\ : std_logic;
signal \DUT.uart_inst0.N_81_mux_i_i_0\ : std_logic;
signal \DUT.uart_inst0.N_81_mux_i_i_a5_0_5_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_81_mux_i_i_a5_1_5\ : std_logic;
signal \DUT.uart_inst0.m8_e_2\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_0_s1\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_1_s1\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_2_s1\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_3_s1\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_4_s1\ : std_logic;
signal \DUT.uart_inst0.m9_3\ : std_logic;
signal \DUT.uart_inst0.m9_4\ : std_logic;
signal \DUT.uart_inst0.N_8\ : std_logic;
signal \DUT.uart_inst0.N_81_mux_i_i_0_0\ : std_logic;
signal \DUT.uart_inst0.N_81_mux_i_i_a5_0_5_0\ : std_logic;
signal \DUT.uart_inst0.m4_3_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_18_mux\ : std_logic;
signal \DUT.uart_inst0.N_297_cascade_\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.N_15_3\ : std_logic;
signal \DUT.uart_inst0.g0_0_i_a3_3_cascade_\ : std_logic;
signal \DUT.uart_inst0.g0_0_i_a3_4\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_2\ : std_logic;
signal \wPllLocked_i\ : std_logic;
signal \bfn_8_18_0_\ : std_logic;
signal \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0\ : std_logic;
signal \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_awe3_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.un1_i11_i_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.un1_rFifoCount_1_axb_2\ : std_logic;
signal \DUT.fifo_rx_inst.un1_i11_i\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoCount_RNIK3G92Z0Z_1\ : std_logic;
signal \DUT.fifo_rx_inst.rWritePtr16_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rWritePtr16\ : std_logic;
signal \DUT.fifo_rx_inst.rWritePtrZ0Z_0\ : std_logic;
signal \DUT.fifo_rx_inst.rWritePtrZ0Z_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_6\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_5\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_5\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_6\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_5\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_6\ : std_logic;
signal \DUT.uart_inst0.N_81_mux_i_i_a5_1_4\ : std_logic;
signal \DUT.uart_inst0.N_13_0\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_RNO_2Z0Z_2\ : std_logic;
signal \DUT.uart_inst0.G_21_0_1_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.G_9_i_o4_0\ : std_logic;
signal \DUT.uart_inst0.g0_0_3\ : std_logic;
signal \DUT.uart_inst0.G_16_i_a3_0_2_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_45_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_55\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_s1_4\ : std_logic;
signal \DUT.uart_inst0.N_10\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.G_21_0_1\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.N_45\ : std_logic;
signal \DUT.uart_inst0.recv_state_ns_0_0_0\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_s1_2\ : std_logic;
signal \DUT.uart_inst0.G_16_i_a3_0_3\ : std_logic;
signal \DUT.uart_inst0.g1_1\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_s1_1\ : std_logic;
signal \DUT.uart_inst0.N_81_mux_i_i_a5_1_5_0\ : std_logic;
signal \DUT.uart_inst0.N_81_mux_i_i_a5_1_3\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_s1_3\ : std_logic;
signal \DUT.uart_inst0.N_300_cascade_\ : std_logic;
signal \DUT.uart_inst0.G_16_i_a3_3_cascade_\ : std_logic;
signal \DUT.uart_inst0.G_16_i_a3_4\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.N_11_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_awe3_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.un1_i11_i\ : std_logic;
signal \DUT.fifo_tx_inst.un1_i11_i_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ1Z_3\ : std_logic;
signal \DUT.uart_inst0.N_13_mux\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_s1_5\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.N_8_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.m10_0_1\ : std_logic;
signal \DUT.uart_inst0.m11_0\ : std_logic;
signal \DUT.uart_inst0.N_15_mux\ : std_logic;
signal \DUT.uart_inst0.N_11_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa\ : std_logic;
signal \DUT.fifo_rx_inst.N_87_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0\ : std_logic;
signal \DUT.wRcvd\ : std_logic;
signal \DUT.fifo_rx_inst.N_87\ : std_logic;
signal \DUT.fifo_rx_inst.N_92_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoCountZ0Z_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoCountZ0Z_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoCountZ0Z_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_awe2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_awe2_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoDataro_3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoDataro_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_awe0_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDataro_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_awe1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDataro_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_awe2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDataro_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDataro_2\ : std_logic;
signal \DUT.fifo_rx_inst.rTxByte_42_1\ : std_logic;
signal \DUT.fifo_rx_inst.rTxByte_42_0_cascade_\ : std_logic;
signal \N_92_i\ : std_logic;
signal \rFifoDatarff_0_RNIHJV05_cascade_\ : std_logic;
signal \DUT.wRxByte_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_0\ : std_logic;
signal \DUT.wRxByte_1\ : std_logic;
signal \DUT.wRxByte_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_2\ : std_logic;
signal \DUT.wRxByte_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_3\ : std_logic;
signal \DUT.wRxByte_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_4\ : std_logic;
signal \DUT.wRxByte_5\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_5\ : std_logic;
signal \DUT.wRxByte_6\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_6\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_awe3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7\ : std_logic;
signal \P1A3_c\ : std_logic;
signal \fifo_inst.ft2232h_inst.rFifoStateZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_10\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_0\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_11\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_12\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_9\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_13\ : std_logic;
signal \DUT.uart_inst0.un1_N_5_mux_cascade_\ : std_logic;
signal \DUT.uart_inst0.g0_i_o6_0_4_cascade_\ : std_logic;
signal \DUT.uart_inst0.g0_i_o6_0_5\ : std_logic;
signal \DUT.uart_inst0.N_139_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remaining_RNO_1Z0Z_3\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_6\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_7\ : std_logic;
signal \DUT.uart_inst0.N_22_i\ : std_logic;
signal \DUT.uart_inst0.N_79_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_state_ns_i_i_0_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_2\ : std_logic;
signal \DUT.rFifoDatarx_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_\ : std_logic;
signal \DUT.rFifoDatarx_3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoDataro_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoDataro_1\ : std_logic;
signal \DUT.rFifoDataror_1\ : std_logic;
signal \DUT.rFifoDataror_1_cascade_\ : std_logic;
signal \DUT.rFifoDataror_0_0\ : std_logic;
signal \DUT.rFifoDataror_0\ : std_logic;
signal \wPllLocked\ : std_logic;
signal \DUT.fifo_rx_inst.CO0\ : std_logic;
signal \DUT.fifo_rx_inst.un1_i11_2_i\ : std_logic;
signal \DUT.fifo_rx_inst.un1_i11_2_i_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.N_92\ : std_logic;
signal \DUT.fifo_rx_inst.rReadPtrZ0Z_0\ : std_logic;
signal \DUT.fifo_tx_inst.rWritePtrZ0Z_0\ : std_logic;
signal \DUT.fifo_tx_inst.rWritePtrZ0Z_1\ : std_logic;
signal \DUT.fifo_tx_inst.N_83_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.N_88\ : std_logic;
signal \DUT.fifo_tx_inst.N_88_cascade_\ : std_logic;
signal \DUT.rTransmitc\ : std_logic;
signal \DUT.fifo_tx_inst.rWritePtr16\ : std_logic;
signal \DUT.fifo_tx_inst.un1_i11_2_i\ : std_logic;
signal \DUT.fifo_rx_inst.rReadPtrZ0Z_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1\ : std_logic;
signal \N_92_i_0\ : std_logic;
signal \rFifoDatarff_0_RNIHJV05\ : std_logic;
signal \fifo_inst.ft2232h_inst.rFifoStateZ0Z_2\ : std_logic;
signal \P1A4_c\ : std_logic;
signal \fifo_inst.ft2232h_inst.rFifoStateZ0Z_3\ : std_logic;
signal \rTxBusReady\ : std_logic;
signal \fifo_inst.ft2232h_inst.rFifoStateZ0Z_4\ : std_logic;
signal \fifo_inst.ft2232h_inst.rTxRdEnZ0\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_1\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ1Z_1\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_0\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_1\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_2_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_2\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_3\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_4_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_4\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_6\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_5_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_5\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_7\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_6\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_7\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_8\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_9\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_8\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_10\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_9\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_11\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_10\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_11\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_13\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_12\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_14\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_13\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_15\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_14\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_15\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_16\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_16\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_17\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_12\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.N_50\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.N_98_cascade_\ : std_logic;
signal \P1A7_c\ : std_logic;
signal \DUT.uart_inst0.N_82\ : std_logic;
signal \DUT.uart_inst0.N_99\ : std_logic;
signal \DUT.uart_inst0.N_100\ : std_logic;
signal \P1A1_c\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.N_49\ : std_logic;
signal \fifo_inst.ft2232h_inst.rFifoStatec_0\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remainingZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.N_139\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remainingZ0Z_2\ : std_logic;
signal \DUT.rTransmitc_0\ : std_logic;
signal \DUT.uart_inst0.N_85_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_66\ : std_logic;
signal \DUT.uart_inst0.N_22_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remainingZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.N_22\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remainingZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.N_65_i\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.N_85\ : std_logic;
signal \DUT.uart_inst0.N_89\ : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_0\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_1\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_2\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_3\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_4\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_5\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_6\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_7\ : std_logic;
signal \bfn_11_19_0_\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_8\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_9\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_10\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_11\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_12\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_\ : std_logic;
signal \DUT.rFifoDatarx_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_0\ : std_logic;
signal \DUT.rFifoDatarxZ0Z_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1_cascade_\ : std_logic;
signal \DUT.rFifoDatarx_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_4\ : std_logic;
signal \DUT.rFifoDatarx_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_\ : std_logic;
signal \DUT.rFifoDatarx_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_5\ : std_logic;
signal \DUT.fifo_tx_inst.rReadPtrZ0Z_0\ : std_logic;
signal \DUT.fifo_tx_inst.rReadPtrZ0Z_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_6\ : std_logic;
signal \DUT.rFifoDatarx_6\ : std_logic;
signal \DUT.rFifoCount_0\ : std_logic;
signal \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0\ : std_logic;
signal \bfn_11_22_0_\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoCount_RNIBPFMZ0Z_1\ : std_logic;
signal \DUT.rFifoCount_1\ : std_logic;
signal \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0\ : std_logic;
signal \rRxReadZ0\ : std_logic;
signal \DUT.fifo_tx_inst.N_83\ : std_logic;
signal \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1\ : std_logic;
signal \DUT.rFifoCount_2\ : std_logic;
signal \wPllLocked_i_g\ : std_logic;
signal \DUT.wRxByte_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_awe0\ : std_logic;
signal \iRxF_n_c\ : std_logic;
signal \iTxE_n_c\ : std_logic;
signal \fifo_inst.ft2232h_inst.rFifoStateZ0Z_0\ : std_logic;
signal \fifo_inst.ft2232h_inst.N_101\ : std_logic;
signal \DUT.uart_inst0.N_13_cascade_\ : std_logic;
signal \DUT.uart_inst0.g0_i_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.g0_i_a6_0\ : std_logic;
signal \DUT.uart_inst0.g0_i_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.g0_i_a6_3_0\ : std_logic;
signal \DUT.uart_inst0.g0_i_o2_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_77\ : std_logic;
signal \DUT.uart_inst0.g0_i_o2_2\ : std_logic;
signal \DUT.uart_inst0.g0_i_o2_3\ : std_logic;
signal \DUT.uart_inst0.N_11\ : std_logic;
signal \DUT.uart_inst0.g0_11_a4_2\ : std_logic;
signal \DUT.uart_inst0.N_9\ : std_logic;
signal \DUT.uart_inst0.tx_state_ns_i_i_o2_a0_2_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_71_i\ : std_logic;
signal \DUT.uart_inst0.N_8_1\ : std_logic;
signal \DUT.uart_inst0.g0_i_a3_0_cascade_\ : std_logic;
signal \wPllLocked_g\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0\ : std_logic;
signal \DUT.uart_inst0.g0_11_a3_2_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_7\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.N_6_i\ : std_logic;
signal \DUT.rTransmitZ0\ : std_logic;
signal \DUT.tx_state_0\ : std_logic;
signal \DUT.uart_inst0.tx_stateZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.N_11_1\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_9\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_10\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_11\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_8\ : std_logic;
signal \DUT.uart_inst0.N_20\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_12\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_7\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_13\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_6\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_9\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_7\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_8_cascade_\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_6\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_0\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_5_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_6\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_awe3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_1\ : std_logic;
signal \rTxByteZ0Z_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_2\ : std_logic;
signal \rTxByteZ0Z_3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_3\ : std_logic;
signal \rTxByteZ0Z_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_6\ : std_logic;
signal \rTxByteZ0Z_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_7\ : std_logic;
signal \rTxByteZ0Z_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_1\ : std_logic;
signal \rTxByteZ0Z_6\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_6\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_awe0\ : std_logic;
signal \rTxByteZ0Z_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_5\ : std_logic;
signal \rTxByteZ0Z_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_0\ : std_logic;
signal clk_48mhz : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_awe1\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \iClk_wire\ : std_logic;
signal \P1A8_wire\ : std_logic;
signal \ioFifoData_wire\ : std_logic_vector(7 downto 0);
signal \P1A9_wire\ : std_logic;
signal \P1A2_wire\ : std_logic;
signal \P1A4_wire\ : std_logic;
signal \oRx_n_wire\ : std_logic;
signal \iRxF_n_wire\ : std_logic;
signal \P1A3_wire\ : std_logic;
signal \P1A7_wire\ : std_logic;
signal \BTN_N_wire\ : std_logic;
signal \oTx_n_wire\ : std_logic;
signal \iTxE_n_wire\ : std_logic;
signal \P1A1_wire\ : std_logic;
signal \top_pll_inst.top_pll_inst_pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \iClk_wire\ <= iClk;
    P1A8 <= \P1A8_wire\;
    ioFifoData <= \ioFifoData_wire\;
    P1A9 <= \P1A9_wire\;
    P1A2 <= \P1A2_wire\;
    P1A4 <= \P1A4_wire\;
    oRx_n <= \oRx_n_wire\;
    \iRxF_n_wire\ <= iRxF_n;
    P1A3 <= \P1A3_wire\;
    P1A7 <= \P1A7_wire\;
    \BTN_N_wire\ <= BTN_N;
    oTx_n <= \oTx_n_wire\;
    \iTxE_n_wire\ <= iTxE_n;
    \P1A1_wire\ <= P1A1;
    \top_pll_inst.top_pll_inst_pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \top_pll_inst.top_pll_inst_pll\ : PLL40
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "0111111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            PLLOUTGLOBAL => clk_48mhz,
            SDI => \GNDG0\,
            BYPASS => \GNDG0\,
            RESETB => \N__5081\,
            PLLOUTCORE => OPEN,
            LOCK => \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO\,
            SDO => OPEN,
            SCLK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            EXTFEEDBACK => \GNDG0\,
            DYNAMICDELAY => \top_pll_inst.top_pll_inst_pll_DYNAMICDELAY_wire\,
            PLLIN => \N__13526\
        );

    \top_pll_inst.top_pll_inst_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \VCCG0\,
            DIN => '0',
            DOUT => \N__13526\,
            PACKAGEPIN => \iClk_wire\
        );

    \P1A8_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13512\,
            DIN => \N__13511\,
            DOUT => \N__13510\,
            PACKAGEPIN => \P1A8_wire\
        );

    \P1A8_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13512\,
            PADOUT => \N__13511\,
            PADIN => \N__13510\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13503\,
            DIN => \N__13502\,
            DOUT => \N__13501\,
            PACKAGEPIN => \ioFifoData_wire\(1)
        );

    \ioFifoData_obuft_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13503\,
            PADOUT => \N__13502\,
            PADIN => \N__13501\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8698\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A9_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13494\,
            DIN => \N__13493\,
            DOUT => \N__13492\,
            PACKAGEPIN => \P1A9_wire\
        );

    \P1A9_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13494\,
            PADOUT => \N__13493\,
            PADIN => \N__13492\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13485\,
            DIN => \N__13484\,
            DOUT => \N__13483\,
            PACKAGEPIN => \ioFifoData_wire\(4)
        );

    \ioFifoData_obuft_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13485\,
            PADOUT => \N__13484\,
            PADIN => \N__13483\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8743\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A2_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13476\,
            DIN => \N__13475\,
            DOUT => \N__13474\,
            PACKAGEPIN => \P1A2_wire\
        );

    \P1A2_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13476\,
            PADOUT => \N__13475\,
            PADIN => \N__13474\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A4_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13467\,
            DIN => \N__13466\,
            DOUT => \N__13465\,
            PACKAGEPIN => \P1A4_wire\
        );

    \P1A4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13467\,
            PADOUT => \N__13466\,
            PADIN => \N__13465\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8800\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13458\,
            DIN => \N__13457\,
            DOUT => \N__13456\,
            PACKAGEPIN => \ioFifoData_wire\(0)
        );

    \ioFifoData_obuft_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13458\,
            PADOUT => \N__13457\,
            PADIN => \N__13456\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8722\,
            DIN0 => OPEN,
            DOUT0 => \N__12841\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \oRx_n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13449\,
            DIN => \N__13448\,
            DOUT => \N__13447\,
            PACKAGEPIN => \oRx_n_wire\
        );

    \oRx_n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13449\,
            PADOUT => \N__13448\,
            PADIN => \N__13447\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7550\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13440\,
            DIN => \N__13439\,
            DOUT => \N__13438\,
            PACKAGEPIN => \ioFifoData_wire\(7)
        );

    \ioFifoData_obuft_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13440\,
            PADOUT => \N__13439\,
            PADIN => \N__13438\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8751\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \iRxF_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13431\,
            DIN => \N__13430\,
            DOUT => \N__13429\,
            PACKAGEPIN => \iRxF_n_wire\
        );

    \iRxF_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13431\,
            PADOUT => \N__13430\,
            PADIN => \N__13429\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \iRxF_n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13422\,
            DIN => \N__13421\,
            DOUT => \N__13420\,
            PACKAGEPIN => \P1A3_wire\
        );

    \P1A3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13422\,
            PADOUT => \N__13421\,
            PADIN => \N__13420\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7546\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A7_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13413\,
            DIN => \N__13412\,
            DOUT => \N__13411\,
            PACKAGEPIN => \P1A7_wire\
        );

    \P1A7_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13413\,
            PADOUT => \N__13412\,
            PADIN => \N__13411\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9461\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BTN_N_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13404\,
            DIN => \N__13403\,
            DOUT => \N__13402\,
            PACKAGEPIN => \BTN_N_wire\
        );

    \BTN_N_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13404\,
            PADOUT => \N__13403\,
            PADIN => \N__13402\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \BTN_N_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13395\,
            DIN => \N__13394\,
            DOUT => \N__13393\,
            PACKAGEPIN => \ioFifoData_wire\(3)
        );

    \ioFifoData_obuft_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13395\,
            PADOUT => \N__13394\,
            PADIN => \N__13393\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8752\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13386\,
            DIN => \N__13385\,
            DOUT => \N__13384\,
            PACKAGEPIN => \ioFifoData_wire\(6)
        );

    \ioFifoData_obuft_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13386\,
            PADOUT => \N__13385\,
            PADIN => \N__13384\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8750\,
            DIN0 => OPEN,
            DOUT0 => \N__12840\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13377\,
            DIN => \N__13376\,
            DOUT => \N__13375\,
            PACKAGEPIN => \ioFifoData_wire\(5)
        );

    \ioFifoData_obuft_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13377\,
            PADOUT => \N__13376\,
            PADIN => \N__13375\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8728\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \oTx_n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13368\,
            DIN => \N__13367\,
            DOUT => \N__13366\,
            PACKAGEPIN => \oTx_n_wire\
        );

    \oTx_n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13368\,
            PADOUT => \N__13367\,
            PADIN => \N__13366\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8804\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \iTxE_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13359\,
            DIN => \N__13358\,
            DOUT => \N__13357\,
            PACKAGEPIN => \iTxE_n_wire\
        );

    \iTxE_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13359\,
            PADOUT => \N__13358\,
            PADIN => \N__13357\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \iTxE_n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13350\,
            DIN => \N__13349\,
            DOUT => \N__13348\,
            PACKAGEPIN => \ioFifoData_wire\(2)
        );

    \ioFifoData_obuft_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13350\,
            PADOUT => \N__13349\,
            PADIN => \N__13348\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8753\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13341\,
            DIN => \N__13340\,
            DOUT => \N__13339\,
            PACKAGEPIN => \P1A1_wire\
        );

    \P1A1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13341\,
            PADOUT => \N__13340\,
            PADIN => \N__13339\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \P1A1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__3179\ : InMux
    port map (
            O => \N__13322\,
            I => \N__13316\
        );

    \I__3178\ : InMux
    port map (
            O => \N__13321\,
            I => \N__13313\
        );

    \I__3177\ : InMux
    port map (
            O => \N__13320\,
            I => \N__13310\
        );

    \I__3176\ : InMux
    port map (
            O => \N__13319\,
            I => \N__13307\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__13316\,
            I => \N__13302\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__13313\,
            I => \N__13302\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__13310\,
            I => \N__13299\
        );

    \I__3172\ : LocalMux
    port map (
            O => \N__13307\,
            I => \N__13296\
        );

    \I__3171\ : Span4Mux_v
    port map (
            O => \N__13302\,
            I => \N__13293\
        );

    \I__3170\ : Span4Mux_v
    port map (
            O => \N__13299\,
            I => \N__13288\
        );

    \I__3169\ : Span4Mux_v
    port map (
            O => \N__13296\,
            I => \N__13288\
        );

    \I__3168\ : Odrv4
    port map (
            O => \N__13293\,
            I => \rTxByteZ0Z_7\
        );

    \I__3167\ : Odrv4
    port map (
            O => \N__13288\,
            I => \rTxByteZ0Z_7\
        );

    \I__3166\ : InMux
    port map (
            O => \N__13283\,
            I => \N__13280\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__13280\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_7\
        );

    \I__3164\ : InMux
    port map (
            O => \N__13277\,
            I => \N__13271\
        );

    \I__3163\ : InMux
    port map (
            O => \N__13276\,
            I => \N__13268\
        );

    \I__3162\ : InMux
    port map (
            O => \N__13275\,
            I => \N__13265\
        );

    \I__3161\ : InMux
    port map (
            O => \N__13274\,
            I => \N__13262\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__13271\,
            I => \N__13259\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__13268\,
            I => \N__13254\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__13265\,
            I => \N__13254\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__13262\,
            I => \N__13251\
        );

    \I__3156\ : Span4Mux_v
    port map (
            O => \N__13259\,
            I => \N__13248\
        );

    \I__3155\ : Span4Mux_v
    port map (
            O => \N__13254\,
            I => \N__13245\
        );

    \I__3154\ : Span4Mux_h
    port map (
            O => \N__13251\,
            I => \N__13242\
        );

    \I__3153\ : Odrv4
    port map (
            O => \N__13248\,
            I => \rTxByteZ0Z_1\
        );

    \I__3152\ : Odrv4
    port map (
            O => \N__13245\,
            I => \rTxByteZ0Z_1\
        );

    \I__3151\ : Odrv4
    port map (
            O => \N__13242\,
            I => \rTxByteZ0Z_1\
        );

    \I__3150\ : InMux
    port map (
            O => \N__13235\,
            I => \N__13232\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__13232\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_1\
        );

    \I__3148\ : InMux
    port map (
            O => \N__13229\,
            I => \N__13225\
        );

    \I__3147\ : InMux
    port map (
            O => \N__13228\,
            I => \N__13222\
        );

    \I__3146\ : LocalMux
    port map (
            O => \N__13225\,
            I => \N__13217\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__13222\,
            I => \N__13217\
        );

    \I__3144\ : Span4Mux_v
    port map (
            O => \N__13217\,
            I => \N__13213\
        );

    \I__3143\ : InMux
    port map (
            O => \N__13216\,
            I => \N__13210\
        );

    \I__3142\ : Sp12to4
    port map (
            O => \N__13213\,
            I => \N__13204\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__13210\,
            I => \N__13204\
        );

    \I__3140\ : InMux
    port map (
            O => \N__13209\,
            I => \N__13201\
        );

    \I__3139\ : Odrv12
    port map (
            O => \N__13204\,
            I => \rTxByteZ0Z_6\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__13201\,
            I => \rTxByteZ0Z_6\
        );

    \I__3137\ : InMux
    port map (
            O => \N__13196\,
            I => \N__13193\
        );

    \I__3136\ : LocalMux
    port map (
            O => \N__13193\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_6\
        );

    \I__3135\ : CEMux
    port map (
            O => \N__13190\,
            I => \N__13184\
        );

    \I__3134\ : CEMux
    port map (
            O => \N__13189\,
            I => \N__13181\
        );

    \I__3133\ : CEMux
    port map (
            O => \N__13188\,
            I => \N__13178\
        );

    \I__3132\ : CEMux
    port map (
            O => \N__13187\,
            I => \N__13175\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__13184\,
            I => \N__13172\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__13181\,
            I => \N__13169\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__13178\,
            I => \N__13164\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__13175\,
            I => \N__13164\
        );

    \I__3127\ : Span4Mux_h
    port map (
            O => \N__13172\,
            I => \N__13161\
        );

    \I__3126\ : Span4Mux_v
    port map (
            O => \N__13169\,
            I => \N__13158\
        );

    \I__3125\ : Span4Mux_v
    port map (
            O => \N__13164\,
            I => \N__13153\
        );

    \I__3124\ : Span4Mux_h
    port map (
            O => \N__13161\,
            I => \N__13153\
        );

    \I__3123\ : Odrv4
    port map (
            O => \N__13158\,
            I => \DUT.fifo_tx_inst.rFifoData_awe0\
        );

    \I__3122\ : Odrv4
    port map (
            O => \N__13153\,
            I => \DUT.fifo_tx_inst.rFifoData_awe0\
        );

    \I__3121\ : InMux
    port map (
            O => \N__13148\,
            I => \N__13144\
        );

    \I__3120\ : InMux
    port map (
            O => \N__13147\,
            I => \N__13141\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__13144\,
            I => \N__13137\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__13141\,
            I => \N__13134\
        );

    \I__3117\ : InMux
    port map (
            O => \N__13140\,
            I => \N__13131\
        );

    \I__3116\ : Span4Mux_v
    port map (
            O => \N__13137\,
            I => \N__13123\
        );

    \I__3115\ : Span4Mux_v
    port map (
            O => \N__13134\,
            I => \N__13123\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__13131\,
            I => \N__13123\
        );

    \I__3113\ : InMux
    port map (
            O => \N__13130\,
            I => \N__13120\
        );

    \I__3112\ : Odrv4
    port map (
            O => \N__13123\,
            I => \rTxByteZ0Z_5\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__13120\,
            I => \rTxByteZ0Z_5\
        );

    \I__3110\ : InMux
    port map (
            O => \N__13115\,
            I => \N__13112\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__13112\,
            I => \N__13109\
        );

    \I__3108\ : Odrv4
    port map (
            O => \N__13109\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_5\
        );

    \I__3107\ : InMux
    port map (
            O => \N__13106\,
            I => \N__13102\
        );

    \I__3106\ : InMux
    port map (
            O => \N__13105\,
            I => \N__13099\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__13102\,
            I => \N__13095\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__13099\,
            I => \N__13092\
        );

    \I__3103\ : InMux
    port map (
            O => \N__13098\,
            I => \N__13089\
        );

    \I__3102\ : Span4Mux_v
    port map (
            O => \N__13095\,
            I => \N__13081\
        );

    \I__3101\ : Span4Mux_h
    port map (
            O => \N__13092\,
            I => \N__13081\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__13089\,
            I => \N__13081\
        );

    \I__3099\ : InMux
    port map (
            O => \N__13088\,
            I => \N__13078\
        );

    \I__3098\ : Span4Mux_h
    port map (
            O => \N__13081\,
            I => \N__13075\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__13078\,
            I => \N__13072\
        );

    \I__3096\ : Odrv4
    port map (
            O => \N__13075\,
            I => \rTxByteZ0Z_0\
        );

    \I__3095\ : Odrv4
    port map (
            O => \N__13072\,
            I => \rTxByteZ0Z_0\
        );

    \I__3094\ : CascadeMux
    port map (
            O => \N__13067\,
            I => \N__13064\
        );

    \I__3093\ : InMux
    port map (
            O => \N__13064\,
            I => \N__13061\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__13061\,
            I => \N__13058\
        );

    \I__3091\ : Odrv4
    port map (
            O => \N__13058\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_0\
        );

    \I__3090\ : ClkMux
    port map (
            O => \N__13055\,
            I => \N__12887\
        );

    \I__3089\ : ClkMux
    port map (
            O => \N__13054\,
            I => \N__12887\
        );

    \I__3088\ : ClkMux
    port map (
            O => \N__13053\,
            I => \N__12887\
        );

    \I__3087\ : ClkMux
    port map (
            O => \N__13052\,
            I => \N__12887\
        );

    \I__3086\ : ClkMux
    port map (
            O => \N__13051\,
            I => \N__12887\
        );

    \I__3085\ : ClkMux
    port map (
            O => \N__13050\,
            I => \N__12887\
        );

    \I__3084\ : ClkMux
    port map (
            O => \N__13049\,
            I => \N__12887\
        );

    \I__3083\ : ClkMux
    port map (
            O => \N__13048\,
            I => \N__12887\
        );

    \I__3082\ : ClkMux
    port map (
            O => \N__13047\,
            I => \N__12887\
        );

    \I__3081\ : ClkMux
    port map (
            O => \N__13046\,
            I => \N__12887\
        );

    \I__3080\ : ClkMux
    port map (
            O => \N__13045\,
            I => \N__12887\
        );

    \I__3079\ : ClkMux
    port map (
            O => \N__13044\,
            I => \N__12887\
        );

    \I__3078\ : ClkMux
    port map (
            O => \N__13043\,
            I => \N__12887\
        );

    \I__3077\ : ClkMux
    port map (
            O => \N__13042\,
            I => \N__12887\
        );

    \I__3076\ : ClkMux
    port map (
            O => \N__13041\,
            I => \N__12887\
        );

    \I__3075\ : ClkMux
    port map (
            O => \N__13040\,
            I => \N__12887\
        );

    \I__3074\ : ClkMux
    port map (
            O => \N__13039\,
            I => \N__12887\
        );

    \I__3073\ : ClkMux
    port map (
            O => \N__13038\,
            I => \N__12887\
        );

    \I__3072\ : ClkMux
    port map (
            O => \N__13037\,
            I => \N__12887\
        );

    \I__3071\ : ClkMux
    port map (
            O => \N__13036\,
            I => \N__12887\
        );

    \I__3070\ : ClkMux
    port map (
            O => \N__13035\,
            I => \N__12887\
        );

    \I__3069\ : ClkMux
    port map (
            O => \N__13034\,
            I => \N__12887\
        );

    \I__3068\ : ClkMux
    port map (
            O => \N__13033\,
            I => \N__12887\
        );

    \I__3067\ : ClkMux
    port map (
            O => \N__13032\,
            I => \N__12887\
        );

    \I__3066\ : ClkMux
    port map (
            O => \N__13031\,
            I => \N__12887\
        );

    \I__3065\ : ClkMux
    port map (
            O => \N__13030\,
            I => \N__12887\
        );

    \I__3064\ : ClkMux
    port map (
            O => \N__13029\,
            I => \N__12887\
        );

    \I__3063\ : ClkMux
    port map (
            O => \N__13028\,
            I => \N__12887\
        );

    \I__3062\ : ClkMux
    port map (
            O => \N__13027\,
            I => \N__12887\
        );

    \I__3061\ : ClkMux
    port map (
            O => \N__13026\,
            I => \N__12887\
        );

    \I__3060\ : ClkMux
    port map (
            O => \N__13025\,
            I => \N__12887\
        );

    \I__3059\ : ClkMux
    port map (
            O => \N__13024\,
            I => \N__12887\
        );

    \I__3058\ : ClkMux
    port map (
            O => \N__13023\,
            I => \N__12887\
        );

    \I__3057\ : ClkMux
    port map (
            O => \N__13022\,
            I => \N__12887\
        );

    \I__3056\ : ClkMux
    port map (
            O => \N__13021\,
            I => \N__12887\
        );

    \I__3055\ : ClkMux
    port map (
            O => \N__13020\,
            I => \N__12887\
        );

    \I__3054\ : ClkMux
    port map (
            O => \N__13019\,
            I => \N__12887\
        );

    \I__3053\ : ClkMux
    port map (
            O => \N__13018\,
            I => \N__12887\
        );

    \I__3052\ : ClkMux
    port map (
            O => \N__13017\,
            I => \N__12887\
        );

    \I__3051\ : ClkMux
    port map (
            O => \N__13016\,
            I => \N__12887\
        );

    \I__3050\ : ClkMux
    port map (
            O => \N__13015\,
            I => \N__12887\
        );

    \I__3049\ : ClkMux
    port map (
            O => \N__13014\,
            I => \N__12887\
        );

    \I__3048\ : ClkMux
    port map (
            O => \N__13013\,
            I => \N__12887\
        );

    \I__3047\ : ClkMux
    port map (
            O => \N__13012\,
            I => \N__12887\
        );

    \I__3046\ : ClkMux
    port map (
            O => \N__13011\,
            I => \N__12887\
        );

    \I__3045\ : ClkMux
    port map (
            O => \N__13010\,
            I => \N__12887\
        );

    \I__3044\ : ClkMux
    port map (
            O => \N__13009\,
            I => \N__12887\
        );

    \I__3043\ : ClkMux
    port map (
            O => \N__13008\,
            I => \N__12887\
        );

    \I__3042\ : ClkMux
    port map (
            O => \N__13007\,
            I => \N__12887\
        );

    \I__3041\ : ClkMux
    port map (
            O => \N__13006\,
            I => \N__12887\
        );

    \I__3040\ : ClkMux
    port map (
            O => \N__13005\,
            I => \N__12887\
        );

    \I__3039\ : ClkMux
    port map (
            O => \N__13004\,
            I => \N__12887\
        );

    \I__3038\ : ClkMux
    port map (
            O => \N__13003\,
            I => \N__12887\
        );

    \I__3037\ : ClkMux
    port map (
            O => \N__13002\,
            I => \N__12887\
        );

    \I__3036\ : ClkMux
    port map (
            O => \N__13001\,
            I => \N__12887\
        );

    \I__3035\ : ClkMux
    port map (
            O => \N__13000\,
            I => \N__12887\
        );

    \I__3034\ : GlobalMux
    port map (
            O => \N__12887\,
            I => clk_48mhz
        );

    \I__3033\ : CEMux
    port map (
            O => \N__12884\,
            I => \N__12880\
        );

    \I__3032\ : CEMux
    port map (
            O => \N__12883\,
            I => \N__12876\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__12880\,
            I => \N__12873\
        );

    \I__3030\ : CEMux
    port map (
            O => \N__12879\,
            I => \N__12870\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__12876\,
            I => \N__12867\
        );

    \I__3028\ : Span4Mux_v
    port map (
            O => \N__12873\,
            I => \N__12862\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__12870\,
            I => \N__12862\
        );

    \I__3026\ : Span4Mux_h
    port map (
            O => \N__12867\,
            I => \N__12856\
        );

    \I__3025\ : Span4Mux_v
    port map (
            O => \N__12862\,
            I => \N__12856\
        );

    \I__3024\ : InMux
    port map (
            O => \N__12861\,
            I => \N__12853\
        );

    \I__3023\ : Odrv4
    port map (
            O => \N__12856\,
            I => \DUT.fifo_tx_inst.rFifoData_awe1\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__12853\,
            I => \DUT.fifo_tx_inst.rFifoData_awe1\
        );

    \I__3021\ : CascadeMux
    port map (
            O => \N__12848\,
            I => \N__12837\
        );

    \I__3020\ : CascadeMux
    port map (
            O => \N__12847\,
            I => \N__12834\
        );

    \I__3019\ : CascadeMux
    port map (
            O => \N__12846\,
            I => \N__12831\
        );

    \I__3018\ : CascadeMux
    port map (
            O => \N__12845\,
            I => \N__12828\
        );

    \I__3017\ : CascadeMux
    port map (
            O => \N__12844\,
            I => \N__12825\
        );

    \I__3016\ : CascadeMux
    port map (
            O => \N__12843\,
            I => \N__12822\
        );

    \I__3015\ : CascadeMux
    port map (
            O => \N__12842\,
            I => \N__12819\
        );

    \I__3014\ : IoInMux
    port map (
            O => \N__12841\,
            I => \N__12808\
        );

    \I__3013\ : IoInMux
    port map (
            O => \N__12840\,
            I => \N__12804\
        );

    \I__3012\ : InMux
    port map (
            O => \N__12837\,
            I => \N__12797\
        );

    \I__3011\ : InMux
    port map (
            O => \N__12834\,
            I => \N__12797\
        );

    \I__3010\ : InMux
    port map (
            O => \N__12831\,
            I => \N__12797\
        );

    \I__3009\ : InMux
    port map (
            O => \N__12828\,
            I => \N__12788\
        );

    \I__3008\ : InMux
    port map (
            O => \N__12825\,
            I => \N__12788\
        );

    \I__3007\ : InMux
    port map (
            O => \N__12822\,
            I => \N__12788\
        );

    \I__3006\ : InMux
    port map (
            O => \N__12819\,
            I => \N__12788\
        );

    \I__3005\ : CascadeMux
    port map (
            O => \N__12818\,
            I => \N__12785\
        );

    \I__3004\ : CascadeMux
    port map (
            O => \N__12817\,
            I => \N__12782\
        );

    \I__3003\ : CascadeMux
    port map (
            O => \N__12816\,
            I => \N__12779\
        );

    \I__3002\ : CascadeMux
    port map (
            O => \N__12815\,
            I => \N__12776\
        );

    \I__3001\ : CascadeMux
    port map (
            O => \N__12814\,
            I => \N__12773\
        );

    \I__3000\ : CascadeMux
    port map (
            O => \N__12813\,
            I => \N__12770\
        );

    \I__2999\ : CascadeMux
    port map (
            O => \N__12812\,
            I => \N__12767\
        );

    \I__2998\ : CascadeMux
    port map (
            O => \N__12811\,
            I => \N__12764\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__12808\,
            I => \N__12753\
        );

    \I__2996\ : CascadeMux
    port map (
            O => \N__12807\,
            I => \N__12748\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__12804\,
            I => \N__12744\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__12797\,
            I => \N__12736\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__12788\,
            I => \N__12736\
        );

    \I__2992\ : InMux
    port map (
            O => \N__12785\,
            I => \N__12727\
        );

    \I__2991\ : InMux
    port map (
            O => \N__12782\,
            I => \N__12727\
        );

    \I__2990\ : InMux
    port map (
            O => \N__12779\,
            I => \N__12727\
        );

    \I__2989\ : InMux
    port map (
            O => \N__12776\,
            I => \N__12727\
        );

    \I__2988\ : InMux
    port map (
            O => \N__12773\,
            I => \N__12718\
        );

    \I__2987\ : InMux
    port map (
            O => \N__12770\,
            I => \N__12718\
        );

    \I__2986\ : InMux
    port map (
            O => \N__12767\,
            I => \N__12718\
        );

    \I__2985\ : InMux
    port map (
            O => \N__12764\,
            I => \N__12718\
        );

    \I__2984\ : CascadeMux
    port map (
            O => \N__12763\,
            I => \N__12715\
        );

    \I__2983\ : CascadeMux
    port map (
            O => \N__12762\,
            I => \N__12712\
        );

    \I__2982\ : CascadeMux
    port map (
            O => \N__12761\,
            I => \N__12709\
        );

    \I__2981\ : CascadeMux
    port map (
            O => \N__12760\,
            I => \N__12706\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__12759\,
            I => \N__12703\
        );

    \I__2979\ : CascadeMux
    port map (
            O => \N__12758\,
            I => \N__12699\
        );

    \I__2978\ : CascadeMux
    port map (
            O => \N__12757\,
            I => \N__12696\
        );

    \I__2977\ : CascadeMux
    port map (
            O => \N__12756\,
            I => \N__12692\
        );

    \I__2976\ : IoSpan4Mux
    port map (
            O => \N__12753\,
            I => \N__12689\
        );

    \I__2975\ : InMux
    port map (
            O => \N__12752\,
            I => \N__12686\
        );

    \I__2974\ : InMux
    port map (
            O => \N__12751\,
            I => \N__12679\
        );

    \I__2973\ : InMux
    port map (
            O => \N__12748\,
            I => \N__12679\
        );

    \I__2972\ : InMux
    port map (
            O => \N__12747\,
            I => \N__12679\
        );

    \I__2971\ : Span4Mux_s0_v
    port map (
            O => \N__12744\,
            I => \N__12676\
        );

    \I__2970\ : CascadeMux
    port map (
            O => \N__12743\,
            I => \N__12673\
        );

    \I__2969\ : CascadeMux
    port map (
            O => \N__12742\,
            I => \N__12670\
        );

    \I__2968\ : CascadeMux
    port map (
            O => \N__12741\,
            I => \N__12667\
        );

    \I__2967\ : Span4Mux_v
    port map (
            O => \N__12736\,
            I => \N__12660\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__12727\,
            I => \N__12660\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__12718\,
            I => \N__12660\
        );

    \I__2964\ : InMux
    port map (
            O => \N__12715\,
            I => \N__12657\
        );

    \I__2963\ : InMux
    port map (
            O => \N__12712\,
            I => \N__12648\
        );

    \I__2962\ : InMux
    port map (
            O => \N__12709\,
            I => \N__12648\
        );

    \I__2961\ : InMux
    port map (
            O => \N__12706\,
            I => \N__12648\
        );

    \I__2960\ : InMux
    port map (
            O => \N__12703\,
            I => \N__12648\
        );

    \I__2959\ : InMux
    port map (
            O => \N__12702\,
            I => \N__12637\
        );

    \I__2958\ : InMux
    port map (
            O => \N__12699\,
            I => \N__12637\
        );

    \I__2957\ : InMux
    port map (
            O => \N__12696\,
            I => \N__12637\
        );

    \I__2956\ : InMux
    port map (
            O => \N__12695\,
            I => \N__12637\
        );

    \I__2955\ : InMux
    port map (
            O => \N__12692\,
            I => \N__12637\
        );

    \I__2954\ : Span4Mux_s2_v
    port map (
            O => \N__12689\,
            I => \N__12633\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__12686\,
            I => \N__12628\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__12679\,
            I => \N__12628\
        );

    \I__2951\ : Span4Mux_h
    port map (
            O => \N__12676\,
            I => \N__12625\
        );

    \I__2950\ : InMux
    port map (
            O => \N__12673\,
            I => \N__12618\
        );

    \I__2949\ : InMux
    port map (
            O => \N__12670\,
            I => \N__12618\
        );

    \I__2948\ : InMux
    port map (
            O => \N__12667\,
            I => \N__12618\
        );

    \I__2947\ : Span4Mux_h
    port map (
            O => \N__12660\,
            I => \N__12611\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__12657\,
            I => \N__12611\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__12648\,
            I => \N__12611\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__12637\,
            I => \N__12608\
        );

    \I__2943\ : InMux
    port map (
            O => \N__12636\,
            I => \N__12605\
        );

    \I__2942\ : Sp12to4
    port map (
            O => \N__12633\,
            I => \N__12602\
        );

    \I__2941\ : Sp12to4
    port map (
            O => \N__12628\,
            I => \N__12599\
        );

    \I__2940\ : Span4Mux_v
    port map (
            O => \N__12625\,
            I => \N__12596\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__12618\,
            I => \N__12587\
        );

    \I__2938\ : Span4Mux_v
    port map (
            O => \N__12611\,
            I => \N__12587\
        );

    \I__2937\ : Span4Mux_v
    port map (
            O => \N__12608\,
            I => \N__12587\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__12605\,
            I => \N__12587\
        );

    \I__2935\ : Span12Mux_s10_v
    port map (
            O => \N__12602\,
            I => \N__12584\
        );

    \I__2934\ : Span12Mux_v
    port map (
            O => \N__12599\,
            I => \N__12581\
        );

    \I__2933\ : Span4Mux_v
    port map (
            O => \N__12596\,
            I => \N__12576\
        );

    \I__2932\ : Span4Mux_h
    port map (
            O => \N__12587\,
            I => \N__12576\
        );

    \I__2931\ : Odrv12
    port map (
            O => \N__12584\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2930\ : Odrv12
    port map (
            O => \N__12581\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2929\ : Odrv4
    port map (
            O => \N__12576\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2928\ : InMux
    port map (
            O => \N__12569\,
            I => \N__12566\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__12566\,
            I => \N__12563\
        );

    \I__2926\ : Span4Mux_h
    port map (
            O => \N__12563\,
            I => \N__12560\
        );

    \I__2925\ : Odrv4
    port map (
            O => \N__12560\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_4\
        );

    \I__2924\ : InMux
    port map (
            O => \N__12557\,
            I => \N__12554\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__12554\,
            I => \N__12551\
        );

    \I__2922\ : Span4Mux_h
    port map (
            O => \N__12551\,
            I => \N__12548\
        );

    \I__2921\ : Odrv4
    port map (
            O => \N__12548\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_5\
        );

    \I__2920\ : InMux
    port map (
            O => \N__12545\,
            I => \N__12542\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__12542\,
            I => \N__12539\
        );

    \I__2918\ : Span4Mux_h
    port map (
            O => \N__12539\,
            I => \N__12536\
        );

    \I__2917\ : Odrv4
    port map (
            O => \N__12536\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_6\
        );

    \I__2916\ : InMux
    port map (
            O => \N__12533\,
            I => \N__12530\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__12530\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_7\
        );

    \I__2914\ : CEMux
    port map (
            O => \N__12527\,
            I => \N__12524\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__12524\,
            I => \N__12520\
        );

    \I__2912\ : InMux
    port map (
            O => \N__12523\,
            I => \N__12517\
        );

    \I__2911\ : Span4Mux_v
    port map (
            O => \N__12520\,
            I => \N__12514\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__12517\,
            I => \N__12511\
        );

    \I__2909\ : Odrv4
    port map (
            O => \N__12514\,
            I => \DUT.fifo_tx_inst.rFifoData_awe3\
        );

    \I__2908\ : Odrv12
    port map (
            O => \N__12511\,
            I => \DUT.fifo_tx_inst.rFifoData_awe3\
        );

    \I__2907\ : InMux
    port map (
            O => \N__12506\,
            I => \N__12503\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__12503\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_1\
        );

    \I__2905\ : InMux
    port map (
            O => \N__12500\,
            I => \N__12494\
        );

    \I__2904\ : InMux
    port map (
            O => \N__12499\,
            I => \N__12491\
        );

    \I__2903\ : InMux
    port map (
            O => \N__12498\,
            I => \N__12488\
        );

    \I__2902\ : InMux
    port map (
            O => \N__12497\,
            I => \N__12485\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__12494\,
            I => \N__12480\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__12491\,
            I => \N__12480\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__12488\,
            I => \N__12477\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__12485\,
            I => \N__12474\
        );

    \I__2897\ : Span4Mux_h
    port map (
            O => \N__12480\,
            I => \N__12471\
        );

    \I__2896\ : Span4Mux_h
    port map (
            O => \N__12477\,
            I => \N__12466\
        );

    \I__2895\ : Span4Mux_h
    port map (
            O => \N__12474\,
            I => \N__12466\
        );

    \I__2894\ : Odrv4
    port map (
            O => \N__12471\,
            I => \rTxByteZ0Z_2\
        );

    \I__2893\ : Odrv4
    port map (
            O => \N__12466\,
            I => \rTxByteZ0Z_2\
        );

    \I__2892\ : CascadeMux
    port map (
            O => \N__12461\,
            I => \N__12458\
        );

    \I__2891\ : InMux
    port map (
            O => \N__12458\,
            I => \N__12455\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__12455\,
            I => \N__12452\
        );

    \I__2889\ : Span4Mux_h
    port map (
            O => \N__12452\,
            I => \N__12449\
        );

    \I__2888\ : Odrv4
    port map (
            O => \N__12449\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_2\
        );

    \I__2887\ : InMux
    port map (
            O => \N__12446\,
            I => \N__12442\
        );

    \I__2886\ : InMux
    port map (
            O => \N__12445\,
            I => \N__12439\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__12442\,
            I => \N__12435\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__12439\,
            I => \N__12432\
        );

    \I__2883\ : InMux
    port map (
            O => \N__12438\,
            I => \N__12429\
        );

    \I__2882\ : Span4Mux_h
    port map (
            O => \N__12435\,
            I => \N__12422\
        );

    \I__2881\ : Span4Mux_v
    port map (
            O => \N__12432\,
            I => \N__12422\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__12429\,
            I => \N__12422\
        );

    \I__2879\ : Span4Mux_h
    port map (
            O => \N__12422\,
            I => \N__12418\
        );

    \I__2878\ : InMux
    port map (
            O => \N__12421\,
            I => \N__12415\
        );

    \I__2877\ : Odrv4
    port map (
            O => \N__12418\,
            I => \rTxByteZ0Z_3\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__12415\,
            I => \rTxByteZ0Z_3\
        );

    \I__2875\ : InMux
    port map (
            O => \N__12410\,
            I => \N__12407\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__12407\,
            I => \N__12404\
        );

    \I__2873\ : Span4Mux_h
    port map (
            O => \N__12404\,
            I => \N__12401\
        );

    \I__2872\ : Odrv4
    port map (
            O => \N__12401\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_3\
        );

    \I__2871\ : InMux
    port map (
            O => \N__12398\,
            I => \N__12394\
        );

    \I__2870\ : InMux
    port map (
            O => \N__12397\,
            I => \N__12391\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__12394\,
            I => \N__12385\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__12391\,
            I => \N__12385\
        );

    \I__2867\ : InMux
    port map (
            O => \N__12390\,
            I => \N__12382\
        );

    \I__2866\ : Span4Mux_v
    port map (
            O => \N__12385\,
            I => \N__12376\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__12382\,
            I => \N__12376\
        );

    \I__2864\ : InMux
    port map (
            O => \N__12381\,
            I => \N__12373\
        );

    \I__2863\ : Odrv4
    port map (
            O => \N__12376\,
            I => \rTxByteZ0Z_4\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__12373\,
            I => \rTxByteZ0Z_4\
        );

    \I__2861\ : CascadeMux
    port map (
            O => \N__12368\,
            I => \N__12365\
        );

    \I__2860\ : InMux
    port map (
            O => \N__12365\,
            I => \N__12362\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__12362\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_4\
        );

    \I__2858\ : CascadeMux
    port map (
            O => \N__12359\,
            I => \N__12356\
        );

    \I__2857\ : InMux
    port map (
            O => \N__12356\,
            I => \N__12353\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__12353\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_6\
        );

    \I__2855\ : InMux
    port map (
            O => \N__12350\,
            I => \N__12346\
        );

    \I__2854\ : InMux
    port map (
            O => \N__12349\,
            I => \N__12343\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__12346\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_2\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__12343\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_2\
        );

    \I__2851\ : InMux
    port map (
            O => \N__12338\,
            I => \N__12334\
        );

    \I__2850\ : InMux
    port map (
            O => \N__12337\,
            I => \N__12331\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__12334\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_4\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__12331\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_4\
        );

    \I__2847\ : CascadeMux
    port map (
            O => \N__12326\,
            I => \N__12322\
        );

    \I__2846\ : InMux
    port map (
            O => \N__12325\,
            I => \N__12319\
        );

    \I__2845\ : InMux
    port map (
            O => \N__12322\,
            I => \N__12316\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__12319\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_5\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__12316\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_5\
        );

    \I__2842\ : InMux
    port map (
            O => \N__12311\,
            I => \N__12307\
        );

    \I__2841\ : InMux
    port map (
            O => \N__12310\,
            I => \N__12304\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__12307\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_3\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__12304\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_3\
        );

    \I__2838\ : InMux
    port map (
            O => \N__12299\,
            I => \N__12295\
        );

    \I__2837\ : InMux
    port map (
            O => \N__12298\,
            I => \N__12292\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__12295\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_12\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__12292\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_12\
        );

    \I__2834\ : InMux
    port map (
            O => \N__12287\,
            I => \N__12283\
        );

    \I__2833\ : InMux
    port map (
            O => \N__12286\,
            I => \N__12280\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__12283\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_7\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__12280\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_7\
        );

    \I__2830\ : CascadeMux
    port map (
            O => \N__12275\,
            I => \N__12271\
        );

    \I__2829\ : InMux
    port map (
            O => \N__12274\,
            I => \N__12268\
        );

    \I__2828\ : InMux
    port map (
            O => \N__12271\,
            I => \N__12265\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__12268\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_13\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__12265\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_13\
        );

    \I__2825\ : InMux
    port map (
            O => \N__12260\,
            I => \N__12256\
        );

    \I__2824\ : InMux
    port map (
            O => \N__12259\,
            I => \N__12253\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__12256\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_6\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__12253\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_6\
        );

    \I__2821\ : InMux
    port map (
            O => \N__12248\,
            I => \N__12245\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__12245\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_9\
        );

    \I__2819\ : InMux
    port map (
            O => \N__12242\,
            I => \N__12239\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__12239\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_7\
        );

    \I__2817\ : CascadeMux
    port map (
            O => \N__12236\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_8_cascade_\
        );

    \I__2816\ : InMux
    port map (
            O => \N__12233\,
            I => \N__12230\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__12230\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_6\
        );

    \I__2814\ : InMux
    port map (
            O => \N__12227\,
            I => \N__12218\
        );

    \I__2813\ : InMux
    port map (
            O => \N__12226\,
            I => \N__12208\
        );

    \I__2812\ : InMux
    port map (
            O => \N__12225\,
            I => \N__12208\
        );

    \I__2811\ : InMux
    port map (
            O => \N__12224\,
            I => \N__12208\
        );

    \I__2810\ : InMux
    port map (
            O => \N__12223\,
            I => \N__12205\
        );

    \I__2809\ : InMux
    port map (
            O => \N__12222\,
            I => \N__12200\
        );

    \I__2808\ : InMux
    port map (
            O => \N__12221\,
            I => \N__12200\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__12218\,
            I => \N__12196\
        );

    \I__2806\ : InMux
    port map (
            O => \N__12217\,
            I => \N__12189\
        );

    \I__2805\ : InMux
    port map (
            O => \N__12216\,
            I => \N__12189\
        );

    \I__2804\ : InMux
    port map (
            O => \N__12215\,
            I => \N__12189\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__12208\,
            I => \N__12182\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__12205\,
            I => \N__12182\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__12200\,
            I => \N__12182\
        );

    \I__2800\ : InMux
    port map (
            O => \N__12199\,
            I => \N__12179\
        );

    \I__2799\ : Odrv4
    port map (
            O => \N__12196\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__12189\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0\
        );

    \I__2797\ : Odrv4
    port map (
            O => \N__12182\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__12179\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0\
        );

    \I__2795\ : InMux
    port map (
            O => \N__12170\,
            I => \N__12159\
        );

    \I__2794\ : InMux
    port map (
            O => \N__12169\,
            I => \N__12159\
        );

    \I__2793\ : InMux
    port map (
            O => \N__12168\,
            I => \N__12159\
        );

    \I__2792\ : InMux
    port map (
            O => \N__12167\,
            I => \N__12148\
        );

    \I__2791\ : InMux
    port map (
            O => \N__12166\,
            I => \N__12148\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__12159\,
            I => \N__12145\
        );

    \I__2789\ : InMux
    port map (
            O => \N__12158\,
            I => \N__12142\
        );

    \I__2788\ : InMux
    port map (
            O => \N__12157\,
            I => \N__12137\
        );

    \I__2787\ : InMux
    port map (
            O => \N__12156\,
            I => \N__12137\
        );

    \I__2786\ : InMux
    port map (
            O => \N__12155\,
            I => \N__12130\
        );

    \I__2785\ : InMux
    port map (
            O => \N__12154\,
            I => \N__12130\
        );

    \I__2784\ : InMux
    port map (
            O => \N__12153\,
            I => \N__12130\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__12148\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__2782\ : Odrv4
    port map (
            O => \N__12145\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__12142\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__12137\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__12130\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__2778\ : CascadeMux
    port map (
            O => \N__12119\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0_cascade_\
        );

    \I__2777\ : InMux
    port map (
            O => \N__12116\,
            I => \N__12113\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__12113\,
            I => \N__12110\
        );

    \I__2775\ : Odrv12
    port map (
            O => \N__12110\,
            I => \DUT.uart_inst0.N_5_0\
        );

    \I__2774\ : InMux
    port map (
            O => \N__12107\,
            I => \N__12104\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__12104\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_0\
        );

    \I__2772\ : InMux
    port map (
            O => \N__12101\,
            I => \N__12098\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__12098\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_1\
        );

    \I__2770\ : InMux
    port map (
            O => \N__12095\,
            I => \N__12092\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__12092\,
            I => \N__12089\
        );

    \I__2768\ : Odrv4
    port map (
            O => \N__12089\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_2\
        );

    \I__2767\ : InMux
    port map (
            O => \N__12086\,
            I => \N__12083\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__12083\,
            I => \N__12080\
        );

    \I__2765\ : Odrv4
    port map (
            O => \N__12080\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_3\
        );

    \I__2764\ : CascadeMux
    port map (
            O => \N__12077\,
            I => \DUT.uart_inst0.g0_i_a3_0_cascade_\
        );

    \I__2763\ : CascadeMux
    port map (
            O => \N__12074\,
            I => \N__12067\
        );

    \I__2762\ : CascadeMux
    port map (
            O => \N__12073\,
            I => \N__12056\
        );

    \I__2761\ : InMux
    port map (
            O => \N__12072\,
            I => \N__12053\
        );

    \I__2760\ : InMux
    port map (
            O => \N__12071\,
            I => \N__12050\
        );

    \I__2759\ : InMux
    port map (
            O => \N__12070\,
            I => \N__12047\
        );

    \I__2758\ : InMux
    port map (
            O => \N__12067\,
            I => \N__12044\
        );

    \I__2757\ : InMux
    port map (
            O => \N__12066\,
            I => \N__12041\
        );

    \I__2756\ : InMux
    port map (
            O => \N__12065\,
            I => \N__12036\
        );

    \I__2755\ : InMux
    port map (
            O => \N__12064\,
            I => \N__12036\
        );

    \I__2754\ : InMux
    port map (
            O => \N__12063\,
            I => \N__12031\
        );

    \I__2753\ : InMux
    port map (
            O => \N__12062\,
            I => \N__12031\
        );

    \I__2752\ : InMux
    port map (
            O => \N__12061\,
            I => \N__12028\
        );

    \I__2751\ : InMux
    port map (
            O => \N__12060\,
            I => \N__12025\
        );

    \I__2750\ : InMux
    port map (
            O => \N__12059\,
            I => \N__12022\
        );

    \I__2749\ : InMux
    port map (
            O => \N__12056\,
            I => \N__12019\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__12053\,
            I => \N__12016\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__12050\,
            I => \N__12013\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__12047\,
            I => \N__12010\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__12044\,
            I => \N__12007\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__12041\,
            I => \N__12004\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__12036\,
            I => \N__12001\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__12031\,
            I => \N__11997\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__12028\,
            I => \N__11994\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__12025\,
            I => \N__11990\
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__12022\,
            I => \N__11986\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__12019\,
            I => \N__11982\
        );

    \I__2737\ : Glb2LocalMux
    port map (
            O => \N__12016\,
            I => \N__11930\
        );

    \I__2736\ : Glb2LocalMux
    port map (
            O => \N__12013\,
            I => \N__11930\
        );

    \I__2735\ : Glb2LocalMux
    port map (
            O => \N__12010\,
            I => \N__11930\
        );

    \I__2734\ : Glb2LocalMux
    port map (
            O => \N__12007\,
            I => \N__11930\
        );

    \I__2733\ : Glb2LocalMux
    port map (
            O => \N__12004\,
            I => \N__11930\
        );

    \I__2732\ : Glb2LocalMux
    port map (
            O => \N__12001\,
            I => \N__11930\
        );

    \I__2731\ : CEMux
    port map (
            O => \N__12000\,
            I => \N__11930\
        );

    \I__2730\ : Glb2LocalMux
    port map (
            O => \N__11997\,
            I => \N__11930\
        );

    \I__2729\ : Glb2LocalMux
    port map (
            O => \N__11994\,
            I => \N__11930\
        );

    \I__2728\ : CEMux
    port map (
            O => \N__11993\,
            I => \N__11930\
        );

    \I__2727\ : Glb2LocalMux
    port map (
            O => \N__11990\,
            I => \N__11930\
        );

    \I__2726\ : CEMux
    port map (
            O => \N__11989\,
            I => \N__11930\
        );

    \I__2725\ : Glb2LocalMux
    port map (
            O => \N__11986\,
            I => \N__11930\
        );

    \I__2724\ : CEMux
    port map (
            O => \N__11985\,
            I => \N__11930\
        );

    \I__2723\ : Glb2LocalMux
    port map (
            O => \N__11982\,
            I => \N__11930\
        );

    \I__2722\ : CEMux
    port map (
            O => \N__11981\,
            I => \N__11930\
        );

    \I__2721\ : CEMux
    port map (
            O => \N__11980\,
            I => \N__11930\
        );

    \I__2720\ : CEMux
    port map (
            O => \N__11979\,
            I => \N__11930\
        );

    \I__2719\ : CEMux
    port map (
            O => \N__11978\,
            I => \N__11930\
        );

    \I__2718\ : CEMux
    port map (
            O => \N__11977\,
            I => \N__11930\
        );

    \I__2717\ : CEMux
    port map (
            O => \N__11976\,
            I => \N__11930\
        );

    \I__2716\ : CEMux
    port map (
            O => \N__11975\,
            I => \N__11930\
        );

    \I__2715\ : GlobalMux
    port map (
            O => \N__11930\,
            I => \N__11927\
        );

    \I__2714\ : gio2CtrlBuf
    port map (
            O => \N__11927\,
            I => \wPllLocked_g\
        );

    \I__2713\ : InMux
    port map (
            O => \N__11924\,
            I => \N__11921\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__11921\,
            I => \N__11915\
        );

    \I__2711\ : CascadeMux
    port map (
            O => \N__11920\,
            I => \N__11912\
        );

    \I__2710\ : InMux
    port map (
            O => \N__11919\,
            I => \N__11907\
        );

    \I__2709\ : InMux
    port map (
            O => \N__11918\,
            I => \N__11904\
        );

    \I__2708\ : Span4Mux_h
    port map (
            O => \N__11915\,
            I => \N__11901\
        );

    \I__2707\ : InMux
    port map (
            O => \N__11912\,
            I => \N__11894\
        );

    \I__2706\ : InMux
    port map (
            O => \N__11911\,
            I => \N__11894\
        );

    \I__2705\ : InMux
    port map (
            O => \N__11910\,
            I => \N__11894\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__11907\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_4\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__11904\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_4\
        );

    \I__2702\ : Odrv4
    port map (
            O => \N__11901\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_4\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__11894\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_4\
        );

    \I__2700\ : InMux
    port map (
            O => \N__11885\,
            I => \N__11875\
        );

    \I__2699\ : InMux
    port map (
            O => \N__11884\,
            I => \N__11872\
        );

    \I__2698\ : CascadeMux
    port map (
            O => \N__11883\,
            I => \N__11869\
        );

    \I__2697\ : InMux
    port map (
            O => \N__11882\,
            I => \N__11861\
        );

    \I__2696\ : InMux
    port map (
            O => \N__11881\,
            I => \N__11861\
        );

    \I__2695\ : InMux
    port map (
            O => \N__11880\,
            I => \N__11861\
        );

    \I__2694\ : InMux
    port map (
            O => \N__11879\,
            I => \N__11856\
        );

    \I__2693\ : InMux
    port map (
            O => \N__11878\,
            I => \N__11856\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__11875\,
            I => \N__11853\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__11872\,
            I => \N__11850\
        );

    \I__2690\ : InMux
    port map (
            O => \N__11869\,
            I => \N__11845\
        );

    \I__2689\ : InMux
    port map (
            O => \N__11868\,
            I => \N__11845\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__11861\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__11856\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__2686\ : Odrv4
    port map (
            O => \N__11853\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__2685\ : Odrv4
    port map (
            O => \N__11850\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__11845\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__2683\ : InMux
    port map (
            O => \N__11834\,
            I => \N__11830\
        );

    \I__2682\ : CascadeMux
    port map (
            O => \N__11833\,
            I => \N__11826\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__11830\,
            I => \N__11823\
        );

    \I__2680\ : CascadeMux
    port map (
            O => \N__11829\,
            I => \N__11818\
        );

    \I__2679\ : InMux
    port map (
            O => \N__11826\,
            I => \N__11815\
        );

    \I__2678\ : Span4Mux_h
    port map (
            O => \N__11823\,
            I => \N__11812\
        );

    \I__2677\ : InMux
    port map (
            O => \N__11822\,
            I => \N__11809\
        );

    \I__2676\ : InMux
    port map (
            O => \N__11821\,
            I => \N__11804\
        );

    \I__2675\ : InMux
    port map (
            O => \N__11818\,
            I => \N__11804\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__11815\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_5\
        );

    \I__2673\ : Odrv4
    port map (
            O => \N__11812\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_5\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__11809\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_5\
        );

    \I__2671\ : LocalMux
    port map (
            O => \N__11804\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_5\
        );

    \I__2670\ : InMux
    port map (
            O => \N__11795\,
            I => \N__11792\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__11792\,
            I => \DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0\
        );

    \I__2668\ : CascadeMux
    port map (
            O => \N__11789\,
            I => \DUT.uart_inst0.g0_11_a3_2_cascade_\
        );

    \I__2667\ : InMux
    port map (
            O => \N__11786\,
            I => \N__11783\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__11783\,
            I => \N__11780\
        );

    \I__2665\ : Odrv4
    port map (
            O => \N__11780\,
            I => \DUT.uart_inst0.N_7\
        );

    \I__2664\ : InMux
    port map (
            O => \N__11777\,
            I => \N__11774\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__11774\,
            I => \N__11769\
        );

    \I__2662\ : InMux
    port map (
            O => \N__11773\,
            I => \N__11760\
        );

    \I__2661\ : InMux
    port map (
            O => \N__11772\,
            I => \N__11757\
        );

    \I__2660\ : Span4Mux_h
    port map (
            O => \N__11769\,
            I => \N__11754\
        );

    \I__2659\ : InMux
    port map (
            O => \N__11768\,
            I => \N__11745\
        );

    \I__2658\ : InMux
    port map (
            O => \N__11767\,
            I => \N__11745\
        );

    \I__2657\ : InMux
    port map (
            O => \N__11766\,
            I => \N__11745\
        );

    \I__2656\ : InMux
    port map (
            O => \N__11765\,
            I => \N__11745\
        );

    \I__2655\ : InMux
    port map (
            O => \N__11764\,
            I => \N__11740\
        );

    \I__2654\ : InMux
    port map (
            O => \N__11763\,
            I => \N__11740\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__11760\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__11757\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__2651\ : Odrv4
    port map (
            O => \N__11754\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__11745\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__11740\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__2648\ : CascadeMux
    port map (
            O => \N__11729\,
            I => \N__11725\
        );

    \I__2647\ : CascadeMux
    port map (
            O => \N__11728\,
            I => \N__11720\
        );

    \I__2646\ : InMux
    port map (
            O => \N__11725\,
            I => \N__11714\
        );

    \I__2645\ : InMux
    port map (
            O => \N__11724\,
            I => \N__11705\
        );

    \I__2644\ : InMux
    port map (
            O => \N__11723\,
            I => \N__11705\
        );

    \I__2643\ : InMux
    port map (
            O => \N__11720\,
            I => \N__11705\
        );

    \I__2642\ : InMux
    port map (
            O => \N__11719\,
            I => \N__11705\
        );

    \I__2641\ : InMux
    port map (
            O => \N__11718\,
            I => \N__11700\
        );

    \I__2640\ : InMux
    port map (
            O => \N__11717\,
            I => \N__11700\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__11714\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_2\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__11705\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_2\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__11700\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_2\
        );

    \I__2636\ : InMux
    port map (
            O => \N__11693\,
            I => \N__11690\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__11690\,
            I => \DUT.uart_inst0.N_6_i\
        );

    \I__2634\ : InMux
    port map (
            O => \N__11687\,
            I => \N__11681\
        );

    \I__2633\ : InMux
    port map (
            O => \N__11686\,
            I => \N__11677\
        );

    \I__2632\ : InMux
    port map (
            O => \N__11685\,
            I => \N__11672\
        );

    \I__2631\ : InMux
    port map (
            O => \N__11684\,
            I => \N__11672\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__11681\,
            I => \N__11669\
        );

    \I__2629\ : InMux
    port map (
            O => \N__11680\,
            I => \N__11666\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__11677\,
            I => \N__11657\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__11672\,
            I => \N__11652\
        );

    \I__2626\ : Span4Mux_v
    port map (
            O => \N__11669\,
            I => \N__11652\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__11666\,
            I => \N__11649\
        );

    \I__2624\ : InMux
    port map (
            O => \N__11665\,
            I => \N__11638\
        );

    \I__2623\ : InMux
    port map (
            O => \N__11664\,
            I => \N__11638\
        );

    \I__2622\ : InMux
    port map (
            O => \N__11663\,
            I => \N__11638\
        );

    \I__2621\ : InMux
    port map (
            O => \N__11662\,
            I => \N__11638\
        );

    \I__2620\ : InMux
    port map (
            O => \N__11661\,
            I => \N__11638\
        );

    \I__2619\ : InMux
    port map (
            O => \N__11660\,
            I => \N__11633\
        );

    \I__2618\ : Span4Mux_h
    port map (
            O => \N__11657\,
            I => \N__11628\
        );

    \I__2617\ : Span4Mux_v
    port map (
            O => \N__11652\,
            I => \N__11628\
        );

    \I__2616\ : Span4Mux_v
    port map (
            O => \N__11649\,
            I => \N__11623\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__11638\,
            I => \N__11623\
        );

    \I__2614\ : InMux
    port map (
            O => \N__11637\,
            I => \N__11618\
        );

    \I__2613\ : InMux
    port map (
            O => \N__11636\,
            I => \N__11618\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__11633\,
            I => \DUT.rTransmitZ0\
        );

    \I__2611\ : Odrv4
    port map (
            O => \N__11628\,
            I => \DUT.rTransmitZ0\
        );

    \I__2610\ : Odrv4
    port map (
            O => \N__11623\,
            I => \DUT.rTransmitZ0\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__11618\,
            I => \DUT.rTransmitZ0\
        );

    \I__2608\ : InMux
    port map (
            O => \N__11609\,
            I => \N__11590\
        );

    \I__2607\ : InMux
    port map (
            O => \N__11608\,
            I => \N__11585\
        );

    \I__2606\ : InMux
    port map (
            O => \N__11607\,
            I => \N__11585\
        );

    \I__2605\ : InMux
    port map (
            O => \N__11606\,
            I => \N__11582\
        );

    \I__2604\ : InMux
    port map (
            O => \N__11605\,
            I => \N__11577\
        );

    \I__2603\ : InMux
    port map (
            O => \N__11604\,
            I => \N__11577\
        );

    \I__2602\ : CascadeMux
    port map (
            O => \N__11603\,
            I => \N__11573\
        );

    \I__2601\ : CascadeMux
    port map (
            O => \N__11602\,
            I => \N__11570\
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__11601\,
            I => \N__11567\
        );

    \I__2599\ : CascadeMux
    port map (
            O => \N__11600\,
            I => \N__11561\
        );

    \I__2598\ : CascadeMux
    port map (
            O => \N__11599\,
            I => \N__11558\
        );

    \I__2597\ : CascadeMux
    port map (
            O => \N__11598\,
            I => \N__11555\
        );

    \I__2596\ : CascadeMux
    port map (
            O => \N__11597\,
            I => \N__11552\
        );

    \I__2595\ : CascadeMux
    port map (
            O => \N__11596\,
            I => \N__11549\
        );

    \I__2594\ : CascadeMux
    port map (
            O => \N__11595\,
            I => \N__11542\
        );

    \I__2593\ : CascadeMux
    port map (
            O => \N__11594\,
            I => \N__11538\
        );

    \I__2592\ : CascadeMux
    port map (
            O => \N__11593\,
            I => \N__11533\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__11590\,
            I => \N__11530\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__11585\,
            I => \N__11527\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__11582\,
            I => \N__11524\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__11577\,
            I => \N__11521\
        );

    \I__2587\ : InMux
    port map (
            O => \N__11576\,
            I => \N__11508\
        );

    \I__2586\ : InMux
    port map (
            O => \N__11573\,
            I => \N__11508\
        );

    \I__2585\ : InMux
    port map (
            O => \N__11570\,
            I => \N__11508\
        );

    \I__2584\ : InMux
    port map (
            O => \N__11567\,
            I => \N__11508\
        );

    \I__2583\ : InMux
    port map (
            O => \N__11566\,
            I => \N__11508\
        );

    \I__2582\ : InMux
    port map (
            O => \N__11565\,
            I => \N__11508\
        );

    \I__2581\ : InMux
    port map (
            O => \N__11564\,
            I => \N__11505\
        );

    \I__2580\ : InMux
    port map (
            O => \N__11561\,
            I => \N__11500\
        );

    \I__2579\ : InMux
    port map (
            O => \N__11558\,
            I => \N__11500\
        );

    \I__2578\ : InMux
    port map (
            O => \N__11555\,
            I => \N__11483\
        );

    \I__2577\ : InMux
    port map (
            O => \N__11552\,
            I => \N__11483\
        );

    \I__2576\ : InMux
    port map (
            O => \N__11549\,
            I => \N__11483\
        );

    \I__2575\ : InMux
    port map (
            O => \N__11548\,
            I => \N__11483\
        );

    \I__2574\ : InMux
    port map (
            O => \N__11547\,
            I => \N__11483\
        );

    \I__2573\ : InMux
    port map (
            O => \N__11546\,
            I => \N__11483\
        );

    \I__2572\ : InMux
    port map (
            O => \N__11545\,
            I => \N__11483\
        );

    \I__2571\ : InMux
    port map (
            O => \N__11542\,
            I => \N__11483\
        );

    \I__2570\ : InMux
    port map (
            O => \N__11541\,
            I => \N__11480\
        );

    \I__2569\ : InMux
    port map (
            O => \N__11538\,
            I => \N__11477\
        );

    \I__2568\ : InMux
    port map (
            O => \N__11537\,
            I => \N__11472\
        );

    \I__2567\ : InMux
    port map (
            O => \N__11536\,
            I => \N__11472\
        );

    \I__2566\ : InMux
    port map (
            O => \N__11533\,
            I => \N__11469\
        );

    \I__2565\ : Span4Mux_v
    port map (
            O => \N__11530\,
            I => \N__11462\
        );

    \I__2564\ : Span4Mux_v
    port map (
            O => \N__11527\,
            I => \N__11462\
        );

    \I__2563\ : Span4Mux_v
    port map (
            O => \N__11524\,
            I => \N__11462\
        );

    \I__2562\ : Span4Mux_v
    port map (
            O => \N__11521\,
            I => \N__11457\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__11508\,
            I => \N__11457\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__11505\,
            I => \DUT.tx_state_0\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__11500\,
            I => \DUT.tx_state_0\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__11483\,
            I => \DUT.tx_state_0\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__11480\,
            I => \DUT.tx_state_0\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__11477\,
            I => \DUT.tx_state_0\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__11472\,
            I => \DUT.tx_state_0\
        );

    \I__2554\ : LocalMux
    port map (
            O => \N__11469\,
            I => \DUT.tx_state_0\
        );

    \I__2553\ : Odrv4
    port map (
            O => \N__11462\,
            I => \DUT.tx_state_0\
        );

    \I__2552\ : Odrv4
    port map (
            O => \N__11457\,
            I => \DUT.tx_state_0\
        );

    \I__2551\ : InMux
    port map (
            O => \N__11438\,
            I => \N__11434\
        );

    \I__2550\ : InMux
    port map (
            O => \N__11437\,
            I => \N__11428\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__11434\,
            I => \N__11425\
        );

    \I__2548\ : InMux
    port map (
            O => \N__11433\,
            I => \N__11420\
        );

    \I__2547\ : InMux
    port map (
            O => \N__11432\,
            I => \N__11420\
        );

    \I__2546\ : InMux
    port map (
            O => \N__11431\,
            I => \N__11417\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__11428\,
            I => \N__11403\
        );

    \I__2544\ : Span4Mux_h
    port map (
            O => \N__11425\,
            I => \N__11398\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__11420\,
            I => \N__11398\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__11417\,
            I => \N__11395\
        );

    \I__2541\ : InMux
    port map (
            O => \N__11416\,
            I => \N__11388\
        );

    \I__2540\ : InMux
    port map (
            O => \N__11415\,
            I => \N__11388\
        );

    \I__2539\ : InMux
    port map (
            O => \N__11414\,
            I => \N__11388\
        );

    \I__2538\ : InMux
    port map (
            O => \N__11413\,
            I => \N__11377\
        );

    \I__2537\ : InMux
    port map (
            O => \N__11412\,
            I => \N__11377\
        );

    \I__2536\ : InMux
    port map (
            O => \N__11411\,
            I => \N__11377\
        );

    \I__2535\ : InMux
    port map (
            O => \N__11410\,
            I => \N__11377\
        );

    \I__2534\ : InMux
    port map (
            O => \N__11409\,
            I => \N__11377\
        );

    \I__2533\ : InMux
    port map (
            O => \N__11408\,
            I => \N__11374\
        );

    \I__2532\ : InMux
    port map (
            O => \N__11407\,
            I => \N__11371\
        );

    \I__2531\ : InMux
    port map (
            O => \N__11406\,
            I => \N__11368\
        );

    \I__2530\ : Span4Mux_v
    port map (
            O => \N__11403\,
            I => \N__11361\
        );

    \I__2529\ : Span4Mux_v
    port map (
            O => \N__11398\,
            I => \N__11361\
        );

    \I__2528\ : Span4Mux_v
    port map (
            O => \N__11395\,
            I => \N__11361\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__11388\,
            I => \N__11358\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__11377\,
            I => \N__11355\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__11374\,
            I => \DUT.uart_inst0.tx_stateZ0Z_1\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__11371\,
            I => \DUT.uart_inst0.tx_stateZ0Z_1\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__11368\,
            I => \DUT.uart_inst0.tx_stateZ0Z_1\
        );

    \I__2522\ : Odrv4
    port map (
            O => \N__11361\,
            I => \DUT.uart_inst0.tx_stateZ0Z_1\
        );

    \I__2521\ : Odrv4
    port map (
            O => \N__11358\,
            I => \DUT.uart_inst0.tx_stateZ0Z_1\
        );

    \I__2520\ : Odrv4
    port map (
            O => \N__11355\,
            I => \DUT.uart_inst0.tx_stateZ0Z_1\
        );

    \I__2519\ : InMux
    port map (
            O => \N__11342\,
            I => \N__11339\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__11339\,
            I => \N__11336\
        );

    \I__2517\ : Odrv4
    port map (
            O => \N__11336\,
            I => \DUT.uart_inst0.N_11_1\
        );

    \I__2516\ : CascadeMux
    port map (
            O => \N__11333\,
            I => \N__11330\
        );

    \I__2515\ : InMux
    port map (
            O => \N__11330\,
            I => \N__11326\
        );

    \I__2514\ : InMux
    port map (
            O => \N__11329\,
            I => \N__11323\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__11326\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_9\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__11323\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_9\
        );

    \I__2511\ : InMux
    port map (
            O => \N__11318\,
            I => \N__11314\
        );

    \I__2510\ : InMux
    port map (
            O => \N__11317\,
            I => \N__11311\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__11314\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_10\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__11311\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_10\
        );

    \I__2507\ : CascadeMux
    port map (
            O => \N__11306\,
            I => \N__11302\
        );

    \I__2506\ : CascadeMux
    port map (
            O => \N__11305\,
            I => \N__11299\
        );

    \I__2505\ : InMux
    port map (
            O => \N__11302\,
            I => \N__11296\
        );

    \I__2504\ : InMux
    port map (
            O => \N__11299\,
            I => \N__11293\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__11296\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_11\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__11293\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_11\
        );

    \I__2501\ : InMux
    port map (
            O => \N__11288\,
            I => \N__11284\
        );

    \I__2500\ : InMux
    port map (
            O => \N__11287\,
            I => \N__11281\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__11284\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_8\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__11281\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_8\
        );

    \I__2497\ : SRMux
    port map (
            O => \N__11276\,
            I => \N__11273\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__11273\,
            I => \N__11269\
        );

    \I__2495\ : SRMux
    port map (
            O => \N__11272\,
            I => \N__11265\
        );

    \I__2494\ : Span4Mux_h
    port map (
            O => \N__11269\,
            I => \N__11262\
        );

    \I__2493\ : SRMux
    port map (
            O => \N__11268\,
            I => \N__11259\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__11265\,
            I => \DUT.uart_inst0.N_20\
        );

    \I__2491\ : Odrv4
    port map (
            O => \N__11262\,
            I => \DUT.uart_inst0.N_20\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__11259\,
            I => \DUT.uart_inst0.N_20\
        );

    \I__2489\ : InMux
    port map (
            O => \N__11252\,
            I => \N__11248\
        );

    \I__2488\ : InMux
    port map (
            O => \N__11251\,
            I => \N__11245\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__11248\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_1\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__11245\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_1\
        );

    \I__2485\ : InMux
    port map (
            O => \N__11240\,
            I => \N__11235\
        );

    \I__2484\ : InMux
    port map (
            O => \N__11239\,
            I => \N__11230\
        );

    \I__2483\ : InMux
    port map (
            O => \N__11238\,
            I => \N__11230\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__11235\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_0\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__11230\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_0\
        );

    \I__2480\ : CascadeMux
    port map (
            O => \N__11225\,
            I => \DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0_cascade_\
        );

    \I__2479\ : InMux
    port map (
            O => \N__11222\,
            I => \N__11218\
        );

    \I__2478\ : InMux
    port map (
            O => \N__11221\,
            I => \N__11215\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__11218\,
            I => \DUT.uart_inst0.N_77\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__11215\,
            I => \DUT.uart_inst0.N_77\
        );

    \I__2475\ : InMux
    port map (
            O => \N__11210\,
            I => \N__11207\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__11207\,
            I => \DUT.uart_inst0.g0_i_o2_2\
        );

    \I__2473\ : InMux
    port map (
            O => \N__11204\,
            I => \N__11201\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__11201\,
            I => \DUT.uart_inst0.g0_i_o2_3\
        );

    \I__2471\ : CascadeMux
    port map (
            O => \N__11198\,
            I => \N__11195\
        );

    \I__2470\ : InMux
    port map (
            O => \N__11195\,
            I => \N__11192\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__11192\,
            I => \N__11189\
        );

    \I__2468\ : Span4Mux_h
    port map (
            O => \N__11189\,
            I => \N__11186\
        );

    \I__2467\ : Odrv4
    port map (
            O => \N__11186\,
            I => \DUT.uart_inst0.N_11\
        );

    \I__2466\ : InMux
    port map (
            O => \N__11183\,
            I => \N__11180\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__11180\,
            I => \N__11177\
        );

    \I__2464\ : Span4Mux_h
    port map (
            O => \N__11177\,
            I => \N__11174\
        );

    \I__2463\ : Odrv4
    port map (
            O => \N__11174\,
            I => \DUT.uart_inst0.g0_11_a4_2\
        );

    \I__2462\ : CascadeMux
    port map (
            O => \N__11171\,
            I => \N__11168\
        );

    \I__2461\ : InMux
    port map (
            O => \N__11168\,
            I => \N__11165\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__11165\,
            I => \N__11162\
        );

    \I__2459\ : Span4Mux_v
    port map (
            O => \N__11162\,
            I => \N__11159\
        );

    \I__2458\ : Span4Mux_h
    port map (
            O => \N__11159\,
            I => \N__11156\
        );

    \I__2457\ : Odrv4
    port map (
            O => \N__11156\,
            I => \DUT.uart_inst0.N_9\
        );

    \I__2456\ : CascadeMux
    port map (
            O => \N__11153\,
            I => \DUT.uart_inst0.tx_state_ns_i_i_o2_a0_2_0_cascade_\
        );

    \I__2455\ : InMux
    port map (
            O => \N__11150\,
            I => \N__11146\
        );

    \I__2454\ : InMux
    port map (
            O => \N__11149\,
            I => \N__11143\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__11146\,
            I => \DUT.uart_inst0.N_71_i\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__11143\,
            I => \DUT.uart_inst0.N_71_i\
        );

    \I__2451\ : CascadeMux
    port map (
            O => \N__11138\,
            I => \N__11135\
        );

    \I__2450\ : InMux
    port map (
            O => \N__11135\,
            I => \N__11132\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__11132\,
            I => \N__11129\
        );

    \I__2448\ : Span4Mux_h
    port map (
            O => \N__11129\,
            I => \N__11126\
        );

    \I__2447\ : Odrv4
    port map (
            O => \N__11126\,
            I => \DUT.uart_inst0.N_8_1\
        );

    \I__2446\ : InMux
    port map (
            O => \N__11123\,
            I => \N__11117\
        );

    \I__2445\ : InMux
    port map (
            O => \N__11122\,
            I => \N__11112\
        );

    \I__2444\ : InMux
    port map (
            O => \N__11121\,
            I => \N__11112\
        );

    \I__2443\ : InMux
    port map (
            O => \N__11120\,
            I => \N__11109\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__11117\,
            I => \N__11105\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__11112\,
            I => \N__11100\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__11109\,
            I => \N__11100\
        );

    \I__2439\ : InMux
    port map (
            O => \N__11108\,
            I => \N__11097\
        );

    \I__2438\ : Span4Mux_v
    port map (
            O => \N__11105\,
            I => \N__11094\
        );

    \I__2437\ : Span4Mux_v
    port map (
            O => \N__11100\,
            I => \N__11089\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__11097\,
            I => \N__11089\
        );

    \I__2435\ : Sp12to4
    port map (
            O => \N__11094\,
            I => \N__11086\
        );

    \I__2434\ : Span4Mux_v
    port map (
            O => \N__11089\,
            I => \N__11083\
        );

    \I__2433\ : Span12Mux_h
    port map (
            O => \N__11086\,
            I => \N__11080\
        );

    \I__2432\ : Sp12to4
    port map (
            O => \N__11083\,
            I => \N__11077\
        );

    \I__2431\ : Span12Mux_v
    port map (
            O => \N__11080\,
            I => \N__11074\
        );

    \I__2430\ : Span12Mux_h
    port map (
            O => \N__11077\,
            I => \N__11071\
        );

    \I__2429\ : Odrv12
    port map (
            O => \N__11074\,
            I => \iRxF_n_c\
        );

    \I__2428\ : Odrv12
    port map (
            O => \N__11071\,
            I => \iRxF_n_c\
        );

    \I__2427\ : InMux
    port map (
            O => \N__11066\,
            I => \N__11062\
        );

    \I__2426\ : InMux
    port map (
            O => \N__11065\,
            I => \N__11058\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__11062\,
            I => \N__11055\
        );

    \I__2424\ : InMux
    port map (
            O => \N__11061\,
            I => \N__11052\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__11058\,
            I => \N__11049\
        );

    \I__2422\ : Span4Mux_v
    port map (
            O => \N__11055\,
            I => \N__11044\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__11052\,
            I => \N__11044\
        );

    \I__2420\ : Span4Mux_v
    port map (
            O => \N__11049\,
            I => \N__11041\
        );

    \I__2419\ : Span4Mux_v
    port map (
            O => \N__11044\,
            I => \N__11038\
        );

    \I__2418\ : Sp12to4
    port map (
            O => \N__11041\,
            I => \N__11035\
        );

    \I__2417\ : Sp12to4
    port map (
            O => \N__11038\,
            I => \N__11032\
        );

    \I__2416\ : Span12Mux_h
    port map (
            O => \N__11035\,
            I => \N__11029\
        );

    \I__2415\ : Span12Mux_h
    port map (
            O => \N__11032\,
            I => \N__11026\
        );

    \I__2414\ : Span12Mux_v
    port map (
            O => \N__11029\,
            I => \N__11023\
        );

    \I__2413\ : Span12Mux_v
    port map (
            O => \N__11026\,
            I => \N__11020\
        );

    \I__2412\ : Odrv12
    port map (
            O => \N__11023\,
            I => \iTxE_n_c\
        );

    \I__2411\ : Odrv12
    port map (
            O => \N__11020\,
            I => \iTxE_n_c\
        );

    \I__2410\ : InMux
    port map (
            O => \N__11015\,
            I => \N__11012\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__11012\,
            I => \N__11006\
        );

    \I__2408\ : InMux
    port map (
            O => \N__11011\,
            I => \N__11000\
        );

    \I__2407\ : InMux
    port map (
            O => \N__11010\,
            I => \N__11000\
        );

    \I__2406\ : InMux
    port map (
            O => \N__11009\,
            I => \N__10997\
        );

    \I__2405\ : Span4Mux_v
    port map (
            O => \N__11006\,
            I => \N__10994\
        );

    \I__2404\ : InMux
    port map (
            O => \N__11005\,
            I => \N__10991\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__11000\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_0\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__10997\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_0\
        );

    \I__2401\ : Odrv4
    port map (
            O => \N__10994\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_0\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__10991\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_0\
        );

    \I__2399\ : InMux
    port map (
            O => \N__10982\,
            I => \N__10979\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__10979\,
            I => \fifo_inst.ft2232h_inst.N_101\
        );

    \I__2397\ : CascadeMux
    port map (
            O => \N__10976\,
            I => \DUT.uart_inst0.N_13_cascade_\
        );

    \I__2396\ : CascadeMux
    port map (
            O => \N__10973\,
            I => \DUT.uart_inst0.g0_i_0_cascade_\
        );

    \I__2395\ : InMux
    port map (
            O => \N__10970\,
            I => \N__10967\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__10967\,
            I => \N__10964\
        );

    \I__2393\ : Odrv4
    port map (
            O => \N__10964\,
            I => \DUT.uart_inst0.g0_i_a6_0\
        );

    \I__2392\ : CascadeMux
    port map (
            O => \N__10961\,
            I => \DUT.uart_inst0.g0_i_1_cascade_\
        );

    \I__2391\ : InMux
    port map (
            O => \N__10958\,
            I => \N__10955\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__10955\,
            I => \DUT.uart_inst0.g0_i_a6_3_0\
        );

    \I__2389\ : CascadeMux
    port map (
            O => \N__10952\,
            I => \DUT.uart_inst0.g0_i_o2_1_cascade_\
        );

    \I__2388\ : InMux
    port map (
            O => \N__10949\,
            I => \N__10946\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__10946\,
            I => \N__10943\
        );

    \I__2386\ : Span4Mux_v
    port map (
            O => \N__10943\,
            I => \N__10940\
        );

    \I__2385\ : Odrv4
    port map (
            O => \N__10940\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_5\
        );

    \I__2384\ : CascadeMux
    port map (
            O => \N__10937\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_\
        );

    \I__2383\ : InMux
    port map (
            O => \N__10934\,
            I => \N__10931\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__10931\,
            I => \N__10928\
        );

    \I__2381\ : Span4Mux_h
    port map (
            O => \N__10928\,
            I => \N__10925\
        );

    \I__2380\ : Odrv4
    port map (
            O => \N__10925\,
            I => \DUT.rFifoDatarx_5\
        );

    \I__2379\ : InMux
    port map (
            O => \N__10922\,
            I => \N__10919\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__10919\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_5\
        );

    \I__2377\ : CascadeMux
    port map (
            O => \N__10916\,
            I => \N__10911\
        );

    \I__2376\ : InMux
    port map (
            O => \N__10915\,
            I => \N__10896\
        );

    \I__2375\ : InMux
    port map (
            O => \N__10914\,
            I => \N__10896\
        );

    \I__2374\ : InMux
    port map (
            O => \N__10911\,
            I => \N__10893\
        );

    \I__2373\ : InMux
    port map (
            O => \N__10910\,
            I => \N__10886\
        );

    \I__2372\ : InMux
    port map (
            O => \N__10909\,
            I => \N__10886\
        );

    \I__2371\ : InMux
    port map (
            O => \N__10908\,
            I => \N__10886\
        );

    \I__2370\ : InMux
    port map (
            O => \N__10907\,
            I => \N__10879\
        );

    \I__2369\ : InMux
    port map (
            O => \N__10906\,
            I => \N__10879\
        );

    \I__2368\ : InMux
    port map (
            O => \N__10905\,
            I => \N__10879\
        );

    \I__2367\ : InMux
    port map (
            O => \N__10904\,
            I => \N__10872\
        );

    \I__2366\ : InMux
    port map (
            O => \N__10903\,
            I => \N__10872\
        );

    \I__2365\ : InMux
    port map (
            O => \N__10902\,
            I => \N__10872\
        );

    \I__2364\ : InMux
    port map (
            O => \N__10901\,
            I => \N__10869\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__10896\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__10893\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__10886\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__10879\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__10872\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__10869\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__2357\ : CascadeMux
    port map (
            O => \N__10856\,
            I => \N__10843\
        );

    \I__2356\ : CascadeMux
    port map (
            O => \N__10855\,
            I => \N__10836\
        );

    \I__2355\ : CascadeMux
    port map (
            O => \N__10854\,
            I => \N__10833\
        );

    \I__2354\ : CascadeMux
    port map (
            O => \N__10853\,
            I => \N__10827\
        );

    \I__2353\ : CascadeMux
    port map (
            O => \N__10852\,
            I => \N__10822\
        );

    \I__2352\ : InMux
    port map (
            O => \N__10851\,
            I => \N__10819\
        );

    \I__2351\ : InMux
    port map (
            O => \N__10850\,
            I => \N__10816\
        );

    \I__2350\ : InMux
    port map (
            O => \N__10849\,
            I => \N__10803\
        );

    \I__2349\ : InMux
    port map (
            O => \N__10848\,
            I => \N__10803\
        );

    \I__2348\ : InMux
    port map (
            O => \N__10847\,
            I => \N__10803\
        );

    \I__2347\ : InMux
    port map (
            O => \N__10846\,
            I => \N__10803\
        );

    \I__2346\ : InMux
    port map (
            O => \N__10843\,
            I => \N__10803\
        );

    \I__2345\ : InMux
    port map (
            O => \N__10842\,
            I => \N__10803\
        );

    \I__2344\ : InMux
    port map (
            O => \N__10841\,
            I => \N__10790\
        );

    \I__2343\ : InMux
    port map (
            O => \N__10840\,
            I => \N__10790\
        );

    \I__2342\ : InMux
    port map (
            O => \N__10839\,
            I => \N__10790\
        );

    \I__2341\ : InMux
    port map (
            O => \N__10836\,
            I => \N__10790\
        );

    \I__2340\ : InMux
    port map (
            O => \N__10833\,
            I => \N__10790\
        );

    \I__2339\ : InMux
    port map (
            O => \N__10832\,
            I => \N__10790\
        );

    \I__2338\ : InMux
    port map (
            O => \N__10831\,
            I => \N__10779\
        );

    \I__2337\ : InMux
    port map (
            O => \N__10830\,
            I => \N__10779\
        );

    \I__2336\ : InMux
    port map (
            O => \N__10827\,
            I => \N__10779\
        );

    \I__2335\ : InMux
    port map (
            O => \N__10826\,
            I => \N__10779\
        );

    \I__2334\ : InMux
    port map (
            O => \N__10825\,
            I => \N__10779\
        );

    \I__2333\ : InMux
    port map (
            O => \N__10822\,
            I => \N__10776\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__10819\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__10816\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__10803\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__10790\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__10779\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__10776\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__2326\ : CascadeMux
    port map (
            O => \N__10763\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_\
        );

    \I__2325\ : InMux
    port map (
            O => \N__10760\,
            I => \N__10757\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__10757\,
            I => \N__10754\
        );

    \I__2323\ : Span4Mux_h
    port map (
            O => \N__10754\,
            I => \N__10751\
        );

    \I__2322\ : Odrv4
    port map (
            O => \N__10751\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_6\
        );

    \I__2321\ : InMux
    port map (
            O => \N__10748\,
            I => \N__10745\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__10745\,
            I => \N__10742\
        );

    \I__2319\ : Span4Mux_v
    port map (
            O => \N__10742\,
            I => \N__10739\
        );

    \I__2318\ : Odrv4
    port map (
            O => \N__10739\,
            I => \DUT.rFifoDatarx_6\
        );

    \I__2317\ : CascadeMux
    port map (
            O => \N__10736\,
            I => \N__10731\
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__10735\,
            I => \N__10726\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__10734\,
            I => \N__10723\
        );

    \I__2314\ : InMux
    port map (
            O => \N__10731\,
            I => \N__10718\
        );

    \I__2313\ : InMux
    port map (
            O => \N__10730\,
            I => \N__10718\
        );

    \I__2312\ : InMux
    port map (
            O => \N__10729\,
            I => \N__10715\
        );

    \I__2311\ : InMux
    port map (
            O => \N__10726\,
            I => \N__10710\
        );

    \I__2310\ : InMux
    port map (
            O => \N__10723\,
            I => \N__10710\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__10718\,
            I => \DUT.rFifoCount_0\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__10715\,
            I => \DUT.rFifoCount_0\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__10710\,
            I => \DUT.rFifoCount_0\
        );

    \I__2306\ : CascadeMux
    port map (
            O => \N__10703\,
            I => \N__10700\
        );

    \I__2305\ : InMux
    port map (
            O => \N__10700\,
            I => \N__10697\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__10697\,
            I => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0\
        );

    \I__2303\ : CascadeMux
    port map (
            O => \N__10694\,
            I => \N__10691\
        );

    \I__2302\ : InMux
    port map (
            O => \N__10691\,
            I => \N__10688\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__10688\,
            I => \DUT.fifo_tx_inst.rFifoCount_RNIBPFMZ0Z_1\
        );

    \I__2300\ : InMux
    port map (
            O => \N__10685\,
            I => \N__10679\
        );

    \I__2299\ : InMux
    port map (
            O => \N__10684\,
            I => \N__10672\
        );

    \I__2298\ : InMux
    port map (
            O => \N__10683\,
            I => \N__10672\
        );

    \I__2297\ : InMux
    port map (
            O => \N__10682\,
            I => \N__10672\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__10679\,
            I => \DUT.rFifoCount_1\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__10672\,
            I => \DUT.rFifoCount_1\
        );

    \I__2294\ : InMux
    port map (
            O => \N__10667\,
            I => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0\
        );

    \I__2293\ : InMux
    port map (
            O => \N__10664\,
            I => \N__10660\
        );

    \I__2292\ : InMux
    port map (
            O => \N__10663\,
            I => \N__10649\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__10660\,
            I => \N__10644\
        );

    \I__2290\ : InMux
    port map (
            O => \N__10659\,
            I => \N__10633\
        );

    \I__2289\ : InMux
    port map (
            O => \N__10658\,
            I => \N__10633\
        );

    \I__2288\ : InMux
    port map (
            O => \N__10657\,
            I => \N__10633\
        );

    \I__2287\ : InMux
    port map (
            O => \N__10656\,
            I => \N__10633\
        );

    \I__2286\ : InMux
    port map (
            O => \N__10655\,
            I => \N__10633\
        );

    \I__2285\ : InMux
    port map (
            O => \N__10654\,
            I => \N__10630\
        );

    \I__2284\ : InMux
    port map (
            O => \N__10653\,
            I => \N__10627\
        );

    \I__2283\ : InMux
    port map (
            O => \N__10652\,
            I => \N__10624\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__10649\,
            I => \N__10621\
        );

    \I__2281\ : InMux
    port map (
            O => \N__10648\,
            I => \N__10616\
        );

    \I__2280\ : InMux
    port map (
            O => \N__10647\,
            I => \N__10616\
        );

    \I__2279\ : Span4Mux_h
    port map (
            O => \N__10644\,
            I => \N__10611\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__10633\,
            I => \N__10611\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__10630\,
            I => \rRxReadZ0\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__10627\,
            I => \rRxReadZ0\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__10624\,
            I => \rRxReadZ0\
        );

    \I__2274\ : Odrv4
    port map (
            O => \N__10621\,
            I => \rRxReadZ0\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__10616\,
            I => \rRxReadZ0\
        );

    \I__2272\ : Odrv4
    port map (
            O => \N__10611\,
            I => \rRxReadZ0\
        );

    \I__2271\ : InMux
    port map (
            O => \N__10598\,
            I => \N__10589\
        );

    \I__2270\ : InMux
    port map (
            O => \N__10597\,
            I => \N__10589\
        );

    \I__2269\ : InMux
    port map (
            O => \N__10596\,
            I => \N__10586\
        );

    \I__2268\ : InMux
    port map (
            O => \N__10595\,
            I => \N__10581\
        );

    \I__2267\ : InMux
    port map (
            O => \N__10594\,
            I => \N__10581\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__10589\,
            I => \DUT.fifo_tx_inst.N_83\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__10586\,
            I => \DUT.fifo_tx_inst.N_83\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__10581\,
            I => \DUT.fifo_tx_inst.N_83\
        );

    \I__2263\ : InMux
    port map (
            O => \N__10574\,
            I => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1\
        );

    \I__2262\ : InMux
    port map (
            O => \N__10571\,
            I => \N__10568\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__10568\,
            I => \N__10564\
        );

    \I__2260\ : CascadeMux
    port map (
            O => \N__10567\,
            I => \N__10561\
        );

    \I__2259\ : Span4Mux_h
    port map (
            O => \N__10564\,
            I => \N__10558\
        );

    \I__2258\ : InMux
    port map (
            O => \N__10561\,
            I => \N__10550\
        );

    \I__2257\ : Span4Mux_v
    port map (
            O => \N__10558\,
            I => \N__10547\
        );

    \I__2256\ : InMux
    port map (
            O => \N__10557\,
            I => \N__10536\
        );

    \I__2255\ : InMux
    port map (
            O => \N__10556\,
            I => \N__10536\
        );

    \I__2254\ : InMux
    port map (
            O => \N__10555\,
            I => \N__10536\
        );

    \I__2253\ : InMux
    port map (
            O => \N__10554\,
            I => \N__10536\
        );

    \I__2252\ : InMux
    port map (
            O => \N__10553\,
            I => \N__10536\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__10550\,
            I => \DUT.rFifoCount_2\
        );

    \I__2250\ : Odrv4
    port map (
            O => \N__10547\,
            I => \DUT.rFifoCount_2\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__10536\,
            I => \DUT.rFifoCount_2\
        );

    \I__2248\ : SRMux
    port map (
            O => \N__10529\,
            I => \N__10502\
        );

    \I__2247\ : SRMux
    port map (
            O => \N__10528\,
            I => \N__10502\
        );

    \I__2246\ : SRMux
    port map (
            O => \N__10527\,
            I => \N__10502\
        );

    \I__2245\ : SRMux
    port map (
            O => \N__10526\,
            I => \N__10502\
        );

    \I__2244\ : SRMux
    port map (
            O => \N__10525\,
            I => \N__10502\
        );

    \I__2243\ : SRMux
    port map (
            O => \N__10524\,
            I => \N__10502\
        );

    \I__2242\ : SRMux
    port map (
            O => \N__10523\,
            I => \N__10502\
        );

    \I__2241\ : SRMux
    port map (
            O => \N__10522\,
            I => \N__10502\
        );

    \I__2240\ : SRMux
    port map (
            O => \N__10521\,
            I => \N__10502\
        );

    \I__2239\ : GlobalMux
    port map (
            O => \N__10502\,
            I => \N__10499\
        );

    \I__2238\ : gio2CtrlBuf
    port map (
            O => \N__10499\,
            I => \wPllLocked_i_g\
        );

    \I__2237\ : InMux
    port map (
            O => \N__10496\,
            I => \N__10493\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__10493\,
            I => \N__10487\
        );

    \I__2235\ : InMux
    port map (
            O => \N__10492\,
            I => \N__10484\
        );

    \I__2234\ : InMux
    port map (
            O => \N__10491\,
            I => \N__10481\
        );

    \I__2233\ : InMux
    port map (
            O => \N__10490\,
            I => \N__10478\
        );

    \I__2232\ : Span4Mux_h
    port map (
            O => \N__10487\,
            I => \N__10473\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__10484\,
            I => \N__10473\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__10481\,
            I => \N__10470\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__10478\,
            I => \N__10466\
        );

    \I__2228\ : Span4Mux_v
    port map (
            O => \N__10473\,
            I => \N__10461\
        );

    \I__2227\ : Span4Mux_h
    port map (
            O => \N__10470\,
            I => \N__10461\
        );

    \I__2226\ : InMux
    port map (
            O => \N__10469\,
            I => \N__10458\
        );

    \I__2225\ : Odrv12
    port map (
            O => \N__10466\,
            I => \DUT.wRxByte_7\
        );

    \I__2224\ : Odrv4
    port map (
            O => \N__10461\,
            I => \DUT.wRxByte_7\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__10458\,
            I => \DUT.wRxByte_7\
        );

    \I__2222\ : InMux
    port map (
            O => \N__10451\,
            I => \N__10448\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__10448\,
            I => \N__10445\
        );

    \I__2220\ : Odrv4
    port map (
            O => \N__10445\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_7\
        );

    \I__2219\ : CEMux
    port map (
            O => \N__10442\,
            I => \N__10438\
        );

    \I__2218\ : CEMux
    port map (
            O => \N__10441\,
            I => \N__10434\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__10438\,
            I => \N__10431\
        );

    \I__2216\ : CEMux
    port map (
            O => \N__10437\,
            I => \N__10428\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__10434\,
            I => \N__10425\
        );

    \I__2214\ : Span4Mux_v
    port map (
            O => \N__10431\,
            I => \N__10421\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__10428\,
            I => \N__10418\
        );

    \I__2212\ : Span4Mux_h
    port map (
            O => \N__10425\,
            I => \N__10415\
        );

    \I__2211\ : InMux
    port map (
            O => \N__10424\,
            I => \N__10412\
        );

    \I__2210\ : Odrv4
    port map (
            O => \N__10421\,
            I => \DUT.fifo_rx_inst.rFifoData_awe0\
        );

    \I__2209\ : Odrv4
    port map (
            O => \N__10418\,
            I => \DUT.fifo_rx_inst.rFifoData_awe0\
        );

    \I__2208\ : Odrv4
    port map (
            O => \N__10415\,
            I => \DUT.fifo_rx_inst.rFifoData_awe0\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__10412\,
            I => \DUT.fifo_rx_inst.rFifoData_awe0\
        );

    \I__2206\ : CascadeMux
    port map (
            O => \N__10403\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_\
        );

    \I__2205\ : InMux
    port map (
            O => \N__10400\,
            I => \N__10397\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__10397\,
            I => \N__10394\
        );

    \I__2203\ : Span4Mux_h
    port map (
            O => \N__10394\,
            I => \N__10391\
        );

    \I__2202\ : Odrv4
    port map (
            O => \N__10391\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_0\
        );

    \I__2201\ : InMux
    port map (
            O => \N__10388\,
            I => \N__10385\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__10385\,
            I => \N__10382\
        );

    \I__2199\ : Span4Mux_v
    port map (
            O => \N__10382\,
            I => \N__10379\
        );

    \I__2198\ : Odrv4
    port map (
            O => \N__10379\,
            I => \DUT.rFifoDatarxZ0Z_0\
        );

    \I__2197\ : InMux
    port map (
            O => \N__10376\,
            I => \N__10373\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__10373\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_0\
        );

    \I__2195\ : InMux
    port map (
            O => \N__10370\,
            I => \N__10367\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__10367\,
            I => \N__10364\
        );

    \I__2193\ : Span4Mux_h
    port map (
            O => \N__10364\,
            I => \N__10361\
        );

    \I__2192\ : Odrv4
    port map (
            O => \N__10361\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_1\
        );

    \I__2191\ : CascadeMux
    port map (
            O => \N__10358\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1_cascade_\
        );

    \I__2190\ : InMux
    port map (
            O => \N__10355\,
            I => \N__10352\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__10352\,
            I => \N__10349\
        );

    \I__2188\ : Span4Mux_v
    port map (
            O => \N__10349\,
            I => \N__10346\
        );

    \I__2187\ : Odrv4
    port map (
            O => \N__10346\,
            I => \DUT.rFifoDatarx_1\
        );

    \I__2186\ : CascadeMux
    port map (
            O => \N__10343\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_\
        );

    \I__2185\ : InMux
    port map (
            O => \N__10340\,
            I => \N__10337\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__10337\,
            I => \N__10334\
        );

    \I__2183\ : Span4Mux_v
    port map (
            O => \N__10334\,
            I => \N__10331\
        );

    \I__2182\ : Odrv4
    port map (
            O => \N__10331\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_4\
        );

    \I__2181\ : InMux
    port map (
            O => \N__10328\,
            I => \N__10325\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__10325\,
            I => \N__10322\
        );

    \I__2179\ : Span4Mux_h
    port map (
            O => \N__10322\,
            I => \N__10319\
        );

    \I__2178\ : Odrv4
    port map (
            O => \N__10319\,
            I => \DUT.rFifoDatarx_4\
        );

    \I__2177\ : InMux
    port map (
            O => \N__10316\,
            I => \N__10313\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__10313\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_4\
        );

    \I__2175\ : InMux
    port map (
            O => \N__10310\,
            I => \bfn_11_19_0_\
        );

    \I__2174\ : InMux
    port map (
            O => \N__10307\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_8\
        );

    \I__2173\ : InMux
    port map (
            O => \N__10304\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_9\
        );

    \I__2172\ : InMux
    port map (
            O => \N__10301\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_10\
        );

    \I__2171\ : InMux
    port map (
            O => \N__10298\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_11\
        );

    \I__2170\ : InMux
    port map (
            O => \N__10295\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_12\
        );

    \I__2169\ : InMux
    port map (
            O => \N__10292\,
            I => \N__10289\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__10289\,
            I => \N__10286\
        );

    \I__2167\ : Odrv12
    port map (
            O => \N__10286\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_7\
        );

    \I__2166\ : CascadeMux
    port map (
            O => \N__10283\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_\
        );

    \I__2165\ : InMux
    port map (
            O => \N__10280\,
            I => \N__10277\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__10277\,
            I => \N__10274\
        );

    \I__2163\ : Odrv4
    port map (
            O => \N__10274\,
            I => \DUT.rFifoDatarx_7\
        );

    \I__2162\ : InMux
    port map (
            O => \N__10271\,
            I => \N__10268\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__10268\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_7\
        );

    \I__2160\ : SRMux
    port map (
            O => \N__10265\,
            I => \N__10262\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__10262\,
            I => \N__10259\
        );

    \I__2158\ : Span4Mux_h
    port map (
            O => \N__10259\,
            I => \N__10256\
        );

    \I__2157\ : Span4Mux_h
    port map (
            O => \N__10256\,
            I => \N__10253\
        );

    \I__2156\ : Odrv4
    port map (
            O => \N__10253\,
            I => \DUT.uart_inst0.N_65_i\
        );

    \I__2155\ : CascadeMux
    port map (
            O => \N__10250\,
            I => \N__10247\
        );

    \I__2154\ : InMux
    port map (
            O => \N__10247\,
            I => \N__10243\
        );

    \I__2153\ : InMux
    port map (
            O => \N__10246\,
            I => \N__10240\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__10243\,
            I => \DUT.uart_inst0.tx_dataZ0Z_0\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__10240\,
            I => \DUT.uart_inst0.tx_dataZ0Z_0\
        );

    \I__2150\ : InMux
    port map (
            O => \N__10235\,
            I => \N__10229\
        );

    \I__2149\ : InMux
    port map (
            O => \N__10234\,
            I => \N__10226\
        );

    \I__2148\ : InMux
    port map (
            O => \N__10233\,
            I => \N__10223\
        );

    \I__2147\ : InMux
    port map (
            O => \N__10232\,
            I => \N__10220\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__10229\,
            I => \DUT.uart_inst0.N_85\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__10226\,
            I => \DUT.uart_inst0.N_85\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__10223\,
            I => \DUT.uart_inst0.N_85\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__10220\,
            I => \DUT.uart_inst0.N_85\
        );

    \I__2142\ : InMux
    port map (
            O => \N__10211\,
            I => \N__10208\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__10208\,
            I => \DUT.uart_inst0.N_89\
        );

    \I__2140\ : InMux
    port map (
            O => \N__10205\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_0\
        );

    \I__2139\ : InMux
    port map (
            O => \N__10202\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_1\
        );

    \I__2138\ : InMux
    port map (
            O => \N__10199\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_2\
        );

    \I__2137\ : InMux
    port map (
            O => \N__10196\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_3\
        );

    \I__2136\ : InMux
    port map (
            O => \N__10193\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_4\
        );

    \I__2135\ : InMux
    port map (
            O => \N__10190\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_5\
        );

    \I__2134\ : InMux
    port map (
            O => \N__10187\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_6\
        );

    \I__2133\ : CascadeMux
    port map (
            O => \N__10184\,
            I => \N__10181\
        );

    \I__2132\ : InMux
    port map (
            O => \N__10181\,
            I => \N__10175\
        );

    \I__2131\ : InMux
    port map (
            O => \N__10180\,
            I => \N__10175\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__10175\,
            I => \DUT.uart_inst0.N_100\
        );

    \I__2129\ : CascadeMux
    port map (
            O => \N__10172\,
            I => \N__10166\
        );

    \I__2128\ : CascadeMux
    port map (
            O => \N__10171\,
            I => \N__10162\
        );

    \I__2127\ : InMux
    port map (
            O => \N__10170\,
            I => \N__10158\
        );

    \I__2126\ : InMux
    port map (
            O => \N__10169\,
            I => \N__10155\
        );

    \I__2125\ : InMux
    port map (
            O => \N__10166\,
            I => \N__10150\
        );

    \I__2124\ : InMux
    port map (
            O => \N__10165\,
            I => \N__10150\
        );

    \I__2123\ : InMux
    port map (
            O => \N__10162\,
            I => \N__10147\
        );

    \I__2122\ : CascadeMux
    port map (
            O => \N__10161\,
            I => \N__10142\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__10158\,
            I => \N__10137\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__10155\,
            I => \N__10134\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__10150\,
            I => \N__10129\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__10147\,
            I => \N__10129\
        );

    \I__2117\ : InMux
    port map (
            O => \N__10146\,
            I => \N__10126\
        );

    \I__2116\ : InMux
    port map (
            O => \N__10145\,
            I => \N__10123\
        );

    \I__2115\ : InMux
    port map (
            O => \N__10142\,
            I => \N__10120\
        );

    \I__2114\ : InMux
    port map (
            O => \N__10141\,
            I => \N__10117\
        );

    \I__2113\ : CascadeMux
    port map (
            O => \N__10140\,
            I => \N__10112\
        );

    \I__2112\ : Span4Mux_v
    port map (
            O => \N__10137\,
            I => \N__10108\
        );

    \I__2111\ : Span4Mux_v
    port map (
            O => \N__10134\,
            I => \N__10105\
        );

    \I__2110\ : Span4Mux_v
    port map (
            O => \N__10129\,
            I => \N__10102\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__10126\,
            I => \N__10095\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__10123\,
            I => \N__10095\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__10120\,
            I => \N__10095\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__10117\,
            I => \N__10092\
        );

    \I__2105\ : InMux
    port map (
            O => \N__10116\,
            I => \N__10085\
        );

    \I__2104\ : InMux
    port map (
            O => \N__10115\,
            I => \N__10085\
        );

    \I__2103\ : InMux
    port map (
            O => \N__10112\,
            I => \N__10085\
        );

    \I__2102\ : InMux
    port map (
            O => \N__10111\,
            I => \N__10082\
        );

    \I__2101\ : Span4Mux_v
    port map (
            O => \N__10108\,
            I => \N__10075\
        );

    \I__2100\ : Span4Mux_v
    port map (
            O => \N__10105\,
            I => \N__10075\
        );

    \I__2099\ : Span4Mux_v
    port map (
            O => \N__10102\,
            I => \N__10075\
        );

    \I__2098\ : Span4Mux_v
    port map (
            O => \N__10095\,
            I => \N__10072\
        );

    \I__2097\ : Span4Mux_h
    port map (
            O => \N__10092\,
            I => \N__10067\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__10085\,
            I => \N__10067\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__10082\,
            I => \N__10064\
        );

    \I__2094\ : Sp12to4
    port map (
            O => \N__10075\,
            I => \N__10061\
        );

    \I__2093\ : Span4Mux_v
    port map (
            O => \N__10072\,
            I => \N__10056\
        );

    \I__2092\ : Span4Mux_v
    port map (
            O => \N__10067\,
            I => \N__10056\
        );

    \I__2091\ : Span12Mux_v
    port map (
            O => \N__10064\,
            I => \N__10049\
        );

    \I__2090\ : Span12Mux_h
    port map (
            O => \N__10061\,
            I => \N__10049\
        );

    \I__2089\ : Sp12to4
    port map (
            O => \N__10056\,
            I => \N__10049\
        );

    \I__2088\ : Odrv12
    port map (
            O => \N__10049\,
            I => \P1A1_c\
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__10046\,
            I => \N__10042\
        );

    \I__2086\ : CascadeMux
    port map (
            O => \N__10045\,
            I => \N__10036\
        );

    \I__2085\ : InMux
    port map (
            O => \N__10042\,
            I => \N__10032\
        );

    \I__2084\ : InMux
    port map (
            O => \N__10041\,
            I => \N__10029\
        );

    \I__2083\ : InMux
    port map (
            O => \N__10040\,
            I => \N__10026\
        );

    \I__2082\ : InMux
    port map (
            O => \N__10039\,
            I => \N__10023\
        );

    \I__2081\ : InMux
    port map (
            O => \N__10036\,
            I => \N__10020\
        );

    \I__2080\ : CascadeMux
    port map (
            O => \N__10035\,
            I => \N__10016\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__10032\,
            I => \N__10013\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__10029\,
            I => \N__10010\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__10026\,
            I => \N__10007\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__10023\,
            I => \N__10004\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__10020\,
            I => \N__10001\
        );

    \I__2074\ : InMux
    port map (
            O => \N__10019\,
            I => \N__9998\
        );

    \I__2073\ : InMux
    port map (
            O => \N__10016\,
            I => \N__9995\
        );

    \I__2072\ : Span4Mux_v
    port map (
            O => \N__10013\,
            I => \N__9988\
        );

    \I__2071\ : Span4Mux_h
    port map (
            O => \N__10010\,
            I => \N__9988\
        );

    \I__2070\ : Span4Mux_v
    port map (
            O => \N__10007\,
            I => \N__9988\
        );

    \I__2069\ : Odrv12
    port map (
            O => \N__10004\,
            I => \DUT.uart_inst0.recv_stateZ0Z_5\
        );

    \I__2068\ : Odrv12
    port map (
            O => \N__10001\,
            I => \DUT.uart_inst0.recv_stateZ0Z_5\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__9998\,
            I => \DUT.uart_inst0.recv_stateZ0Z_5\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__9995\,
            I => \DUT.uart_inst0.recv_stateZ0Z_5\
        );

    \I__2065\ : Odrv4
    port map (
            O => \N__9988\,
            I => \DUT.uart_inst0.recv_stateZ0Z_5\
        );

    \I__2064\ : InMux
    port map (
            O => \N__9977\,
            I => \N__9973\
        );

    \I__2063\ : InMux
    port map (
            O => \N__9976\,
            I => \N__9970\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__9973\,
            I => \N__9965\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__9970\,
            I => \N__9962\
        );

    \I__2060\ : InMux
    port map (
            O => \N__9969\,
            I => \N__9959\
        );

    \I__2059\ : InMux
    port map (
            O => \N__9968\,
            I => \N__9956\
        );

    \I__2058\ : Span4Mux_h
    port map (
            O => \N__9965\,
            I => \N__9953\
        );

    \I__2057\ : Span4Mux_h
    port map (
            O => \N__9962\,
            I => \N__9950\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__9959\,
            I => \N__9947\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__9956\,
            I => \DUT.uart_inst0.recv_stateZ0Z_0\
        );

    \I__2054\ : Odrv4
    port map (
            O => \N__9953\,
            I => \DUT.uart_inst0.recv_stateZ0Z_0\
        );

    \I__2053\ : Odrv4
    port map (
            O => \N__9950\,
            I => \DUT.uart_inst0.recv_stateZ0Z_0\
        );

    \I__2052\ : Odrv4
    port map (
            O => \N__9947\,
            I => \DUT.uart_inst0.recv_stateZ0Z_0\
        );

    \I__2051\ : InMux
    port map (
            O => \N__9938\,
            I => \N__9933\
        );

    \I__2050\ : InMux
    port map (
            O => \N__9937\,
            I => \N__9928\
        );

    \I__2049\ : InMux
    port map (
            O => \N__9936\,
            I => \N__9928\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__9933\,
            I => \N__9925\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__9928\,
            I => \N__9922\
        );

    \I__2046\ : Span12Mux_v
    port map (
            O => \N__9925\,
            I => \N__9919\
        );

    \I__2045\ : Span4Mux_h
    port map (
            O => \N__9922\,
            I => \N__9916\
        );

    \I__2044\ : Odrv12
    port map (
            O => \N__9919\,
            I => \DUT.uart_inst0.N_49\
        );

    \I__2043\ : Odrv4
    port map (
            O => \N__9916\,
            I => \DUT.uart_inst0.N_49\
        );

    \I__2042\ : InMux
    port map (
            O => \N__9911\,
            I => \N__9908\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__9908\,
            I => \N__9905\
        );

    \I__2040\ : Odrv12
    port map (
            O => \N__9905\,
            I => \fifo_inst.ft2232h_inst.rFifoStatec_0\
        );

    \I__2039\ : CascadeMux
    port map (
            O => \N__9902\,
            I => \N__9898\
        );

    \I__2038\ : CascadeMux
    port map (
            O => \N__9901\,
            I => \N__9893\
        );

    \I__2037\ : InMux
    port map (
            O => \N__9898\,
            I => \N__9890\
        );

    \I__2036\ : InMux
    port map (
            O => \N__9897\,
            I => \N__9883\
        );

    \I__2035\ : InMux
    port map (
            O => \N__9896\,
            I => \N__9883\
        );

    \I__2034\ : InMux
    port map (
            O => \N__9893\,
            I => \N__9883\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__9890\,
            I => \N__9880\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__9883\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_3\
        );

    \I__2031\ : Odrv4
    port map (
            O => \N__9880\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_3\
        );

    \I__2030\ : InMux
    port map (
            O => \N__9875\,
            I => \N__9865\
        );

    \I__2029\ : InMux
    port map (
            O => \N__9874\,
            I => \N__9865\
        );

    \I__2028\ : InMux
    port map (
            O => \N__9873\,
            I => \N__9865\
        );

    \I__2027\ : InMux
    port map (
            O => \N__9872\,
            I => \N__9862\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__9865\,
            I => \DUT.uart_inst0.N_139\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__9862\,
            I => \DUT.uart_inst0.N_139\
        );

    \I__2024\ : CascadeMux
    port map (
            O => \N__9857\,
            I => \N__9853\
        );

    \I__2023\ : InMux
    port map (
            O => \N__9856\,
            I => \N__9845\
        );

    \I__2022\ : InMux
    port map (
            O => \N__9853\,
            I => \N__9845\
        );

    \I__2021\ : InMux
    port map (
            O => \N__9852\,
            I => \N__9845\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__9845\,
            I => \N__9840\
        );

    \I__2019\ : InMux
    port map (
            O => \N__9844\,
            I => \N__9835\
        );

    \I__2018\ : InMux
    port map (
            O => \N__9843\,
            I => \N__9835\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__9840\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_2\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__9835\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_2\
        );

    \I__2015\ : InMux
    port map (
            O => \N__9830\,
            I => \N__9826\
        );

    \I__2014\ : InMux
    port map (
            O => \N__9829\,
            I => \N__9822\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__9826\,
            I => \N__9819\
        );

    \I__2012\ : InMux
    port map (
            O => \N__9825\,
            I => \N__9816\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__9822\,
            I => \DUT.rTransmitc_0\
        );

    \I__2010\ : Odrv4
    port map (
            O => \N__9819\,
            I => \DUT.rTransmitc_0\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__9816\,
            I => \DUT.rTransmitc_0\
        );

    \I__2008\ : CascadeMux
    port map (
            O => \N__9809\,
            I => \DUT.uart_inst0.N_85_cascade_\
        );

    \I__2007\ : InMux
    port map (
            O => \N__9806\,
            I => \N__9803\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__9803\,
            I => \N__9798\
        );

    \I__2005\ : InMux
    port map (
            O => \N__9802\,
            I => \N__9795\
        );

    \I__2004\ : InMux
    port map (
            O => \N__9801\,
            I => \N__9792\
        );

    \I__2003\ : Odrv4
    port map (
            O => \N__9798\,
            I => \DUT.uart_inst0.N_66\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__9795\,
            I => \DUT.uart_inst0.N_66\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__9792\,
            I => \DUT.uart_inst0.N_66\
        );

    \I__2000\ : CascadeMux
    port map (
            O => \N__9785\,
            I => \DUT.uart_inst0.N_22_cascade_\
        );

    \I__1999\ : InMux
    port map (
            O => \N__9782\,
            I => \N__9773\
        );

    \I__1998\ : InMux
    port map (
            O => \N__9781\,
            I => \N__9773\
        );

    \I__1997\ : InMux
    port map (
            O => \N__9780\,
            I => \N__9773\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__9773\,
            I => \N__9766\
        );

    \I__1995\ : InMux
    port map (
            O => \N__9772\,
            I => \N__9757\
        );

    \I__1994\ : InMux
    port map (
            O => \N__9771\,
            I => \N__9757\
        );

    \I__1993\ : InMux
    port map (
            O => \N__9770\,
            I => \N__9757\
        );

    \I__1992\ : InMux
    port map (
            O => \N__9769\,
            I => \N__9757\
        );

    \I__1991\ : Odrv4
    port map (
            O => \N__9766\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_0\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__9757\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_0\
        );

    \I__1989\ : InMux
    port map (
            O => \N__9752\,
            I => \N__9749\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__9749\,
            I => \N__9744\
        );

    \I__1987\ : InMux
    port map (
            O => \N__9748\,
            I => \N__9739\
        );

    \I__1986\ : InMux
    port map (
            O => \N__9747\,
            I => \N__9739\
        );

    \I__1985\ : Odrv4
    port map (
            O => \N__9744\,
            I => \DUT.uart_inst0.N_22\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__9739\,
            I => \DUT.uart_inst0.N_22\
        );

    \I__1983\ : InMux
    port map (
            O => \N__9734\,
            I => \N__9723\
        );

    \I__1982\ : InMux
    port map (
            O => \N__9733\,
            I => \N__9723\
        );

    \I__1981\ : InMux
    port map (
            O => \N__9732\,
            I => \N__9723\
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__9731\,
            I => \N__9720\
        );

    \I__1979\ : CascadeMux
    port map (
            O => \N__9730\,
            I => \N__9717\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__9723\,
            I => \N__9713\
        );

    \I__1977\ : InMux
    port map (
            O => \N__9720\,
            I => \N__9706\
        );

    \I__1976\ : InMux
    port map (
            O => \N__9717\,
            I => \N__9706\
        );

    \I__1975\ : InMux
    port map (
            O => \N__9716\,
            I => \N__9706\
        );

    \I__1974\ : Odrv4
    port map (
            O => \N__9713\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_1\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__9706\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_1\
        );

    \I__1972\ : InMux
    port map (
            O => \N__9701\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_16\
        );

    \I__1971\ : CascadeMux
    port map (
            O => \N__9698\,
            I => \N__9694\
        );

    \I__1970\ : InMux
    port map (
            O => \N__9697\,
            I => \N__9691\
        );

    \I__1969\ : InMux
    port map (
            O => \N__9694\,
            I => \N__9688\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__9691\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_17\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__9688\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_17\
        );

    \I__1966\ : InMux
    port map (
            O => \N__9683\,
            I => \N__9680\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__9680\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO\
        );

    \I__1964\ : InMux
    port map (
            O => \N__9677\,
            I => \N__9672\
        );

    \I__1963\ : InMux
    port map (
            O => \N__9676\,
            I => \N__9669\
        );

    \I__1962\ : InMux
    port map (
            O => \N__9675\,
            I => \N__9666\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__9672\,
            I => \N__9661\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__9669\,
            I => \N__9661\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__9666\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_12\
        );

    \I__1958\ : Odrv4
    port map (
            O => \N__9661\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_12\
        );

    \I__1957\ : InMux
    port map (
            O => \N__9656\,
            I => \N__9653\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__9653\,
            I => \N__9650\
        );

    \I__1955\ : Odrv12
    port map (
            O => \N__9650\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO\
        );

    \I__1954\ : InMux
    port map (
            O => \N__9647\,
            I => \N__9642\
        );

    \I__1953\ : InMux
    port map (
            O => \N__9646\,
            I => \N__9639\
        );

    \I__1952\ : InMux
    port map (
            O => \N__9645\,
            I => \N__9636\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__9642\,
            I => \N__9633\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__9639\,
            I => \N__9630\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__9636\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_2\
        );

    \I__1948\ : Odrv4
    port map (
            O => \N__9633\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_2\
        );

    \I__1947\ : Odrv4
    port map (
            O => \N__9630\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_2\
        );

    \I__1946\ : InMux
    port map (
            O => \N__9623\,
            I => \N__9620\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__9620\,
            I => \N__9617\
        );

    \I__1944\ : Odrv4
    port map (
            O => \N__9617\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO\
        );

    \I__1943\ : CascadeMux
    port map (
            O => \N__9614\,
            I => \N__9602\
        );

    \I__1942\ : CascadeMux
    port map (
            O => \N__9613\,
            I => \N__9596\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__9612\,
            I => \N__9592\
        );

    \I__1940\ : InMux
    port map (
            O => \N__9611\,
            I => \N__9581\
        );

    \I__1939\ : InMux
    port map (
            O => \N__9610\,
            I => \N__9581\
        );

    \I__1938\ : InMux
    port map (
            O => \N__9609\,
            I => \N__9581\
        );

    \I__1937\ : InMux
    port map (
            O => \N__9608\,
            I => \N__9581\
        );

    \I__1936\ : InMux
    port map (
            O => \N__9607\,
            I => \N__9567\
        );

    \I__1935\ : InMux
    port map (
            O => \N__9606\,
            I => \N__9567\
        );

    \I__1934\ : InMux
    port map (
            O => \N__9605\,
            I => \N__9567\
        );

    \I__1933\ : InMux
    port map (
            O => \N__9602\,
            I => \N__9567\
        );

    \I__1932\ : InMux
    port map (
            O => \N__9601\,
            I => \N__9567\
        );

    \I__1931\ : InMux
    port map (
            O => \N__9600\,
            I => \N__9567\
        );

    \I__1930\ : InMux
    port map (
            O => \N__9599\,
            I => \N__9551\
        );

    \I__1929\ : InMux
    port map (
            O => \N__9596\,
            I => \N__9551\
        );

    \I__1928\ : InMux
    port map (
            O => \N__9595\,
            I => \N__9551\
        );

    \I__1927\ : InMux
    port map (
            O => \N__9592\,
            I => \N__9551\
        );

    \I__1926\ : InMux
    port map (
            O => \N__9591\,
            I => \N__9551\
        );

    \I__1925\ : InMux
    port map (
            O => \N__9590\,
            I => \N__9551\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__9581\,
            I => \N__9548\
        );

    \I__1923\ : InMux
    port map (
            O => \N__9580\,
            I => \N__9545\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__9567\,
            I => \N__9542\
        );

    \I__1921\ : InMux
    port map (
            O => \N__9566\,
            I => \N__9536\
        );

    \I__1920\ : InMux
    port map (
            O => \N__9565\,
            I => \N__9533\
        );

    \I__1919\ : InMux
    port map (
            O => \N__9564\,
            I => \N__9530\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__9551\,
            I => \N__9527\
        );

    \I__1917\ : Span4Mux_h
    port map (
            O => \N__9548\,
            I => \N__9524\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__9545\,
            I => \N__9519\
        );

    \I__1915\ : Span4Mux_h
    port map (
            O => \N__9542\,
            I => \N__9519\
        );

    \I__1914\ : InMux
    port map (
            O => \N__9541\,
            I => \N__9516\
        );

    \I__1913\ : InMux
    port map (
            O => \N__9540\,
            I => \N__9511\
        );

    \I__1912\ : InMux
    port map (
            O => \N__9539\,
            I => \N__9511\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__9536\,
            I => \N__9506\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__9533\,
            I => \N__9506\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__9530\,
            I => \DUT.uart_inst0.N_50\
        );

    \I__1908\ : Odrv4
    port map (
            O => \N__9527\,
            I => \DUT.uart_inst0.N_50\
        );

    \I__1907\ : Odrv4
    port map (
            O => \N__9524\,
            I => \DUT.uart_inst0.N_50\
        );

    \I__1906\ : Odrv4
    port map (
            O => \N__9519\,
            I => \DUT.uart_inst0.N_50\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__9516\,
            I => \DUT.uart_inst0.N_50\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__9511\,
            I => \DUT.uart_inst0.N_50\
        );

    \I__1903\ : Odrv4
    port map (
            O => \N__9506\,
            I => \DUT.uart_inst0.N_50\
        );

    \I__1902\ : CascadeMux
    port map (
            O => \N__9491\,
            I => \N__9487\
        );

    \I__1901\ : InMux
    port map (
            O => \N__9490\,
            I => \N__9483\
        );

    \I__1900\ : InMux
    port map (
            O => \N__9487\,
            I => \N__9480\
        );

    \I__1899\ : InMux
    port map (
            O => \N__9486\,
            I => \N__9477\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__9483\,
            I => \N__9474\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__9480\,
            I => \N__9471\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__9477\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_4\
        );

    \I__1895\ : Odrv4
    port map (
            O => \N__9474\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_4\
        );

    \I__1894\ : Odrv4
    port map (
            O => \N__9471\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_4\
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__9464\,
            I => \DUT.uart_inst0.N_98_cascade_\
        );

    \I__1892\ : IoInMux
    port map (
            O => \N__9461\,
            I => \N__9458\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__9458\,
            I => \N__9455\
        );

    \I__1890\ : Span4Mux_s3_v
    port map (
            O => \N__9455\,
            I => \N__9452\
        );

    \I__1889\ : Span4Mux_v
    port map (
            O => \N__9452\,
            I => \N__9449\
        );

    \I__1888\ : Span4Mux_v
    port map (
            O => \N__9449\,
            I => \N__9445\
        );

    \I__1887\ : InMux
    port map (
            O => \N__9448\,
            I => \N__9442\
        );

    \I__1886\ : Span4Mux_v
    port map (
            O => \N__9445\,
            I => \N__9439\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__9442\,
            I => \N__9436\
        );

    \I__1884\ : Odrv4
    port map (
            O => \N__9439\,
            I => \P1A7_c\
        );

    \I__1883\ : Odrv4
    port map (
            O => \N__9436\,
            I => \P1A7_c\
        );

    \I__1882\ : InMux
    port map (
            O => \N__9431\,
            I => \N__9428\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__9428\,
            I => \DUT.uart_inst0.N_82\
        );

    \I__1880\ : InMux
    port map (
            O => \N__9425\,
            I => \N__9419\
        );

    \I__1879\ : InMux
    port map (
            O => \N__9424\,
            I => \N__9419\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__9419\,
            I => \DUT.uart_inst0.N_99\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__9416\,
            I => \N__9411\
        );

    \I__1876\ : InMux
    port map (
            O => \N__9415\,
            I => \N__9408\
        );

    \I__1875\ : InMux
    port map (
            O => \N__9414\,
            I => \N__9403\
        );

    \I__1874\ : InMux
    port map (
            O => \N__9411\,
            I => \N__9403\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__9408\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_9\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__9403\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_9\
        );

    \I__1871\ : CascadeMux
    port map (
            O => \N__9398\,
            I => \N__9395\
        );

    \I__1870\ : InMux
    port map (
            O => \N__9395\,
            I => \N__9392\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__9392\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO\
        );

    \I__1868\ : InMux
    port map (
            O => \N__9389\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_8\
        );

    \I__1867\ : InMux
    port map (
            O => \N__9386\,
            I => \N__9381\
        );

    \I__1866\ : InMux
    port map (
            O => \N__9385\,
            I => \N__9378\
        );

    \I__1865\ : InMux
    port map (
            O => \N__9384\,
            I => \N__9375\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__9381\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_10\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__9378\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_10\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__9375\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_10\
        );

    \I__1861\ : InMux
    port map (
            O => \N__9368\,
            I => \N__9365\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__9365\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO\
        );

    \I__1859\ : InMux
    port map (
            O => \N__9362\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_9\
        );

    \I__1858\ : InMux
    port map (
            O => \N__9359\,
            I => \N__9354\
        );

    \I__1857\ : InMux
    port map (
            O => \N__9358\,
            I => \N__9351\
        );

    \I__1856\ : InMux
    port map (
            O => \N__9357\,
            I => \N__9348\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__9354\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_11\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__9351\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_11\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__9348\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_11\
        );

    \I__1852\ : InMux
    port map (
            O => \N__9341\,
            I => \N__9338\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__9338\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO\
        );

    \I__1850\ : InMux
    port map (
            O => \N__9335\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_10\
        );

    \I__1849\ : InMux
    port map (
            O => \N__9332\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_11\
        );

    \I__1848\ : InMux
    port map (
            O => \N__9329\,
            I => \N__9324\
        );

    \I__1847\ : InMux
    port map (
            O => \N__9328\,
            I => \N__9319\
        );

    \I__1846\ : InMux
    port map (
            O => \N__9327\,
            I => \N__9319\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__9324\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_13\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__9319\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_13\
        );

    \I__1843\ : InMux
    port map (
            O => \N__9314\,
            I => \N__9311\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__9311\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO\
        );

    \I__1841\ : InMux
    port map (
            O => \N__9308\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_12\
        );

    \I__1840\ : InMux
    port map (
            O => \N__9305\,
            I => \N__9300\
        );

    \I__1839\ : InMux
    port map (
            O => \N__9304\,
            I => \N__9297\
        );

    \I__1838\ : InMux
    port map (
            O => \N__9303\,
            I => \N__9294\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__9300\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_14\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__9297\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_14\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__9294\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_14\
        );

    \I__1834\ : InMux
    port map (
            O => \N__9287\,
            I => \N__9284\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__9284\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO\
        );

    \I__1832\ : InMux
    port map (
            O => \N__9281\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_13\
        );

    \I__1831\ : InMux
    port map (
            O => \N__9278\,
            I => \N__9273\
        );

    \I__1830\ : InMux
    port map (
            O => \N__9277\,
            I => \N__9268\
        );

    \I__1829\ : InMux
    port map (
            O => \N__9276\,
            I => \N__9268\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__9273\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_15\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__9268\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_15\
        );

    \I__1826\ : InMux
    port map (
            O => \N__9263\,
            I => \N__9260\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__9260\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO\
        );

    \I__1824\ : InMux
    port map (
            O => \N__9257\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_14\
        );

    \I__1823\ : InMux
    port map (
            O => \N__9254\,
            I => \N__9249\
        );

    \I__1822\ : InMux
    port map (
            O => \N__9253\,
            I => \N__9246\
        );

    \I__1821\ : InMux
    port map (
            O => \N__9252\,
            I => \N__9243\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__9249\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_16\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__9246\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_16\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__9243\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_16\
        );

    \I__1817\ : InMux
    port map (
            O => \N__9236\,
            I => \N__9233\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__9233\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO\
        );

    \I__1815\ : InMux
    port map (
            O => \N__9230\,
            I => \bfn_11_15_0_\
        );

    \I__1814\ : InMux
    port map (
            O => \N__9227\,
            I => \N__9224\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__9224\,
            I => \N__9221\
        );

    \I__1812\ : Span4Mux_h
    port map (
            O => \N__9221\,
            I => \N__9216\
        );

    \I__1811\ : InMux
    port map (
            O => \N__9220\,
            I => \N__9211\
        );

    \I__1810\ : InMux
    port map (
            O => \N__9219\,
            I => \N__9211\
        );

    \I__1809\ : Odrv4
    port map (
            O => \N__9216\,
            I => \DUT.uart_inst0.rx_clk_dividerZ1Z_1\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__9211\,
            I => \DUT.uart_inst0.rx_clk_dividerZ1Z_1\
        );

    \I__1807\ : InMux
    port map (
            O => \N__9206\,
            I => \N__9203\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__9203\,
            I => \N__9200\
        );

    \I__1805\ : Span4Mux_h
    port map (
            O => \N__9200\,
            I => \N__9197\
        );

    \I__1804\ : Odrv4
    port map (
            O => \N__9197\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO\
        );

    \I__1803\ : InMux
    port map (
            O => \N__9194\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_0\
        );

    \I__1802\ : InMux
    port map (
            O => \N__9191\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_1\
        );

    \I__1801\ : InMux
    port map (
            O => \N__9188\,
            I => \N__9185\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__9185\,
            I => \N__9182\
        );

    \I__1799\ : Span4Mux_h
    port map (
            O => \N__9182\,
            I => \N__9177\
        );

    \I__1798\ : InMux
    port map (
            O => \N__9181\,
            I => \N__9172\
        );

    \I__1797\ : InMux
    port map (
            O => \N__9180\,
            I => \N__9172\
        );

    \I__1796\ : Odrv4
    port map (
            O => \N__9177\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_3\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__9172\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_3\
        );

    \I__1794\ : CascadeMux
    port map (
            O => \N__9167\,
            I => \N__9164\
        );

    \I__1793\ : InMux
    port map (
            O => \N__9164\,
            I => \N__9161\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__9161\,
            I => \N__9158\
        );

    \I__1791\ : Span4Mux_v
    port map (
            O => \N__9158\,
            I => \N__9155\
        );

    \I__1790\ : Span4Mux_h
    port map (
            O => \N__9155\,
            I => \N__9152\
        );

    \I__1789\ : Odrv4
    port map (
            O => \N__9152\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_2_THRU_CO\
        );

    \I__1788\ : InMux
    port map (
            O => \N__9149\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_2\
        );

    \I__1787\ : InMux
    port map (
            O => \N__9146\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_3\
        );

    \I__1786\ : InMux
    port map (
            O => \N__9143\,
            I => \N__9138\
        );

    \I__1785\ : InMux
    port map (
            O => \N__9142\,
            I => \N__9133\
        );

    \I__1784\ : InMux
    port map (
            O => \N__9141\,
            I => \N__9133\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__9138\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_5\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__9133\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_5\
        );

    \I__1781\ : InMux
    port map (
            O => \N__9128\,
            I => \N__9125\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__9125\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_4_THRU_CO\
        );

    \I__1779\ : InMux
    port map (
            O => \N__9122\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_4\
        );

    \I__1778\ : CascadeMux
    port map (
            O => \N__9119\,
            I => \N__9115\
        );

    \I__1777\ : InMux
    port map (
            O => \N__9118\,
            I => \N__9111\
        );

    \I__1776\ : InMux
    port map (
            O => \N__9115\,
            I => \N__9106\
        );

    \I__1775\ : InMux
    port map (
            O => \N__9114\,
            I => \N__9106\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__9111\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_6\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__9106\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_6\
        );

    \I__1772\ : InMux
    port map (
            O => \N__9101\,
            I => \N__9098\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__9098\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_5_THRU_CO\
        );

    \I__1770\ : InMux
    port map (
            O => \N__9095\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_5\
        );

    \I__1769\ : InMux
    port map (
            O => \N__9092\,
            I => \N__9087\
        );

    \I__1768\ : InMux
    port map (
            O => \N__9091\,
            I => \N__9084\
        );

    \I__1767\ : InMux
    port map (
            O => \N__9090\,
            I => \N__9081\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__9087\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_7\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__9084\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_7\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__9081\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_7\
        );

    \I__1763\ : InMux
    port map (
            O => \N__9074\,
            I => \N__9071\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__9071\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO\
        );

    \I__1761\ : InMux
    port map (
            O => \N__9068\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_6\
        );

    \I__1760\ : CascadeMux
    port map (
            O => \N__9065\,
            I => \N__9060\
        );

    \I__1759\ : InMux
    port map (
            O => \N__9064\,
            I => \N__9057\
        );

    \I__1758\ : InMux
    port map (
            O => \N__9063\,
            I => \N__9052\
        );

    \I__1757\ : InMux
    port map (
            O => \N__9060\,
            I => \N__9052\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__9057\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_8\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__9052\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_8\
        );

    \I__1754\ : InMux
    port map (
            O => \N__9047\,
            I => \N__9044\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__9044\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO\
        );

    \I__1752\ : InMux
    port map (
            O => \N__9041\,
            I => \bfn_11_14_0_\
        );

    \I__1751\ : CascadeMux
    port map (
            O => \N__9038\,
            I => \N__9035\
        );

    \I__1750\ : InMux
    port map (
            O => \N__9035\,
            I => \N__9029\
        );

    \I__1749\ : InMux
    port map (
            O => \N__9034\,
            I => \N__9029\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__9029\,
            I => \DUT.fifo_tx_inst.un1_i11_2_i\
        );

    \I__1747\ : CascadeMux
    port map (
            O => \N__9026\,
            I => \N__9021\
        );

    \I__1746\ : CascadeMux
    port map (
            O => \N__9025\,
            I => \N__9012\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__9024\,
            I => \N__9006\
        );

    \I__1744\ : InMux
    port map (
            O => \N__9021\,
            I => \N__9000\
        );

    \I__1743\ : InMux
    port map (
            O => \N__9020\,
            I => \N__8995\
        );

    \I__1742\ : InMux
    port map (
            O => \N__9019\,
            I => \N__8995\
        );

    \I__1741\ : InMux
    port map (
            O => \N__9018\,
            I => \N__8978\
        );

    \I__1740\ : InMux
    port map (
            O => \N__9017\,
            I => \N__8978\
        );

    \I__1739\ : InMux
    port map (
            O => \N__9016\,
            I => \N__8978\
        );

    \I__1738\ : InMux
    port map (
            O => \N__9015\,
            I => \N__8978\
        );

    \I__1737\ : InMux
    port map (
            O => \N__9012\,
            I => \N__8978\
        );

    \I__1736\ : InMux
    port map (
            O => \N__9011\,
            I => \N__8978\
        );

    \I__1735\ : InMux
    port map (
            O => \N__9010\,
            I => \N__8978\
        );

    \I__1734\ : InMux
    port map (
            O => \N__9009\,
            I => \N__8978\
        );

    \I__1733\ : InMux
    port map (
            O => \N__9006\,
            I => \N__8969\
        );

    \I__1732\ : InMux
    port map (
            O => \N__9005\,
            I => \N__8969\
        );

    \I__1731\ : InMux
    port map (
            O => \N__9004\,
            I => \N__8969\
        );

    \I__1730\ : CascadeMux
    port map (
            O => \N__9003\,
            I => \N__8965\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__9000\,
            I => \N__8961\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__8995\,
            I => \N__8956\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__8978\,
            I => \N__8956\
        );

    \I__1726\ : InMux
    port map (
            O => \N__8977\,
            I => \N__8953\
        );

    \I__1725\ : InMux
    port map (
            O => \N__8976\,
            I => \N__8950\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__8969\,
            I => \N__8947\
        );

    \I__1723\ : CascadeMux
    port map (
            O => \N__8968\,
            I => \N__8943\
        );

    \I__1722\ : InMux
    port map (
            O => \N__8965\,
            I => \N__8938\
        );

    \I__1721\ : InMux
    port map (
            O => \N__8964\,
            I => \N__8938\
        );

    \I__1720\ : Span4Mux_v
    port map (
            O => \N__8961\,
            I => \N__8935\
        );

    \I__1719\ : Span4Mux_v
    port map (
            O => \N__8956\,
            I => \N__8930\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__8953\,
            I => \N__8930\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__8950\,
            I => \N__8925\
        );

    \I__1716\ : Span4Mux_h
    port map (
            O => \N__8947\,
            I => \N__8925\
        );

    \I__1715\ : InMux
    port map (
            O => \N__8946\,
            I => \N__8920\
        );

    \I__1714\ : InMux
    port map (
            O => \N__8943\,
            I => \N__8920\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__8938\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__1712\ : Odrv4
    port map (
            O => \N__8935\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__1711\ : Odrv4
    port map (
            O => \N__8930\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__1710\ : Odrv4
    port map (
            O => \N__8925\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__8920\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__1708\ : InMux
    port map (
            O => \N__8909\,
            I => \N__8906\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__8906\,
            I => \N__8903\
        );

    \I__1706\ : Span4Mux_v
    port map (
            O => \N__8903\,
            I => \N__8900\
        );

    \I__1705\ : Odrv4
    port map (
            O => \N__8900\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_1\
        );

    \I__1704\ : CascadeMux
    port map (
            O => \N__8897\,
            I => \N__8894\
        );

    \I__1703\ : InMux
    port map (
            O => \N__8894\,
            I => \N__8891\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__8891\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_1\
        );

    \I__1701\ : InMux
    port map (
            O => \N__8888\,
            I => \N__8885\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8885\,
            I => \N__8882\
        );

    \I__1699\ : Odrv12
    port map (
            O => \N__8882\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1\
        );

    \I__1698\ : CEMux
    port map (
            O => \N__8879\,
            I => \N__8874\
        );

    \I__1697\ : CEMux
    port map (
            O => \N__8878\,
            I => \N__8871\
        );

    \I__1696\ : CEMux
    port map (
            O => \N__8877\,
            I => \N__8868\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__8874\,
            I => \N__8865\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__8871\,
            I => \N__8862\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__8868\,
            I => \N__8859\
        );

    \I__1692\ : Odrv4
    port map (
            O => \N__8865\,
            I => \N_92_i_0\
        );

    \I__1691\ : Odrv4
    port map (
            O => \N__8862\,
            I => \N_92_i_0\
        );

    \I__1690\ : Odrv4
    port map (
            O => \N__8859\,
            I => \N_92_i_0\
        );

    \I__1689\ : SRMux
    port map (
            O => \N__8852\,
            I => \N__8848\
        );

    \I__1688\ : SRMux
    port map (
            O => \N__8851\,
            I => \N__8845\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__8848\,
            I => \N__8841\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__8845\,
            I => \N__8838\
        );

    \I__1685\ : SRMux
    port map (
            O => \N__8844\,
            I => \N__8835\
        );

    \I__1684\ : Span4Mux_h
    port map (
            O => \N__8841\,
            I => \N__8832\
        );

    \I__1683\ : Span4Mux_h
    port map (
            O => \N__8838\,
            I => \N__8829\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__8835\,
            I => \N__8826\
        );

    \I__1681\ : Odrv4
    port map (
            O => \N__8832\,
            I => \rFifoDatarff_0_RNIHJV05\
        );

    \I__1680\ : Odrv4
    port map (
            O => \N__8829\,
            I => \rFifoDatarff_0_RNIHJV05\
        );

    \I__1679\ : Odrv4
    port map (
            O => \N__8826\,
            I => \rFifoDatarff_0_RNIHJV05\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__8819\,
            I => \N__8816\
        );

    \I__1677\ : InMux
    port map (
            O => \N__8816\,
            I => \N__8812\
        );

    \I__1676\ : InMux
    port map (
            O => \N__8815\,
            I => \N__8809\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__8812\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_2\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__8809\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_2\
        );

    \I__1673\ : IoInMux
    port map (
            O => \N__8804\,
            I => \N__8801\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__8801\,
            I => \N__8797\
        );

    \I__1671\ : IoInMux
    port map (
            O => \N__8800\,
            I => \N__8794\
        );

    \I__1670\ : IoSpan4Mux
    port map (
            O => \N__8797\,
            I => \N__8791\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__8794\,
            I => \N__8788\
        );

    \I__1668\ : Span4Mux_s2_v
    port map (
            O => \N__8791\,
            I => \N__8785\
        );

    \I__1667\ : IoSpan4Mux
    port map (
            O => \N__8788\,
            I => \N__8782\
        );

    \I__1666\ : Sp12to4
    port map (
            O => \N__8785\,
            I => \N__8779\
        );

    \I__1665\ : Sp12to4
    port map (
            O => \N__8782\,
            I => \N__8776\
        );

    \I__1664\ : Span12Mux_s8_v
    port map (
            O => \N__8779\,
            I => \N__8770\
        );

    \I__1663\ : Span12Mux_s9_v
    port map (
            O => \N__8776\,
            I => \N__8770\
        );

    \I__1662\ : InMux
    port map (
            O => \N__8775\,
            I => \N__8767\
        );

    \I__1661\ : Odrv12
    port map (
            O => \N__8770\,
            I => \P1A4_c\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__8767\,
            I => \P1A4_c\
        );

    \I__1659\ : InMux
    port map (
            O => \N__8762\,
            I => \N__8756\
        );

    \I__1658\ : InMux
    port map (
            O => \N__8761\,
            I => \N__8756\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__8756\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_3\
        );

    \I__1656\ : IoInMux
    port map (
            O => \N__8753\,
            I => \N__8747\
        );

    \I__1655\ : IoInMux
    port map (
            O => \N__8752\,
            I => \N__8744\
        );

    \I__1654\ : IoInMux
    port map (
            O => \N__8751\,
            I => \N__8740\
        );

    \I__1653\ : IoInMux
    port map (
            O => \N__8750\,
            I => \N__8737\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__8747\,
            I => \N__8732\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__8744\,
            I => \N__8732\
        );

    \I__1650\ : IoInMux
    port map (
            O => \N__8743\,
            I => \N__8729\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__8740\,
            I => \N__8723\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__8737\,
            I => \N__8723\
        );

    \I__1647\ : IoSpan4Mux
    port map (
            O => \N__8732\,
            I => \N__8717\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__8729\,
            I => \N__8717\
        );

    \I__1645\ : IoInMux
    port map (
            O => \N__8728\,
            I => \N__8714\
        );

    \I__1644\ : Span4Mux_s2_v
    port map (
            O => \N__8723\,
            I => \N__8711\
        );

    \I__1643\ : IoInMux
    port map (
            O => \N__8722\,
            I => \N__8708\
        );

    \I__1642\ : IoSpan4Mux
    port map (
            O => \N__8717\,
            I => \N__8705\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__8714\,
            I => \N__8702\
        );

    \I__1640\ : Span4Mux_h
    port map (
            O => \N__8711\,
            I => \N__8699\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__8708\,
            I => \N__8695\
        );

    \I__1638\ : Span4Mux_s3_v
    port map (
            O => \N__8705\,
            I => \N__8692\
        );

    \I__1637\ : Span4Mux_s3_v
    port map (
            O => \N__8702\,
            I => \N__8689\
        );

    \I__1636\ : Span4Mux_v
    port map (
            O => \N__8699\,
            I => \N__8686\
        );

    \I__1635\ : IoInMux
    port map (
            O => \N__8698\,
            I => \N__8683\
        );

    \I__1634\ : Span4Mux_s3_v
    port map (
            O => \N__8695\,
            I => \N__8680\
        );

    \I__1633\ : Sp12to4
    port map (
            O => \N__8692\,
            I => \N__8674\
        );

    \I__1632\ : Sp12to4
    port map (
            O => \N__8689\,
            I => \N__8674\
        );

    \I__1631\ : Sp12to4
    port map (
            O => \N__8686\,
            I => \N__8671\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__8683\,
            I => \N__8668\
        );

    \I__1629\ : Span4Mux_v
    port map (
            O => \N__8680\,
            I => \N__8665\
        );

    \I__1628\ : CascadeMux
    port map (
            O => \N__8679\,
            I => \N__8662\
        );

    \I__1627\ : Span12Mux_h
    port map (
            O => \N__8674\,
            I => \N__8659\
        );

    \I__1626\ : Span12Mux_v
    port map (
            O => \N__8671\,
            I => \N__8654\
        );

    \I__1625\ : Span12Mux_s11_v
    port map (
            O => \N__8668\,
            I => \N__8654\
        );

    \I__1624\ : Span4Mux_v
    port map (
            O => \N__8665\,
            I => \N__8651\
        );

    \I__1623\ : InMux
    port map (
            O => \N__8662\,
            I => \N__8648\
        );

    \I__1622\ : Odrv12
    port map (
            O => \N__8659\,
            I => \rTxBusReady\
        );

    \I__1621\ : Odrv12
    port map (
            O => \N__8654\,
            I => \rTxBusReady\
        );

    \I__1620\ : Odrv4
    port map (
            O => \N__8651\,
            I => \rTxBusReady\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__8648\,
            I => \rTxBusReady\
        );

    \I__1618\ : InMux
    port map (
            O => \N__8639\,
            I => \N__8632\
        );

    \I__1617\ : InMux
    port map (
            O => \N__8638\,
            I => \N__8623\
        );

    \I__1616\ : InMux
    port map (
            O => \N__8637\,
            I => \N__8623\
        );

    \I__1615\ : InMux
    port map (
            O => \N__8636\,
            I => \N__8623\
        );

    \I__1614\ : InMux
    port map (
            O => \N__8635\,
            I => \N__8623\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__8632\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_4\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__8623\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_4\
        );

    \I__1611\ : CascadeMux
    port map (
            O => \N__8618\,
            I => \N__8614\
        );

    \I__1610\ : CascadeMux
    port map (
            O => \N__8617\,
            I => \N__8609\
        );

    \I__1609\ : InMux
    port map (
            O => \N__8614\,
            I => \N__8601\
        );

    \I__1608\ : InMux
    port map (
            O => \N__8613\,
            I => \N__8601\
        );

    \I__1607\ : InMux
    port map (
            O => \N__8612\,
            I => \N__8601\
        );

    \I__1606\ : InMux
    port map (
            O => \N__8609\,
            I => \N__8596\
        );

    \I__1605\ : InMux
    port map (
            O => \N__8608\,
            I => \N__8596\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__8601\,
            I => \fifo_inst.ft2232h_inst.rTxRdEnZ0\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__8596\,
            I => \fifo_inst.ft2232h_inst.rTxRdEnZ0\
        );

    \I__1602\ : InMux
    port map (
            O => \N__8591\,
            I => \N__8586\
        );

    \I__1601\ : InMux
    port map (
            O => \N__8590\,
            I => \N__8581\
        );

    \I__1600\ : InMux
    port map (
            O => \N__8589\,
            I => \N__8581\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__8586\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_1\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__8581\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_1\
        );

    \I__1597\ : InMux
    port map (
            O => \N__8576\,
            I => \N__8571\
        );

    \I__1596\ : InMux
    port map (
            O => \N__8575\,
            I => \N__8563\
        );

    \I__1595\ : InMux
    port map (
            O => \N__8574\,
            I => \N__8563\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__8571\,
            I => \N__8560\
        );

    \I__1593\ : CascadeMux
    port map (
            O => \N__8570\,
            I => \N__8557\
        );

    \I__1592\ : InMux
    port map (
            O => \N__8569\,
            I => \N__8552\
        );

    \I__1591\ : InMux
    port map (
            O => \N__8568\,
            I => \N__8552\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__8563\,
            I => \N__8549\
        );

    \I__1589\ : Span4Mux_v
    port map (
            O => \N__8560\,
            I => \N__8546\
        );

    \I__1588\ : InMux
    port map (
            O => \N__8557\,
            I => \N__8543\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__8552\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_0\
        );

    \I__1586\ : Odrv12
    port map (
            O => \N__8549\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_0\
        );

    \I__1585\ : Odrv4
    port map (
            O => \N__8546\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_0\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__8543\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_0\
        );

    \I__1583\ : InMux
    port map (
            O => \N__8534\,
            I => \N__8525\
        );

    \I__1582\ : InMux
    port map (
            O => \N__8533\,
            I => \N__8525\
        );

    \I__1581\ : InMux
    port map (
            O => \N__8532\,
            I => \N__8522\
        );

    \I__1580\ : InMux
    port map (
            O => \N__8531\,
            I => \N__8519\
        );

    \I__1579\ : InMux
    port map (
            O => \N__8530\,
            I => \N__8516\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__8525\,
            I => \N__8511\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__8522\,
            I => \N__8511\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__8519\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_1\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__8516\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_1\
        );

    \I__1574\ : Odrv4
    port map (
            O => \N__8511\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_1\
        );

    \I__1573\ : CascadeMux
    port map (
            O => \N__8504\,
            I => \DUT.fifo_tx_inst.N_83_cascade_\
        );

    \I__1572\ : InMux
    port map (
            O => \N__8501\,
            I => \N__8498\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__8498\,
            I => \DUT.fifo_tx_inst.N_88\
        );

    \I__1570\ : CascadeMux
    port map (
            O => \N__8495\,
            I => \DUT.fifo_tx_inst.N_88_cascade_\
        );

    \I__1569\ : InMux
    port map (
            O => \N__8492\,
            I => \N__8489\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__8489\,
            I => \DUT.rTransmitc\
        );

    \I__1567\ : InMux
    port map (
            O => \N__8486\,
            I => \N__8480\
        );

    \I__1566\ : InMux
    port map (
            O => \N__8485\,
            I => \N__8480\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__8480\,
            I => \N__8477\
        );

    \I__1564\ : Span4Mux_v
    port map (
            O => \N__8477\,
            I => \N__8471\
        );

    \I__1563\ : InMux
    port map (
            O => \N__8476\,
            I => \N__8466\
        );

    \I__1562\ : InMux
    port map (
            O => \N__8475\,
            I => \N__8466\
        );

    \I__1561\ : InMux
    port map (
            O => \N__8474\,
            I => \N__8463\
        );

    \I__1560\ : Odrv4
    port map (
            O => \N__8471\,
            I => \DUT.fifo_tx_inst.rWritePtr16\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__8466\,
            I => \DUT.fifo_tx_inst.rWritePtr16\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__8463\,
            I => \DUT.fifo_tx_inst.rWritePtr16\
        );

    \I__1557\ : InMux
    port map (
            O => \N__8456\,
            I => \N__8453\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__8453\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_3\
        );

    \I__1555\ : InMux
    port map (
            O => \N__8450\,
            I => \N__8446\
        );

    \I__1554\ : InMux
    port map (
            O => \N__8449\,
            I => \N__8443\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__8446\,
            I => \DUT.fifo_tx_inst.rFifoDataro_0\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__8443\,
            I => \DUT.fifo_tx_inst.rFifoDataro_0\
        );

    \I__1551\ : CascadeMux
    port map (
            O => \N__8438\,
            I => \N__8434\
        );

    \I__1550\ : InMux
    port map (
            O => \N__8437\,
            I => \N__8431\
        );

    \I__1549\ : InMux
    port map (
            O => \N__8434\,
            I => \N__8428\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__8431\,
            I => \DUT.fifo_tx_inst.rFifoDataro_1\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__8428\,
            I => \DUT.fifo_tx_inst.rFifoDataro_1\
        );

    \I__1546\ : CascadeMux
    port map (
            O => \N__8423\,
            I => \N__8420\
        );

    \I__1545\ : InMux
    port map (
            O => \N__8420\,
            I => \N__8417\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__8417\,
            I => \DUT.rFifoDataror_1\
        );

    \I__1543\ : CascadeMux
    port map (
            O => \N__8414\,
            I => \DUT.rFifoDataror_1_cascade_\
        );

    \I__1542\ : InMux
    port map (
            O => \N__8411\,
            I => \N__8408\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__8408\,
            I => \N__8404\
        );

    \I__1540\ : InMux
    port map (
            O => \N__8407\,
            I => \N__8401\
        );

    \I__1539\ : Odrv4
    port map (
            O => \N__8404\,
            I => \DUT.rFifoDataror_0_0\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__8401\,
            I => \DUT.rFifoDataror_0_0\
        );

    \I__1537\ : CascadeMux
    port map (
            O => \N__8396\,
            I => \N__8392\
        );

    \I__1536\ : InMux
    port map (
            O => \N__8395\,
            I => \N__8382\
        );

    \I__1535\ : InMux
    port map (
            O => \N__8392\,
            I => \N__8382\
        );

    \I__1534\ : InMux
    port map (
            O => \N__8391\,
            I => \N__8371\
        );

    \I__1533\ : InMux
    port map (
            O => \N__8390\,
            I => \N__8371\
        );

    \I__1532\ : InMux
    port map (
            O => \N__8389\,
            I => \N__8371\
        );

    \I__1531\ : InMux
    port map (
            O => \N__8388\,
            I => \N__8371\
        );

    \I__1530\ : InMux
    port map (
            O => \N__8387\,
            I => \N__8371\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__8382\,
            I => \N__8366\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__8371\,
            I => \N__8366\
        );

    \I__1527\ : Odrv4
    port map (
            O => \N__8366\,
            I => \DUT.rFifoDataror_0\
        );

    \I__1526\ : IoInMux
    port map (
            O => \N__8363\,
            I => \N__8359\
        );

    \I__1525\ : CascadeMux
    port map (
            O => \N__8362\,
            I => \N__8354\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__8359\,
            I => \N__8349\
        );

    \I__1523\ : InMux
    port map (
            O => \N__8358\,
            I => \N__8343\
        );

    \I__1522\ : InMux
    port map (
            O => \N__8357\,
            I => \N__8343\
        );

    \I__1521\ : InMux
    port map (
            O => \N__8354\,
            I => \N__8340\
        );

    \I__1520\ : InMux
    port map (
            O => \N__8353\,
            I => \N__8337\
        );

    \I__1519\ : InMux
    port map (
            O => \N__8352\,
            I => \N__8333\
        );

    \I__1518\ : Span4Mux_s1_v
    port map (
            O => \N__8349\,
            I => \N__8329\
        );

    \I__1517\ : CascadeMux
    port map (
            O => \N__8348\,
            I => \N__8325\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__8343\,
            I => \N__8320\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__8340\,
            I => \N__8320\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__8337\,
            I => \N__8317\
        );

    \I__1513\ : InMux
    port map (
            O => \N__8336\,
            I => \N__8314\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__8333\,
            I => \N__8311\
        );

    \I__1511\ : InMux
    port map (
            O => \N__8332\,
            I => \N__8308\
        );

    \I__1510\ : Sp12to4
    port map (
            O => \N__8329\,
            I => \N__8305\
        );

    \I__1509\ : InMux
    port map (
            O => \N__8328\,
            I => \N__8300\
        );

    \I__1508\ : InMux
    port map (
            O => \N__8325\,
            I => \N__8300\
        );

    \I__1507\ : Span4Mux_v
    port map (
            O => \N__8320\,
            I => \N__8293\
        );

    \I__1506\ : Span4Mux_v
    port map (
            O => \N__8317\,
            I => \N__8293\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__8314\,
            I => \N__8293\
        );

    \I__1504\ : Span4Mux_h
    port map (
            O => \N__8311\,
            I => \N__8290\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__8308\,
            I => \N__8287\
        );

    \I__1502\ : Span12Mux_h
    port map (
            O => \N__8305\,
            I => \N__8284\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__8300\,
            I => \N__8281\
        );

    \I__1500\ : Span4Mux_v
    port map (
            O => \N__8293\,
            I => \N__8278\
        );

    \I__1499\ : Span4Mux_v
    port map (
            O => \N__8290\,
            I => \N__8273\
        );

    \I__1498\ : Span4Mux_h
    port map (
            O => \N__8287\,
            I => \N__8273\
        );

    \I__1497\ : Span12Mux_v
    port map (
            O => \N__8284\,
            I => \N__8268\
        );

    \I__1496\ : Span12Mux_h
    port map (
            O => \N__8281\,
            I => \N__8268\
        );

    \I__1495\ : Sp12to4
    port map (
            O => \N__8278\,
            I => \N__8265\
        );

    \I__1494\ : Sp12to4
    port map (
            O => \N__8273\,
            I => \N__8262\
        );

    \I__1493\ : Span12Mux_v
    port map (
            O => \N__8268\,
            I => \N__8259\
        );

    \I__1492\ : Span12Mux_h
    port map (
            O => \N__8265\,
            I => \N__8256\
        );

    \I__1491\ : Span12Mux_v
    port map (
            O => \N__8262\,
            I => \N__8253\
        );

    \I__1490\ : Odrv12
    port map (
            O => \N__8259\,
            I => \wPllLocked\
        );

    \I__1489\ : Odrv12
    port map (
            O => \N__8256\,
            I => \wPllLocked\
        );

    \I__1488\ : Odrv12
    port map (
            O => \N__8253\,
            I => \wPllLocked\
        );

    \I__1487\ : InMux
    port map (
            O => \N__8246\,
            I => \N__8240\
        );

    \I__1486\ : InMux
    port map (
            O => \N__8245\,
            I => \N__8240\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__8240\,
            I => \DUT.fifo_rx_inst.CO0\
        );

    \I__1484\ : InMux
    port map (
            O => \N__8237\,
            I => \N__8234\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__8234\,
            I => \DUT.fifo_rx_inst.un1_i11_2_i\
        );

    \I__1482\ : CascadeMux
    port map (
            O => \N__8231\,
            I => \DUT.fifo_rx_inst.un1_i11_2_i_cascade_\
        );

    \I__1481\ : InMux
    port map (
            O => \N__8228\,
            I => \N__8224\
        );

    \I__1480\ : InMux
    port map (
            O => \N__8227\,
            I => \N__8218\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__8224\,
            I => \N__8215\
        );

    \I__1478\ : InMux
    port map (
            O => \N__8223\,
            I => \N__8210\
        );

    \I__1477\ : InMux
    port map (
            O => \N__8222\,
            I => \N__8210\
        );

    \I__1476\ : InMux
    port map (
            O => \N__8221\,
            I => \N__8207\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__8218\,
            I => \DUT.fifo_rx_inst.N_92\
        );

    \I__1474\ : Odrv4
    port map (
            O => \N__8215\,
            I => \DUT.fifo_rx_inst.N_92\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__8210\,
            I => \DUT.fifo_rx_inst.N_92\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__8207\,
            I => \DUT.fifo_rx_inst.N_92\
        );

    \I__1471\ : InMux
    port map (
            O => \N__8198\,
            I => \N__8183\
        );

    \I__1470\ : InMux
    port map (
            O => \N__8197\,
            I => \N__8183\
        );

    \I__1469\ : InMux
    port map (
            O => \N__8196\,
            I => \N__8183\
        );

    \I__1468\ : InMux
    port map (
            O => \N__8195\,
            I => \N__8183\
        );

    \I__1467\ : InMux
    port map (
            O => \N__8194\,
            I => \N__8177\
        );

    \I__1466\ : InMux
    port map (
            O => \N__8193\,
            I => \N__8177\
        );

    \I__1465\ : InMux
    port map (
            O => \N__8192\,
            I => \N__8173\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__8183\,
            I => \N__8170\
        );

    \I__1463\ : InMux
    port map (
            O => \N__8182\,
            I => \N__8167\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__8177\,
            I => \N__8164\
        );

    \I__1461\ : InMux
    port map (
            O => \N__8176\,
            I => \N__8158\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__8173\,
            I => \N__8155\
        );

    \I__1459\ : Span4Mux_v
    port map (
            O => \N__8170\,
            I => \N__8150\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__8167\,
            I => \N__8150\
        );

    \I__1457\ : Span4Mux_h
    port map (
            O => \N__8164\,
            I => \N__8147\
        );

    \I__1456\ : InMux
    port map (
            O => \N__8163\,
            I => \N__8144\
        );

    \I__1455\ : InMux
    port map (
            O => \N__8162\,
            I => \N__8139\
        );

    \I__1454\ : InMux
    port map (
            O => \N__8161\,
            I => \N__8139\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__8158\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__1452\ : Odrv4
    port map (
            O => \N__8155\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__1451\ : Odrv4
    port map (
            O => \N__8150\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__1450\ : Odrv4
    port map (
            O => \N__8147\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__8144\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__8139\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__1447\ : CascadeMux
    port map (
            O => \N__8126\,
            I => \DUT.uart_inst0.N_79_cascade_\
        );

    \I__1446\ : InMux
    port map (
            O => \N__8123\,
            I => \N__8120\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__8120\,
            I => \N__8117\
        );

    \I__1444\ : Odrv12
    port map (
            O => \N__8117\,
            I => \DUT.uart_inst0.tx_state_ns_i_i_0_0\
        );

    \I__1443\ : CascadeMux
    port map (
            O => \N__8114\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_\
        );

    \I__1442\ : InMux
    port map (
            O => \N__8111\,
            I => \N__8108\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__8108\,
            I => \N__8105\
        );

    \I__1440\ : Span4Mux_h
    port map (
            O => \N__8105\,
            I => \N__8102\
        );

    \I__1439\ : Odrv4
    port map (
            O => \N__8102\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_2\
        );

    \I__1438\ : InMux
    port map (
            O => \N__8099\,
            I => \N__8096\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__8096\,
            I => \N__8093\
        );

    \I__1436\ : Odrv4
    port map (
            O => \N__8093\,
            I => \DUT.rFifoDatarx_2\
        );

    \I__1435\ : InMux
    port map (
            O => \N__8090\,
            I => \N__8087\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__8087\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_2\
        );

    \I__1433\ : InMux
    port map (
            O => \N__8084\,
            I => \N__8081\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__8081\,
            I => \N__8078\
        );

    \I__1431\ : Span4Mux_h
    port map (
            O => \N__8078\,
            I => \N__8075\
        );

    \I__1430\ : Odrv4
    port map (
            O => \N__8075\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_3\
        );

    \I__1429\ : CascadeMux
    port map (
            O => \N__8072\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_\
        );

    \I__1428\ : InMux
    port map (
            O => \N__8069\,
            I => \N__8066\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__8066\,
            I => \N__8063\
        );

    \I__1426\ : Odrv4
    port map (
            O => \N__8063\,
            I => \DUT.rFifoDatarx_3\
        );

    \I__1425\ : CascadeMux
    port map (
            O => \N__8060\,
            I => \N__8057\
        );

    \I__1424\ : InMux
    port map (
            O => \N__8057\,
            I => \N__8054\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__8054\,
            I => \DUT.uart_inst0.tx_dataZ0Z_1\
        );

    \I__1422\ : InMux
    port map (
            O => \N__8051\,
            I => \N__8048\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__8048\,
            I => \DUT.uart_inst0.tx_dataZ0Z_2\
        );

    \I__1420\ : InMux
    port map (
            O => \N__8045\,
            I => \N__8042\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__8042\,
            I => \DUT.uart_inst0.tx_dataZ0Z_3\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__8039\,
            I => \N__8036\
        );

    \I__1417\ : InMux
    port map (
            O => \N__8036\,
            I => \N__8033\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__8033\,
            I => \DUT.uart_inst0.tx_dataZ0Z_4\
        );

    \I__1415\ : InMux
    port map (
            O => \N__8030\,
            I => \N__8027\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__8027\,
            I => \N__8024\
        );

    \I__1413\ : Odrv4
    port map (
            O => \N__8024\,
            I => \DUT.uart_inst0.tx_dataZ0Z_5\
        );

    \I__1412\ : CascadeMux
    port map (
            O => \N__8021\,
            I => \N__8018\
        );

    \I__1411\ : InMux
    port map (
            O => \N__8018\,
            I => \N__8015\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__8015\,
            I => \DUT.uart_inst0.tx_dataZ0Z_6\
        );

    \I__1409\ : InMux
    port map (
            O => \N__8012\,
            I => \N__8009\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__8009\,
            I => \N__8006\
        );

    \I__1407\ : Odrv4
    port map (
            O => \N__8006\,
            I => \DUT.uart_inst0.tx_dataZ0Z_7\
        );

    \I__1406\ : CEMux
    port map (
            O => \N__8003\,
            I => \N__7999\
        );

    \I__1405\ : CEMux
    port map (
            O => \N__8002\,
            I => \N__7996\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__7999\,
            I => \N__7993\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__7996\,
            I => \N__7990\
        );

    \I__1402\ : Span4Mux_h
    port map (
            O => \N__7993\,
            I => \N__7987\
        );

    \I__1401\ : Odrv4
    port map (
            O => \N__7990\,
            I => \DUT.uart_inst0.N_22_i\
        );

    \I__1400\ : Odrv4
    port map (
            O => \N__7987\,
            I => \DUT.uart_inst0.N_22_i\
        );

    \I__1399\ : CascadeMux
    port map (
            O => \N__7982\,
            I => \DUT.uart_inst0.g0_i_o6_0_4_cascade_\
        );

    \I__1398\ : InMux
    port map (
            O => \N__7979\,
            I => \N__7976\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__7976\,
            I => \DUT.uart_inst0.g0_i_o6_0_5\
        );

    \I__1396\ : CascadeMux
    port map (
            O => \N__7973\,
            I => \DUT.uart_inst0.N_139_0_cascade_\
        );

    \I__1395\ : InMux
    port map (
            O => \N__7970\,
            I => \N__7967\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__7967\,
            I => \DUT.uart_inst0.tx_bits_remaining_RNO_1Z0Z_3\
        );

    \I__1393\ : InMux
    port map (
            O => \N__7964\,
            I => \N__7961\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__7961\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_9\
        );

    \I__1391\ : InMux
    port map (
            O => \N__7958\,
            I => \N__7955\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__7955\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_13\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__7952\,
            I => \DUT.uart_inst0.un1_N_5_mux_cascade_\
        );

    \I__1388\ : InMux
    port map (
            O => \N__7949\,
            I => \N__7946\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__7946\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_1\
        );

    \I__1386\ : InMux
    port map (
            O => \N__7943\,
            I => \N__7940\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__7940\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_10\
        );

    \I__1384\ : InMux
    port map (
            O => \N__7937\,
            I => \N__7930\
        );

    \I__1383\ : InMux
    port map (
            O => \N__7936\,
            I => \N__7930\
        );

    \I__1382\ : InMux
    port map (
            O => \N__7935\,
            I => \N__7927\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__7930\,
            I => \N__7914\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__7927\,
            I => \N__7910\
        );

    \I__1379\ : InMux
    port map (
            O => \N__7926\,
            I => \N__7907\
        );

    \I__1378\ : InMux
    port map (
            O => \N__7925\,
            I => \N__7904\
        );

    \I__1377\ : InMux
    port map (
            O => \N__7924\,
            I => \N__7901\
        );

    \I__1376\ : CascadeMux
    port map (
            O => \N__7923\,
            I => \N__7896\
        );

    \I__1375\ : InMux
    port map (
            O => \N__7922\,
            I => \N__7888\
        );

    \I__1374\ : InMux
    port map (
            O => \N__7921\,
            I => \N__7888\
        );

    \I__1373\ : InMux
    port map (
            O => \N__7920\,
            I => \N__7881\
        );

    \I__1372\ : InMux
    port map (
            O => \N__7919\,
            I => \N__7881\
        );

    \I__1371\ : InMux
    port map (
            O => \N__7918\,
            I => \N__7881\
        );

    \I__1370\ : InMux
    port map (
            O => \N__7917\,
            I => \N__7878\
        );

    \I__1369\ : Span4Mux_h
    port map (
            O => \N__7914\,
            I => \N__7875\
        );

    \I__1368\ : InMux
    port map (
            O => \N__7913\,
            I => \N__7872\
        );

    \I__1367\ : Span4Mux_h
    port map (
            O => \N__7910\,
            I => \N__7863\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__7907\,
            I => \N__7863\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__7904\,
            I => \N__7863\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__7901\,
            I => \N__7863\
        );

    \I__1363\ : InMux
    port map (
            O => \N__7900\,
            I => \N__7858\
        );

    \I__1362\ : InMux
    port map (
            O => \N__7899\,
            I => \N__7858\
        );

    \I__1361\ : InMux
    port map (
            O => \N__7896\,
            I => \N__7851\
        );

    \I__1360\ : InMux
    port map (
            O => \N__7895\,
            I => \N__7851\
        );

    \I__1359\ : InMux
    port map (
            O => \N__7894\,
            I => \N__7851\
        );

    \I__1358\ : InMux
    port map (
            O => \N__7893\,
            I => \N__7848\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__7888\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__7881\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__7878\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__1354\ : Odrv4
    port map (
            O => \N__7875\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__7872\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__1352\ : Odrv4
    port map (
            O => \N__7863\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__7858\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__7851\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__7848\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__1348\ : InMux
    port map (
            O => \N__7829\,
            I => \N__7826\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__7826\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_11\
        );

    \I__1346\ : CascadeMux
    port map (
            O => \N__7823\,
            I => \N__7820\
        );

    \I__1345\ : InMux
    port map (
            O => \N__7820\,
            I => \N__7817\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__7817\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_12\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7814\,
            I => \N__7811\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__7811\,
            I => \N__7806\
        );

    \I__1341\ : InMux
    port map (
            O => \N__7810\,
            I => \N__7803\
        );

    \I__1340\ : InMux
    port map (
            O => \N__7809\,
            I => \N__7799\
        );

    \I__1339\ : Span4Mux_v
    port map (
            O => \N__7806\,
            I => \N__7794\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__7803\,
            I => \N__7794\
        );

    \I__1337\ : InMux
    port map (
            O => \N__7802\,
            I => \N__7791\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__7799\,
            I => \N__7788\
        );

    \I__1335\ : Span4Mux_v
    port map (
            O => \N__7794\,
            I => \N__7784\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__7791\,
            I => \N__7781\
        );

    \I__1333\ : Span4Mux_h
    port map (
            O => \N__7788\,
            I => \N__7778\
        );

    \I__1332\ : InMux
    port map (
            O => \N__7787\,
            I => \N__7775\
        );

    \I__1331\ : Odrv4
    port map (
            O => \N__7784\,
            I => \DUT.wRxByte_3\
        );

    \I__1330\ : Odrv12
    port map (
            O => \N__7781\,
            I => \DUT.wRxByte_3\
        );

    \I__1329\ : Odrv4
    port map (
            O => \N__7778\,
            I => \DUT.wRxByte_3\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__7775\,
            I => \DUT.wRxByte_3\
        );

    \I__1327\ : InMux
    port map (
            O => \N__7766\,
            I => \N__7763\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__7763\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_3\
        );

    \I__1325\ : InMux
    port map (
            O => \N__7760\,
            I => \N__7755\
        );

    \I__1324\ : InMux
    port map (
            O => \N__7759\,
            I => \N__7751\
        );

    \I__1323\ : InMux
    port map (
            O => \N__7758\,
            I => \N__7748\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__7755\,
            I => \N__7745\
        );

    \I__1321\ : InMux
    port map (
            O => \N__7754\,
            I => \N__7742\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__7751\,
            I => \N__7739\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__7748\,
            I => \N__7732\
        );

    \I__1318\ : Span4Mux_h
    port map (
            O => \N__7745\,
            I => \N__7732\
        );

    \I__1317\ : LocalMux
    port map (
            O => \N__7742\,
            I => \N__7732\
        );

    \I__1316\ : Span4Mux_v
    port map (
            O => \N__7739\,
            I => \N__7728\
        );

    \I__1315\ : Span4Mux_v
    port map (
            O => \N__7732\,
            I => \N__7725\
        );

    \I__1314\ : InMux
    port map (
            O => \N__7731\,
            I => \N__7722\
        );

    \I__1313\ : Odrv4
    port map (
            O => \N__7728\,
            I => \DUT.wRxByte_4\
        );

    \I__1312\ : Odrv4
    port map (
            O => \N__7725\,
            I => \DUT.wRxByte_4\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__7722\,
            I => \DUT.wRxByte_4\
        );

    \I__1310\ : InMux
    port map (
            O => \N__7715\,
            I => \N__7712\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__7712\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_4\
        );

    \I__1308\ : InMux
    port map (
            O => \N__7709\,
            I => \N__7704\
        );

    \I__1307\ : InMux
    port map (
            O => \N__7708\,
            I => \N__7700\
        );

    \I__1306\ : InMux
    port map (
            O => \N__7707\,
            I => \N__7697\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__7704\,
            I => \N__7694\
        );

    \I__1304\ : InMux
    port map (
            O => \N__7703\,
            I => \N__7691\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__7700\,
            I => \N__7688\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__7697\,
            I => \N__7681\
        );

    \I__1301\ : Span4Mux_h
    port map (
            O => \N__7694\,
            I => \N__7681\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__7691\,
            I => \N__7681\
        );

    \I__1299\ : Span4Mux_v
    port map (
            O => \N__7688\,
            I => \N__7677\
        );

    \I__1298\ : Span4Mux_v
    port map (
            O => \N__7681\,
            I => \N__7674\
        );

    \I__1297\ : InMux
    port map (
            O => \N__7680\,
            I => \N__7671\
        );

    \I__1296\ : Odrv4
    port map (
            O => \N__7677\,
            I => \DUT.wRxByte_5\
        );

    \I__1295\ : Odrv4
    port map (
            O => \N__7674\,
            I => \DUT.wRxByte_5\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__7671\,
            I => \DUT.wRxByte_5\
        );

    \I__1293\ : InMux
    port map (
            O => \N__7664\,
            I => \N__7661\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__7661\,
            I => \N__7658\
        );

    \I__1291\ : Odrv4
    port map (
            O => \N__7658\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_5\
        );

    \I__1290\ : InMux
    port map (
            O => \N__7655\,
            I => \N__7649\
        );

    \I__1289\ : InMux
    port map (
            O => \N__7654\,
            I => \N__7646\
        );

    \I__1288\ : InMux
    port map (
            O => \N__7653\,
            I => \N__7643\
        );

    \I__1287\ : InMux
    port map (
            O => \N__7652\,
            I => \N__7640\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__7649\,
            I => \N__7637\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__7646\,
            I => \N__7632\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__7643\,
            I => \N__7632\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__7640\,
            I => \N__7629\
        );

    \I__1282\ : Span4Mux_h
    port map (
            O => \N__7637\,
            I => \N__7625\
        );

    \I__1281\ : Span4Mux_v
    port map (
            O => \N__7632\,
            I => \N__7620\
        );

    \I__1280\ : Span4Mux_h
    port map (
            O => \N__7629\,
            I => \N__7620\
        );

    \I__1279\ : InMux
    port map (
            O => \N__7628\,
            I => \N__7617\
        );

    \I__1278\ : Odrv4
    port map (
            O => \N__7625\,
            I => \DUT.wRxByte_6\
        );

    \I__1277\ : Odrv4
    port map (
            O => \N__7620\,
            I => \DUT.wRxByte_6\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__7617\,
            I => \DUT.wRxByte_6\
        );

    \I__1275\ : InMux
    port map (
            O => \N__7610\,
            I => \N__7607\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__7607\,
            I => \N__7604\
        );

    \I__1273\ : Span4Mux_v
    port map (
            O => \N__7604\,
            I => \N__7601\
        );

    \I__1272\ : Odrv4
    port map (
            O => \N__7601\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_6\
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__7598\,
            I => \N__7595\
        );

    \I__1270\ : InMux
    port map (
            O => \N__7595\,
            I => \N__7592\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__7592\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_7\
        );

    \I__1268\ : CEMux
    port map (
            O => \N__7589\,
            I => \N__7586\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__7586\,
            I => \N__7582\
        );

    \I__1266\ : InMux
    port map (
            O => \N__7585\,
            I => \N__7579\
        );

    \I__1265\ : Span4Mux_v
    port map (
            O => \N__7582\,
            I => \N__7576\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__7579\,
            I => \N__7573\
        );

    \I__1263\ : Span4Mux_h
    port map (
            O => \N__7576\,
            I => \N__7570\
        );

    \I__1262\ : Span4Mux_h
    port map (
            O => \N__7573\,
            I => \N__7567\
        );

    \I__1261\ : Odrv4
    port map (
            O => \N__7570\,
            I => \DUT.fifo_rx_inst.rFifoData_awe3\
        );

    \I__1260\ : Odrv4
    port map (
            O => \N__7567\,
            I => \DUT.fifo_rx_inst.rFifoData_awe3\
        );

    \I__1259\ : InMux
    port map (
            O => \N__7562\,
            I => \N__7559\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__7559\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_7\
        );

    \I__1257\ : InMux
    port map (
            O => \N__7556\,
            I => \N__7553\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__7553\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7\
        );

    \I__1255\ : IoInMux
    port map (
            O => \N__7550\,
            I => \N__7547\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__7547\,
            I => \N__7543\
        );

    \I__1253\ : IoInMux
    port map (
            O => \N__7546\,
            I => \N__7540\
        );

    \I__1252\ : IoSpan4Mux
    port map (
            O => \N__7543\,
            I => \N__7537\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__7540\,
            I => \N__7534\
        );

    \I__1250\ : IoSpan4Mux
    port map (
            O => \N__7537\,
            I => \N__7531\
        );

    \I__1249\ : Span4Mux_s3_v
    port map (
            O => \N__7534\,
            I => \N__7528\
        );

    \I__1248\ : Span4Mux_s3_v
    port map (
            O => \N__7531\,
            I => \N__7523\
        );

    \I__1247\ : Span4Mux_h
    port map (
            O => \N__7528\,
            I => \N__7523\
        );

    \I__1246\ : Sp12to4
    port map (
            O => \N__7523\,
            I => \N__7519\
        );

    \I__1245\ : InMux
    port map (
            O => \N__7522\,
            I => \N__7516\
        );

    \I__1244\ : Odrv12
    port map (
            O => \N__7519\,
            I => \P1A3_c\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__7516\,
            I => \P1A3_c\
        );

    \I__1242\ : CEMux
    port map (
            O => \N__7511\,
            I => \N__7508\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__7508\,
            I => \N__7504\
        );

    \I__1240\ : InMux
    port map (
            O => \N__7507\,
            I => \N__7501\
        );

    \I__1239\ : Odrv12
    port map (
            O => \N__7504\,
            I => \DUT.fifo_rx_inst.rFifoData_awe1\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__7501\,
            I => \DUT.fifo_rx_inst.rFifoData_awe1\
        );

    \I__1237\ : InMux
    port map (
            O => \N__7496\,
            I => \N__7490\
        );

    \I__1236\ : InMux
    port map (
            O => \N__7495\,
            I => \N__7490\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__7490\,
            I => \DUT.fifo_rx_inst.rFifoDataro_1\
        );

    \I__1234\ : CEMux
    port map (
            O => \N__7487\,
            I => \N__7484\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__7484\,
            I => \N__7481\
        );

    \I__1232\ : Span4Mux_h
    port map (
            O => \N__7481\,
            I => \N__7477\
        );

    \I__1231\ : InMux
    port map (
            O => \N__7480\,
            I => \N__7474\
        );

    \I__1230\ : Odrv4
    port map (
            O => \N__7477\,
            I => \DUT.fifo_rx_inst.rFifoData_awe2\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__7474\,
            I => \DUT.fifo_rx_inst.rFifoData_awe2\
        );

    \I__1228\ : InMux
    port map (
            O => \N__7469\,
            I => \N__7463\
        );

    \I__1227\ : InMux
    port map (
            O => \N__7468\,
            I => \N__7463\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__7463\,
            I => \DUT.fifo_rx_inst.rFifoDataro_3\
        );

    \I__1225\ : CascadeMux
    port map (
            O => \N__7460\,
            I => \N__7456\
        );

    \I__1224\ : InMux
    port map (
            O => \N__7459\,
            I => \N__7451\
        );

    \I__1223\ : InMux
    port map (
            O => \N__7456\,
            I => \N__7451\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__7451\,
            I => \DUT.fifo_rx_inst.rFifoDataro_2\
        );

    \I__1221\ : InMux
    port map (
            O => \N__7448\,
            I => \N__7445\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__7445\,
            I => \DUT.fifo_rx_inst.rTxByte_42_1\
        );

    \I__1219\ : CascadeMux
    port map (
            O => \N__7442\,
            I => \DUT.fifo_rx_inst.rTxByte_42_0_cascade_\
        );

    \I__1218\ : InMux
    port map (
            O => \N__7439\,
            I => \N__7436\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__7436\,
            I => \N__7433\
        );

    \I__1216\ : Odrv4
    port map (
            O => \N__7433\,
            I => \N_92_i\
        );

    \I__1215\ : CascadeMux
    port map (
            O => \N__7430\,
            I => \rFifoDatarff_0_RNIHJV05_cascade_\
        );

    \I__1214\ : InMux
    port map (
            O => \N__7427\,
            I => \N__7423\
        );

    \I__1213\ : InMux
    port map (
            O => \N__7426\,
            I => \N__7419\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__7423\,
            I => \N__7415\
        );

    \I__1211\ : InMux
    port map (
            O => \N__7422\,
            I => \N__7412\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__7419\,
            I => \N__7409\
        );

    \I__1209\ : InMux
    port map (
            O => \N__7418\,
            I => \N__7406\
        );

    \I__1208\ : Span4Mux_v
    port map (
            O => \N__7415\,
            I => \N__7401\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__7412\,
            I => \N__7401\
        );

    \I__1206\ : Span4Mux_v
    port map (
            O => \N__7409\,
            I => \N__7396\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__7406\,
            I => \N__7396\
        );

    \I__1204\ : Span4Mux_v
    port map (
            O => \N__7401\,
            I => \N__7393\
        );

    \I__1203\ : Span4Mux_h
    port map (
            O => \N__7396\,
            I => \N__7390\
        );

    \I__1202\ : Odrv4
    port map (
            O => \N__7393\,
            I => \DUT.wRxByte_0\
        );

    \I__1201\ : Odrv4
    port map (
            O => \N__7390\,
            I => \DUT.wRxByte_0\
        );

    \I__1200\ : InMux
    port map (
            O => \N__7385\,
            I => \N__7382\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__7382\,
            I => \N__7379\
        );

    \I__1198\ : Odrv4
    port map (
            O => \N__7379\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_0\
        );

    \I__1197\ : InMux
    port map (
            O => \N__7376\,
            I => \N__7371\
        );

    \I__1196\ : InMux
    port map (
            O => \N__7375\,
            I => \N__7367\
        );

    \I__1195\ : InMux
    port map (
            O => \N__7374\,
            I => \N__7364\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__7371\,
            I => \N__7361\
        );

    \I__1193\ : InMux
    port map (
            O => \N__7370\,
            I => \N__7358\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__7367\,
            I => \N__7355\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__7364\,
            I => \N__7352\
        );

    \I__1190\ : Span4Mux_v
    port map (
            O => \N__7361\,
            I => \N__7348\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__7358\,
            I => \N__7345\
        );

    \I__1188\ : Span4Mux_v
    port map (
            O => \N__7355\,
            I => \N__7340\
        );

    \I__1187\ : Span4Mux_h
    port map (
            O => \N__7352\,
            I => \N__7340\
        );

    \I__1186\ : InMux
    port map (
            O => \N__7351\,
            I => \N__7337\
        );

    \I__1185\ : Odrv4
    port map (
            O => \N__7348\,
            I => \DUT.wRxByte_1\
        );

    \I__1184\ : Odrv12
    port map (
            O => \N__7345\,
            I => \DUT.wRxByte_1\
        );

    \I__1183\ : Odrv4
    port map (
            O => \N__7340\,
            I => \DUT.wRxByte_1\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__7337\,
            I => \DUT.wRxByte_1\
        );

    \I__1181\ : InMux
    port map (
            O => \N__7328\,
            I => \N__7323\
        );

    \I__1180\ : InMux
    port map (
            O => \N__7327\,
            I => \N__7320\
        );

    \I__1179\ : InMux
    port map (
            O => \N__7326\,
            I => \N__7316\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__7323\,
            I => \N__7313\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__7320\,
            I => \N__7310\
        );

    \I__1176\ : InMux
    port map (
            O => \N__7319\,
            I => \N__7307\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__7316\,
            I => \N__7304\
        );

    \I__1174\ : Span4Mux_v
    port map (
            O => \N__7313\,
            I => \N__7298\
        );

    \I__1173\ : Span4Mux_h
    port map (
            O => \N__7310\,
            I => \N__7298\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__7307\,
            I => \N__7295\
        );

    \I__1171\ : Span4Mux_h
    port map (
            O => \N__7304\,
            I => \N__7292\
        );

    \I__1170\ : InMux
    port map (
            O => \N__7303\,
            I => \N__7289\
        );

    \I__1169\ : Odrv4
    port map (
            O => \N__7298\,
            I => \DUT.wRxByte_2\
        );

    \I__1168\ : Odrv12
    port map (
            O => \N__7295\,
            I => \DUT.wRxByte_2\
        );

    \I__1167\ : Odrv4
    port map (
            O => \N__7292\,
            I => \DUT.wRxByte_2\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__7289\,
            I => \DUT.wRxByte_2\
        );

    \I__1165\ : InMux
    port map (
            O => \N__7280\,
            I => \N__7277\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__7277\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_2\
        );

    \I__1163\ : InMux
    port map (
            O => \N__7274\,
            I => \N__7268\
        );

    \I__1162\ : InMux
    port map (
            O => \N__7273\,
            I => \N__7259\
        );

    \I__1161\ : InMux
    port map (
            O => \N__7272\,
            I => \N__7259\
        );

    \I__1160\ : InMux
    port map (
            O => \N__7271\,
            I => \N__7256\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__7268\,
            I => \N__7253\
        );

    \I__1158\ : InMux
    port map (
            O => \N__7267\,
            I => \N__7244\
        );

    \I__1157\ : InMux
    port map (
            O => \N__7266\,
            I => \N__7244\
        );

    \I__1156\ : InMux
    port map (
            O => \N__7265\,
            I => \N__7244\
        );

    \I__1155\ : InMux
    port map (
            O => \N__7264\,
            I => \N__7244\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__7259\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__7256\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__7253\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__7244\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\
        );

    \I__1150\ : CascadeMux
    port map (
            O => \N__7235\,
            I => \N__7230\
        );

    \I__1149\ : InMux
    port map (
            O => \N__7234\,
            I => \N__7225\
        );

    \I__1148\ : InMux
    port map (
            O => \N__7233\,
            I => \N__7222\
        );

    \I__1147\ : InMux
    port map (
            O => \N__7230\,
            I => \N__7217\
        );

    \I__1146\ : InMux
    port map (
            O => \N__7229\,
            I => \N__7217\
        );

    \I__1145\ : InMux
    port map (
            O => \N__7228\,
            I => \N__7214\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__7225\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_1\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__7222\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_1\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__7217\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_1\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__7214\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_1\
        );

    \I__1140\ : CEMux
    port map (
            O => \N__7205\,
            I => \N__7202\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__7202\,
            I => \N__7199\
        );

    \I__1138\ : Span4Mux_h
    port map (
            O => \N__7199\,
            I => \N__7196\
        );

    \I__1137\ : Odrv4
    port map (
            O => \N__7196\,
            I => \DUT.fifo_tx_inst.rFifoData_awe2\
        );

    \I__1136\ : CascadeMux
    port map (
            O => \N__7193\,
            I => \DUT.fifo_tx_inst.rFifoData_awe2_cascade_\
        );

    \I__1135\ : InMux
    port map (
            O => \N__7190\,
            I => \N__7184\
        );

    \I__1134\ : InMux
    port map (
            O => \N__7189\,
            I => \N__7184\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__7184\,
            I => \DUT.fifo_tx_inst.rFifoDataro_3\
        );

    \I__1132\ : InMux
    port map (
            O => \N__7181\,
            I => \N__7175\
        );

    \I__1131\ : InMux
    port map (
            O => \N__7180\,
            I => \N__7175\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__7175\,
            I => \DUT.fifo_tx_inst.rFifoDataro_2\
        );

    \I__1129\ : CascadeMux
    port map (
            O => \N__7172\,
            I => \DUT.fifo_tx_inst.rFifoData_awe0_cascade_\
        );

    \I__1128\ : InMux
    port map (
            O => \N__7169\,
            I => \N__7163\
        );

    \I__1127\ : InMux
    port map (
            O => \N__7168\,
            I => \N__7163\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__7163\,
            I => \DUT.fifo_rx_inst.rFifoDataro_0\
        );

    \I__1125\ : CEMux
    port map (
            O => \N__7160\,
            I => \N__7157\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__7157\,
            I => \N__7154\
        );

    \I__1123\ : Odrv12
    port map (
            O => \N__7154\,
            I => \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa\
        );

    \I__1122\ : CascadeMux
    port map (
            O => \N__7151\,
            I => \DUT.fifo_rx_inst.N_87_cascade_\
        );

    \I__1121\ : InMux
    port map (
            O => \N__7148\,
            I => \N__7145\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__7145\,
            I => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0\
        );

    \I__1119\ : InMux
    port map (
            O => \N__7142\,
            I => \N__7135\
        );

    \I__1118\ : CascadeMux
    port map (
            O => \N__7141\,
            I => \N__7132\
        );

    \I__1117\ : InMux
    port map (
            O => \N__7140\,
            I => \N__7127\
        );

    \I__1116\ : InMux
    port map (
            O => \N__7139\,
            I => \N__7122\
        );

    \I__1115\ : InMux
    port map (
            O => \N__7138\,
            I => \N__7122\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__7135\,
            I => \N__7119\
        );

    \I__1113\ : InMux
    port map (
            O => \N__7132\,
            I => \N__7112\
        );

    \I__1112\ : InMux
    port map (
            O => \N__7131\,
            I => \N__7112\
        );

    \I__1111\ : InMux
    port map (
            O => \N__7130\,
            I => \N__7112\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__7127\,
            I => \N__7107\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__7122\,
            I => \N__7107\
        );

    \I__1108\ : Span4Mux_v
    port map (
            O => \N__7119\,
            I => \N__7099\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__7112\,
            I => \N__7099\
        );

    \I__1106\ : Span4Mux_h
    port map (
            O => \N__7107\,
            I => \N__7099\
        );

    \I__1105\ : InMux
    port map (
            O => \N__7106\,
            I => \N__7096\
        );

    \I__1104\ : Sp12to4
    port map (
            O => \N__7099\,
            I => \N__7091\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__7096\,
            I => \N__7091\
        );

    \I__1102\ : Odrv12
    port map (
            O => \N__7091\,
            I => \DUT.wRcvd\
        );

    \I__1101\ : CascadeMux
    port map (
            O => \N__7088\,
            I => \N__7085\
        );

    \I__1100\ : InMux
    port map (
            O => \N__7085\,
            I => \N__7082\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__7082\,
            I => \DUT.fifo_rx_inst.N_87\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__7079\,
            I => \DUT.fifo_rx_inst.N_92_cascade_\
        );

    \I__1097\ : CascadeMux
    port map (
            O => \N__7076\,
            I => \N__7073\
        );

    \I__1096\ : InMux
    port map (
            O => \N__7073\,
            I => \N__7065\
        );

    \I__1095\ : InMux
    port map (
            O => \N__7072\,
            I => \N__7062\
        );

    \I__1094\ : InMux
    port map (
            O => \N__7071\,
            I => \N__7053\
        );

    \I__1093\ : InMux
    port map (
            O => \N__7070\,
            I => \N__7053\
        );

    \I__1092\ : InMux
    port map (
            O => \N__7069\,
            I => \N__7053\
        );

    \I__1091\ : InMux
    port map (
            O => \N__7068\,
            I => \N__7053\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__7065\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_0\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__7062\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_0\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__7053\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_0\
        );

    \I__1087\ : CascadeMux
    port map (
            O => \N__7046\,
            I => \DUT.fifo_tx_inst.rFifoData_awe3_cascade_\
        );

    \I__1086\ : InMux
    port map (
            O => \N__7043\,
            I => \N__7040\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__7040\,
            I => \DUT.fifo_tx_inst.un1_i11_i\
        );

    \I__1084\ : CascadeMux
    port map (
            O => \N__7037\,
            I => \DUT.fifo_tx_inst.un1_i11_i_cascade_\
        );

    \I__1083\ : CascadeMux
    port map (
            O => \N__7034\,
            I => \N__7026\
        );

    \I__1082\ : CascadeMux
    port map (
            O => \N__7033\,
            I => \N__7023\
        );

    \I__1081\ : CascadeMux
    port map (
            O => \N__7032\,
            I => \N__7020\
        );

    \I__1080\ : InMux
    port map (
            O => \N__7031\,
            I => \N__7013\
        );

    \I__1079\ : InMux
    port map (
            O => \N__7030\,
            I => \N__7013\
        );

    \I__1078\ : InMux
    port map (
            O => \N__7029\,
            I => \N__7010\
        );

    \I__1077\ : InMux
    port map (
            O => \N__7026\,
            I => \N__7003\
        );

    \I__1076\ : InMux
    port map (
            O => \N__7023\,
            I => \N__7003\
        );

    \I__1075\ : InMux
    port map (
            O => \N__7020\,
            I => \N__7003\
        );

    \I__1074\ : CascadeMux
    port map (
            O => \N__7019\,
            I => \N__6999\
        );

    \I__1073\ : CascadeMux
    port map (
            O => \N__7018\,
            I => \N__6995\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__7013\,
            I => \N__6986\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__7010\,
            I => \N__6986\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__7003\,
            I => \N__6986\
        );

    \I__1069\ : InMux
    port map (
            O => \N__7002\,
            I => \N__6981\
        );

    \I__1068\ : InMux
    port map (
            O => \N__6999\,
            I => \N__6981\
        );

    \I__1067\ : InMux
    port map (
            O => \N__6998\,
            I => \N__6974\
        );

    \I__1066\ : InMux
    port map (
            O => \N__6995\,
            I => \N__6974\
        );

    \I__1065\ : InMux
    port map (
            O => \N__6994\,
            I => \N__6974\
        );

    \I__1064\ : InMux
    port map (
            O => \N__6993\,
            I => \N__6971\
        );

    \I__1063\ : Span4Mux_v
    port map (
            O => \N__6986\,
            I => \N__6966\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__6981\,
            I => \N__6966\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__6974\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_4\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__6971\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_4\
        );

    \I__1059\ : Odrv4
    port map (
            O => \N__6966\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_4\
        );

    \I__1058\ : CascadeMux
    port map (
            O => \N__6959\,
            I => \N__6956\
        );

    \I__1057\ : InMux
    port map (
            O => \N__6956\,
            I => \N__6948\
        );

    \I__1056\ : InMux
    port map (
            O => \N__6955\,
            I => \N__6948\
        );

    \I__1055\ : InMux
    port map (
            O => \N__6954\,
            I => \N__6942\
        );

    \I__1054\ : InMux
    port map (
            O => \N__6953\,
            I => \N__6942\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__6948\,
            I => \N__6932\
        );

    \I__1052\ : CascadeMux
    port map (
            O => \N__6947\,
            I => \N__6929\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__6942\,
            I => \N__6926\
        );

    \I__1050\ : InMux
    port map (
            O => \N__6941\,
            I => \N__6923\
        );

    \I__1049\ : InMux
    port map (
            O => \N__6940\,
            I => \N__6918\
        );

    \I__1048\ : InMux
    port map (
            O => \N__6939\,
            I => \N__6918\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6938\,
            I => \N__6909\
        );

    \I__1046\ : InMux
    port map (
            O => \N__6937\,
            I => \N__6909\
        );

    \I__1045\ : InMux
    port map (
            O => \N__6936\,
            I => \N__6909\
        );

    \I__1044\ : InMux
    port map (
            O => \N__6935\,
            I => \N__6909\
        );

    \I__1043\ : Span4Mux_h
    port map (
            O => \N__6932\,
            I => \N__6906\
        );

    \I__1042\ : InMux
    port map (
            O => \N__6929\,
            I => \N__6903\
        );

    \I__1041\ : Odrv4
    port map (
            O => \N__6926\,
            I => \DUT.uart_inst0.rx_countdownZ1Z_3\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__6923\,
            I => \DUT.uart_inst0.rx_countdownZ1Z_3\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__6918\,
            I => \DUT.uart_inst0.rx_countdownZ1Z_3\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__6909\,
            I => \DUT.uart_inst0.rx_countdownZ1Z_3\
        );

    \I__1037\ : Odrv4
    port map (
            O => \N__6906\,
            I => \DUT.uart_inst0.rx_countdownZ1Z_3\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__6903\,
            I => \DUT.uart_inst0.rx_countdownZ1Z_3\
        );

    \I__1035\ : CascadeMux
    port map (
            O => \N__6890\,
            I => \N__6886\
        );

    \I__1034\ : CascadeMux
    port map (
            O => \N__6889\,
            I => \N__6883\
        );

    \I__1033\ : InMux
    port map (
            O => \N__6886\,
            I => \N__6880\
        );

    \I__1032\ : InMux
    port map (
            O => \N__6883\,
            I => \N__6877\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__6880\,
            I => \DUT.uart_inst0.N_13_mux\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__6877\,
            I => \DUT.uart_inst0.N_13_mux\
        );

    \I__1029\ : InMux
    port map (
            O => \N__6872\,
            I => \N__6864\
        );

    \I__1028\ : InMux
    port map (
            O => \N__6871\,
            I => \N__6864\
        );

    \I__1027\ : InMux
    port map (
            O => \N__6870\,
            I => \N__6859\
        );

    \I__1026\ : CascadeMux
    port map (
            O => \N__6869\,
            I => \N__6855\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__6864\,
            I => \N__6848\
        );

    \I__1024\ : InMux
    port map (
            O => \N__6863\,
            I => \N__6843\
        );

    \I__1023\ : InMux
    port map (
            O => \N__6862\,
            I => \N__6843\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__6859\,
            I => \N__6840\
        );

    \I__1021\ : InMux
    port map (
            O => \N__6858\,
            I => \N__6837\
        );

    \I__1020\ : InMux
    port map (
            O => \N__6855\,
            I => \N__6834\
        );

    \I__1019\ : InMux
    port map (
            O => \N__6854\,
            I => \N__6831\
        );

    \I__1018\ : InMux
    port map (
            O => \N__6853\,
            I => \N__6828\
        );

    \I__1017\ : InMux
    port map (
            O => \N__6852\,
            I => \N__6823\
        );

    \I__1016\ : InMux
    port map (
            O => \N__6851\,
            I => \N__6823\
        );

    \I__1015\ : Span4Mux_h
    port map (
            O => \N__6848\,
            I => \N__6818\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__6843\,
            I => \N__6818\
        );

    \I__1013\ : Span4Mux_v
    port map (
            O => \N__6840\,
            I => \N__6813\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__6837\,
            I => \N__6813\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__6834\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_2\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__6831\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_2\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__6828\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_2\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__6823\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_2\
        );

    \I__1007\ : Odrv4
    port map (
            O => \N__6818\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_2\
        );

    \I__1006\ : Odrv4
    port map (
            O => \N__6813\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_2\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6800\,
            I => \N__6797\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__6797\,
            I => \N__6785\
        );

    \I__1003\ : CascadeMux
    port map (
            O => \N__6796\,
            I => \N__6782\
        );

    \I__1002\ : InMux
    port map (
            O => \N__6795\,
            I => \N__6777\
        );

    \I__1001\ : InMux
    port map (
            O => \N__6794\,
            I => \N__6768\
        );

    \I__1000\ : InMux
    port map (
            O => \N__6793\,
            I => \N__6768\
        );

    \I__999\ : InMux
    port map (
            O => \N__6792\,
            I => \N__6768\
        );

    \I__998\ : InMux
    port map (
            O => \N__6791\,
            I => \N__6768\
        );

    \I__997\ : InMux
    port map (
            O => \N__6790\,
            I => \N__6765\
        );

    \I__996\ : InMux
    port map (
            O => \N__6789\,
            I => \N__6760\
        );

    \I__995\ : InMux
    port map (
            O => \N__6788\,
            I => \N__6760\
        );

    \I__994\ : Span4Mux_h
    port map (
            O => \N__6785\,
            I => \N__6757\
        );

    \I__993\ : InMux
    port map (
            O => \N__6782\,
            I => \N__6754\
        );

    \I__992\ : InMux
    port map (
            O => \N__6781\,
            I => \N__6749\
        );

    \I__991\ : InMux
    port map (
            O => \N__6780\,
            I => \N__6749\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__6777\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_5\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__6768\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_5\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__6765\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_5\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__6760\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_5\
        );

    \I__986\ : Odrv4
    port map (
            O => \N__6757\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_5\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__6754\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_5\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__6749\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_5\
        );

    \I__983\ : InMux
    port map (
            O => \N__6734\,
            I => \N__6726\
        );

    \I__982\ : CascadeMux
    port map (
            O => \N__6733\,
            I => \N__6723\
        );

    \I__981\ : CascadeMux
    port map (
            O => \N__6732\,
            I => \N__6720\
        );

    \I__980\ : InMux
    port map (
            O => \N__6731\,
            I => \N__6714\
        );

    \I__979\ : InMux
    port map (
            O => \N__6730\,
            I => \N__6714\
        );

    \I__978\ : CascadeMux
    port map (
            O => \N__6729\,
            I => \N__6708\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__6726\,
            I => \N__6705\
        );

    \I__976\ : InMux
    port map (
            O => \N__6723\,
            I => \N__6700\
        );

    \I__975\ : InMux
    port map (
            O => \N__6720\,
            I => \N__6700\
        );

    \I__974\ : InMux
    port map (
            O => \N__6719\,
            I => \N__6692\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__6714\,
            I => \N__6689\
        );

    \I__972\ : InMux
    port map (
            O => \N__6713\,
            I => \N__6680\
        );

    \I__971\ : InMux
    port map (
            O => \N__6712\,
            I => \N__6680\
        );

    \I__970\ : CascadeMux
    port map (
            O => \N__6711\,
            I => \N__6675\
        );

    \I__969\ : InMux
    port map (
            O => \N__6708\,
            I => \N__6672\
        );

    \I__968\ : Span4Mux_h
    port map (
            O => \N__6705\,
            I => \N__6669\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__6700\,
            I => \N__6666\
        );

    \I__966\ : InMux
    port map (
            O => \N__6699\,
            I => \N__6659\
        );

    \I__965\ : InMux
    port map (
            O => \N__6698\,
            I => \N__6659\
        );

    \I__964\ : InMux
    port map (
            O => \N__6697\,
            I => \N__6659\
        );

    \I__963\ : InMux
    port map (
            O => \N__6696\,
            I => \N__6654\
        );

    \I__962\ : InMux
    port map (
            O => \N__6695\,
            I => \N__6654\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__6692\,
            I => \N__6649\
        );

    \I__960\ : Span4Mux_h
    port map (
            O => \N__6689\,
            I => \N__6649\
        );

    \I__959\ : InMux
    port map (
            O => \N__6688\,
            I => \N__6644\
        );

    \I__958\ : InMux
    port map (
            O => \N__6687\,
            I => \N__6644\
        );

    \I__957\ : InMux
    port map (
            O => \N__6686\,
            I => \N__6639\
        );

    \I__956\ : InMux
    port map (
            O => \N__6685\,
            I => \N__6639\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__6680\,
            I => \N__6636\
        );

    \I__954\ : InMux
    port map (
            O => \N__6679\,
            I => \N__6631\
        );

    \I__953\ : InMux
    port map (
            O => \N__6678\,
            I => \N__6631\
        );

    \I__952\ : InMux
    port map (
            O => \N__6675\,
            I => \N__6628\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__6672\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__950\ : Odrv4
    port map (
            O => \N__6669\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__949\ : Odrv4
    port map (
            O => \N__6666\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__6659\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__6654\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__946\ : Odrv4
    port map (
            O => \N__6649\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__6644\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__6639\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__943\ : Odrv4
    port map (
            O => \N__6636\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__6631\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__6628\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__940\ : CascadeMux
    port map (
            O => \N__6605\,
            I => \DUT.uart_inst0.N_8_0_cascade_\
        );

    \I__939\ : InMux
    port map (
            O => \N__6602\,
            I => \N__6599\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__6599\,
            I => \DUT.uart_inst0.m10_0_1\
        );

    \I__937\ : InMux
    port map (
            O => \N__6596\,
            I => \N__6593\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__6593\,
            I => \N__6590\
        );

    \I__935\ : Odrv4
    port map (
            O => \N__6590\,
            I => \DUT.uart_inst0.m11_0\
        );

    \I__934\ : InMux
    port map (
            O => \N__6587\,
            I => \N__6584\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__6584\,
            I => \N__6581\
        );

    \I__932\ : Odrv4
    port map (
            O => \N__6581\,
            I => \DUT.uart_inst0.N_15_mux\
        );

    \I__931\ : CascadeMux
    port map (
            O => \N__6578\,
            I => \DUT.uart_inst0.N_11_0_cascade_\
        );

    \I__930\ : CascadeMux
    port map (
            O => \N__6575\,
            I => \N__6572\
        );

    \I__929\ : InMux
    port map (
            O => \N__6572\,
            I => \N__6569\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__6569\,
            I => \DUT.uart_inst0.N_81_mux_i_i_a5_1_3\
        );

    \I__927\ : CascadeMux
    port map (
            O => \N__6566\,
            I => \N__6555\
        );

    \I__926\ : InMux
    port map (
            O => \N__6565\,
            I => \N__6550\
        );

    \I__925\ : InMux
    port map (
            O => \N__6564\,
            I => \N__6547\
        );

    \I__924\ : InMux
    port map (
            O => \N__6563\,
            I => \N__6542\
        );

    \I__923\ : InMux
    port map (
            O => \N__6562\,
            I => \N__6542\
        );

    \I__922\ : InMux
    port map (
            O => \N__6561\,
            I => \N__6537\
        );

    \I__921\ : InMux
    port map (
            O => \N__6560\,
            I => \N__6537\
        );

    \I__920\ : InMux
    port map (
            O => \N__6559\,
            I => \N__6532\
        );

    \I__919\ : InMux
    port map (
            O => \N__6558\,
            I => \N__6532\
        );

    \I__918\ : InMux
    port map (
            O => \N__6555\,
            I => \N__6525\
        );

    \I__917\ : InMux
    port map (
            O => \N__6554\,
            I => \N__6525\
        );

    \I__916\ : InMux
    port map (
            O => \N__6553\,
            I => \N__6525\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__6550\,
            I => \N__6522\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__6547\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_3\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__6542\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_3\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__6537\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_3\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__6532\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_3\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__6525\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_3\
        );

    \I__909\ : Odrv4
    port map (
            O => \N__6522\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_3\
        );

    \I__908\ : CascadeMux
    port map (
            O => \N__6509\,
            I => \DUT.uart_inst0.N_300_cascade_\
        );

    \I__907\ : CascadeMux
    port map (
            O => \N__6506\,
            I => \DUT.uart_inst0.G_16_i_a3_3_cascade_\
        );

    \I__906\ : InMux
    port map (
            O => \N__6503\,
            I => \N__6500\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__6500\,
            I => \N__6497\
        );

    \I__904\ : Odrv12
    port map (
            O => \N__6497\,
            I => \DUT.uart_inst0.G_16_i_a3_4\
        );

    \I__903\ : InMux
    port map (
            O => \N__6494\,
            I => \N__6488\
        );

    \I__902\ : InMux
    port map (
            O => \N__6493\,
            I => \N__6484\
        );

    \I__901\ : CascadeMux
    port map (
            O => \N__6492\,
            I => \N__6474\
        );

    \I__900\ : InMux
    port map (
            O => \N__6491\,
            I => \N__6471\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__6488\,
            I => \N__6468\
        );

    \I__898\ : InMux
    port map (
            O => \N__6487\,
            I => \N__6465\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__6484\,
            I => \N__6462\
        );

    \I__896\ : InMux
    port map (
            O => \N__6483\,
            I => \N__6455\
        );

    \I__895\ : InMux
    port map (
            O => \N__6482\,
            I => \N__6455\
        );

    \I__894\ : InMux
    port map (
            O => \N__6481\,
            I => \N__6455\
        );

    \I__893\ : InMux
    port map (
            O => \N__6480\,
            I => \N__6446\
        );

    \I__892\ : InMux
    port map (
            O => \N__6479\,
            I => \N__6446\
        );

    \I__891\ : InMux
    port map (
            O => \N__6478\,
            I => \N__6446\
        );

    \I__890\ : InMux
    port map (
            O => \N__6477\,
            I => \N__6446\
        );

    \I__889\ : InMux
    port map (
            O => \N__6474\,
            I => \N__6443\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__6471\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_1\
        );

    \I__887\ : Odrv4
    port map (
            O => \N__6468\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_1\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__6465\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_1\
        );

    \I__885\ : Odrv4
    port map (
            O => \N__6462\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_1\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__6455\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_1\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__6446\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_1\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__6443\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_1\
        );

    \I__881\ : InMux
    port map (
            O => \N__6428\,
            I => \N__6421\
        );

    \I__880\ : InMux
    port map (
            O => \N__6427\,
            I => \N__6416\
        );

    \I__879\ : CascadeMux
    port map (
            O => \N__6426\,
            I => \N__6413\
        );

    \I__878\ : InMux
    port map (
            O => \N__6425\,
            I => \N__6409\
        );

    \I__877\ : CascadeMux
    port map (
            O => \N__6424\,
            I => \N__6406\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__6421\,
            I => \N__6401\
        );

    \I__875\ : CascadeMux
    port map (
            O => \N__6420\,
            I => \N__6397\
        );

    \I__874\ : InMux
    port map (
            O => \N__6419\,
            I => \N__6393\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__6416\,
            I => \N__6390\
        );

    \I__872\ : InMux
    port map (
            O => \N__6413\,
            I => \N__6385\
        );

    \I__871\ : InMux
    port map (
            O => \N__6412\,
            I => \N__6385\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__6409\,
            I => \N__6382\
        );

    \I__869\ : InMux
    port map (
            O => \N__6406\,
            I => \N__6379\
        );

    \I__868\ : InMux
    port map (
            O => \N__6405\,
            I => \N__6374\
        );

    \I__867\ : InMux
    port map (
            O => \N__6404\,
            I => \N__6374\
        );

    \I__866\ : Span4Mux_h
    port map (
            O => \N__6401\,
            I => \N__6371\
        );

    \I__865\ : InMux
    port map (
            O => \N__6400\,
            I => \N__6368\
        );

    \I__864\ : InMux
    port map (
            O => \N__6397\,
            I => \N__6363\
        );

    \I__863\ : InMux
    port map (
            O => \N__6396\,
            I => \N__6363\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__6393\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_5\
        );

    \I__861\ : Odrv4
    port map (
            O => \N__6390\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_5\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__6385\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_5\
        );

    \I__859\ : Odrv4
    port map (
            O => \N__6382\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_5\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__6379\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_5\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__6374\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_5\
        );

    \I__856\ : Odrv4
    port map (
            O => \N__6371\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_5\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__6368\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_5\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__6363\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_5\
        );

    \I__853\ : InMux
    port map (
            O => \N__6344\,
            I => \N__6341\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__6341\,
            I => \N__6338\
        );

    \I__851\ : Odrv12
    port map (
            O => \N__6338\,
            I => \DUT.uart_inst0.N_11_2\
        );

    \I__850\ : CascadeMux
    port map (
            O => \N__6335\,
            I => \N__6329\
        );

    \I__849\ : InMux
    port map (
            O => \N__6334\,
            I => \N__6326\
        );

    \I__848\ : CascadeMux
    port map (
            O => \N__6333\,
            I => \N__6322\
        );

    \I__847\ : CascadeMux
    port map (
            O => \N__6332\,
            I => \N__6317\
        );

    \I__846\ : InMux
    port map (
            O => \N__6329\,
            I => \N__6311\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__6326\,
            I => \N__6308\
        );

    \I__844\ : InMux
    port map (
            O => \N__6325\,
            I => \N__6305\
        );

    \I__843\ : InMux
    port map (
            O => \N__6322\,
            I => \N__6302\
        );

    \I__842\ : InMux
    port map (
            O => \N__6321\,
            I => \N__6297\
        );

    \I__841\ : InMux
    port map (
            O => \N__6320\,
            I => \N__6297\
        );

    \I__840\ : InMux
    port map (
            O => \N__6317\,
            I => \N__6294\
        );

    \I__839\ : InMux
    port map (
            O => \N__6316\,
            I => \N__6287\
        );

    \I__838\ : InMux
    port map (
            O => \N__6315\,
            I => \N__6287\
        );

    \I__837\ : InMux
    port map (
            O => \N__6314\,
            I => \N__6287\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__6311\,
            I => \N__6284\
        );

    \I__835\ : Odrv4
    port map (
            O => \N__6308\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_2\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__6305\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_2\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__6302\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_2\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__6297\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_2\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__6294\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_2\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__6287\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_2\
        );

    \I__829\ : Odrv4
    port map (
            O => \N__6284\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_2\
        );

    \I__828\ : InMux
    port map (
            O => \N__6269\,
            I => \N__6266\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__6266\,
            I => \DUT.uart_inst0.G_16_i_a3_0_3\
        );

    \I__826\ : CascadeMux
    port map (
            O => \N__6263\,
            I => \N__6260\
        );

    \I__825\ : InMux
    port map (
            O => \N__6260\,
            I => \N__6257\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__6257\,
            I => \DUT.uart_inst0.g1_1\
        );

    \I__823\ : CascadeMux
    port map (
            O => \N__6254\,
            I => \N__6245\
        );

    \I__822\ : CascadeMux
    port map (
            O => \N__6253\,
            I => \N__6239\
        );

    \I__821\ : CascadeMux
    port map (
            O => \N__6252\,
            I => \N__6235\
        );

    \I__820\ : InMux
    port map (
            O => \N__6251\,
            I => \N__6231\
        );

    \I__819\ : InMux
    port map (
            O => \N__6250\,
            I => \N__6228\
        );

    \I__818\ : InMux
    port map (
            O => \N__6249\,
            I => \N__6225\
        );

    \I__817\ : InMux
    port map (
            O => \N__6248\,
            I => \N__6220\
        );

    \I__816\ : InMux
    port map (
            O => \N__6245\,
            I => \N__6220\
        );

    \I__815\ : InMux
    port map (
            O => \N__6244\,
            I => \N__6213\
        );

    \I__814\ : InMux
    port map (
            O => \N__6243\,
            I => \N__6213\
        );

    \I__813\ : InMux
    port map (
            O => \N__6242\,
            I => \N__6213\
        );

    \I__812\ : InMux
    port map (
            O => \N__6239\,
            I => \N__6208\
        );

    \I__811\ : InMux
    port map (
            O => \N__6238\,
            I => \N__6208\
        );

    \I__810\ : InMux
    port map (
            O => \N__6235\,
            I => \N__6205\
        );

    \I__809\ : InMux
    port map (
            O => \N__6234\,
            I => \N__6202\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__6231\,
            I => \N__6197\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__6228\,
            I => \N__6197\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__6225\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_1\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__6220\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_1\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__6213\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_1\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__6208\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_1\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__6205\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_1\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__6202\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_1\
        );

    \I__800\ : Odrv4
    port map (
            O => \N__6197\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_1\
        );

    \I__799\ : InMux
    port map (
            O => \N__6182\,
            I => \N__6179\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__6179\,
            I => \DUT.uart_inst0.N_81_mux_i_i_a5_1_5_0\
        );

    \I__797\ : InMux
    port map (
            O => \N__6176\,
            I => \N__6173\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__6173\,
            I => \DUT.uart_inst0.rx_countdown_RNO_2Z0Z_2\
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__6170\,
            I => \DUT.uart_inst0.G_21_0_1_0_cascade_\
        );

    \I__794\ : InMux
    port map (
            O => \N__6167\,
            I => \N__6164\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__6164\,
            I => \DUT.uart_inst0.G_9_i_o4_0\
        );

    \I__792\ : InMux
    port map (
            O => \N__6161\,
            I => \N__6158\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__6158\,
            I => \DUT.uart_inst0.g0_0_3\
        );

    \I__790\ : CascadeMux
    port map (
            O => \N__6155\,
            I => \DUT.uart_inst0.G_16_i_a3_0_2_cascade_\
        );

    \I__789\ : CascadeMux
    port map (
            O => \N__6152\,
            I => \DUT.uart_inst0.N_45_cascade_\
        );

    \I__788\ : InMux
    port map (
            O => \N__6149\,
            I => \N__6146\
        );

    \I__787\ : LocalMux
    port map (
            O => \N__6146\,
            I => \DUT.uart_inst0.N_55\
        );

    \I__786\ : InMux
    port map (
            O => \N__6143\,
            I => \N__6137\
        );

    \I__785\ : CascadeMux
    port map (
            O => \N__6142\,
            I => \N__6133\
        );

    \I__784\ : CascadeMux
    port map (
            O => \N__6141\,
            I => \N__6127\
        );

    \I__783\ : InMux
    port map (
            O => \N__6140\,
            I => \N__6121\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__6137\,
            I => \N__6118\
        );

    \I__781\ : InMux
    port map (
            O => \N__6136\,
            I => \N__6113\
        );

    \I__780\ : InMux
    port map (
            O => \N__6133\,
            I => \N__6113\
        );

    \I__779\ : InMux
    port map (
            O => \N__6132\,
            I => \N__6108\
        );

    \I__778\ : InMux
    port map (
            O => \N__6131\,
            I => \N__6108\
        );

    \I__777\ : InMux
    port map (
            O => \N__6130\,
            I => \N__6103\
        );

    \I__776\ : InMux
    port map (
            O => \N__6127\,
            I => \N__6103\
        );

    \I__775\ : InMux
    port map (
            O => \N__6126\,
            I => \N__6100\
        );

    \I__774\ : InMux
    port map (
            O => \N__6125\,
            I => \N__6095\
        );

    \I__773\ : InMux
    port map (
            O => \N__6124\,
            I => \N__6095\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__6121\,
            I => \N__6092\
        );

    \I__771\ : Odrv4
    port map (
            O => \N__6118\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_4\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__6113\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_4\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__6108\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_4\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__6103\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_4\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__6100\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_4\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__6095\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_4\
        );

    \I__765\ : Odrv4
    port map (
            O => \N__6092\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_4\
        );

    \I__764\ : InMux
    port map (
            O => \N__6077\,
            I => \N__6074\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__6074\,
            I => \DUT.uart_inst0.N_10\
        );

    \I__762\ : CascadeMux
    port map (
            O => \N__6071\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0_cascade_\
        );

    \I__761\ : InMux
    port map (
            O => \N__6068\,
            I => \N__6065\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__6065\,
            I => \DUT.uart_inst0.G_21_0_1\
        );

    \I__759\ : InMux
    port map (
            O => \N__6062\,
            I => \N__6059\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__6059\,
            I => \N__6055\
        );

    \I__757\ : InMux
    port map (
            O => \N__6058\,
            I => \N__6052\
        );

    \I__756\ : Odrv4
    port map (
            O => \N__6055\,
            I => \DUT.uart_inst0.recv_stateZ0Z_4\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__6052\,
            I => \DUT.uart_inst0.recv_stateZ0Z_4\
        );

    \I__754\ : CascadeMux
    port map (
            O => \N__6047\,
            I => \N__6043\
        );

    \I__753\ : InMux
    port map (
            O => \N__6046\,
            I => \N__6039\
        );

    \I__752\ : InMux
    port map (
            O => \N__6043\,
            I => \N__6034\
        );

    \I__751\ : InMux
    port map (
            O => \N__6042\,
            I => \N__6034\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__6039\,
            I => \DUT.uart_inst0.N_45\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__6034\,
            I => \DUT.uart_inst0.N_45\
        );

    \I__748\ : InMux
    port map (
            O => \N__6029\,
            I => \N__6026\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__6026\,
            I => \N__6023\
        );

    \I__746\ : Span4Mux_h
    port map (
            O => \N__6023\,
            I => \N__6020\
        );

    \I__745\ : Odrv4
    port map (
            O => \N__6020\,
            I => \DUT.uart_inst0.recv_state_ns_0_0_0\
        );

    \I__744\ : CascadeMux
    port map (
            O => \N__6017\,
            I => \N__6014\
        );

    \I__743\ : InMux
    port map (
            O => \N__6014\,
            I => \N__6011\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__6011\,
            I => \N__6008\
        );

    \I__741\ : Odrv4
    port map (
            O => \N__6008\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_2\
        );

    \I__740\ : InMux
    port map (
            O => \N__6005\,
            I => \N__6002\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__6002\,
            I => \N__5999\
        );

    \I__738\ : Odrv4
    port map (
            O => \N__5999\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_3\
        );

    \I__737\ : CascadeMux
    port map (
            O => \N__5996\,
            I => \N__5993\
        );

    \I__736\ : InMux
    port map (
            O => \N__5993\,
            I => \N__5990\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__5990\,
            I => \N__5987\
        );

    \I__734\ : Odrv4
    port map (
            O => \N__5987\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_4\
        );

    \I__733\ : CascadeMux
    port map (
            O => \N__5984\,
            I => \N__5981\
        );

    \I__732\ : InMux
    port map (
            O => \N__5981\,
            I => \N__5978\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__5978\,
            I => \N__5975\
        );

    \I__730\ : Odrv4
    port map (
            O => \N__5975\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_5\
        );

    \I__729\ : CascadeMux
    port map (
            O => \N__5972\,
            I => \N__5969\
        );

    \I__728\ : InMux
    port map (
            O => \N__5969\,
            I => \N__5966\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__5966\,
            I => \N__5963\
        );

    \I__726\ : Odrv4
    port map (
            O => \N__5963\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_6\
        );

    \I__725\ : InMux
    port map (
            O => \N__5960\,
            I => \N__5957\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__5957\,
            I => \DUT.uart_inst0.N_81_mux_i_i_a5_1_4\
        );

    \I__723\ : InMux
    port map (
            O => \N__5954\,
            I => \N__5951\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__5951\,
            I => \DUT.uart_inst0.N_13_0\
        );

    \I__721\ : InMux
    port map (
            O => \N__5948\,
            I => \N__5945\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__5945\,
            I => \N__5942\
        );

    \I__719\ : Odrv4
    port map (
            O => \N__5942\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_3\
        );

    \I__718\ : CascadeMux
    port map (
            O => \N__5939\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_\
        );

    \I__717\ : CascadeMux
    port map (
            O => \N__5936\,
            I => \N__5933\
        );

    \I__716\ : InMux
    port map (
            O => \N__5933\,
            I => \N__5930\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__5930\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_0\
        );

    \I__714\ : InMux
    port map (
            O => \N__5927\,
            I => \N__5924\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__5924\,
            I => \N__5921\
        );

    \I__712\ : Span4Mux_v
    port map (
            O => \N__5921\,
            I => \N__5918\
        );

    \I__711\ : Odrv4
    port map (
            O => \N__5918\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_0\
        );

    \I__710\ : CascadeMux
    port map (
            O => \N__5915\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_\
        );

    \I__709\ : InMux
    port map (
            O => \N__5912\,
            I => \N__5909\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__5909\,
            I => \N__5906\
        );

    \I__707\ : Span4Mux_h
    port map (
            O => \N__5906\,
            I => \N__5903\
        );

    \I__706\ : Odrv4
    port map (
            O => \N__5903\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_7\
        );

    \I__705\ : InMux
    port map (
            O => \N__5900\,
            I => \N__5897\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__5897\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_1\
        );

    \I__703\ : InMux
    port map (
            O => \N__5894\,
            I => \N__5891\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__5891\,
            I => \N__5888\
        );

    \I__701\ : Span4Mux_h
    port map (
            O => \N__5888\,
            I => \N__5885\
        );

    \I__700\ : Odrv4
    port map (
            O => \N__5885\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_2\
        );

    \I__699\ : InMux
    port map (
            O => \N__5882\,
            I => \N__5879\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__5879\,
            I => \N__5876\
        );

    \I__697\ : Odrv4
    port map (
            O => \N__5876\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2\
        );

    \I__696\ : InMux
    port map (
            O => \N__5873\,
            I => \N__5870\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__5870\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_0\
        );

    \I__694\ : CascadeMux
    port map (
            O => \N__5867\,
            I => \N__5864\
        );

    \I__693\ : InMux
    port map (
            O => \N__5864\,
            I => \N__5861\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__5861\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_1\
        );

    \I__691\ : InMux
    port map (
            O => \N__5858\,
            I => \N__5850\
        );

    \I__690\ : InMux
    port map (
            O => \N__5857\,
            I => \N__5850\
        );

    \I__689\ : InMux
    port map (
            O => \N__5856\,
            I => \N__5845\
        );

    \I__688\ : InMux
    port map (
            O => \N__5855\,
            I => \N__5845\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__5850\,
            I => \DUT.fifo_rx_inst.rWritePtr16\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__5845\,
            I => \DUT.fifo_rx_inst.rWritePtr16\
        );

    \I__685\ : CascadeMux
    port map (
            O => \N__5840\,
            I => \N__5836\
        );

    \I__684\ : InMux
    port map (
            O => \N__5839\,
            I => \N__5826\
        );

    \I__683\ : InMux
    port map (
            O => \N__5836\,
            I => \N__5826\
        );

    \I__682\ : InMux
    port map (
            O => \N__5835\,
            I => \N__5826\
        );

    \I__681\ : CascadeMux
    port map (
            O => \N__5834\,
            I => \N__5823\
        );

    \I__680\ : CascadeMux
    port map (
            O => \N__5833\,
            I => \N__5819\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__5826\,
            I => \N__5816\
        );

    \I__678\ : InMux
    port map (
            O => \N__5823\,
            I => \N__5809\
        );

    \I__677\ : InMux
    port map (
            O => \N__5822\,
            I => \N__5809\
        );

    \I__676\ : InMux
    port map (
            O => \N__5819\,
            I => \N__5809\
        );

    \I__675\ : Odrv4
    port map (
            O => \N__5816\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_0\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__5809\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_0\
        );

    \I__673\ : InMux
    port map (
            O => \N__5804\,
            I => \N__5793\
        );

    \I__672\ : InMux
    port map (
            O => \N__5803\,
            I => \N__5793\
        );

    \I__671\ : InMux
    port map (
            O => \N__5802\,
            I => \N__5793\
        );

    \I__670\ : InMux
    port map (
            O => \N__5801\,
            I => \N__5788\
        );

    \I__669\ : InMux
    port map (
            O => \N__5800\,
            I => \N__5788\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__5793\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_1\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__5788\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_1\
        );

    \I__666\ : InMux
    port map (
            O => \N__5783\,
            I => \N__5780\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__5780\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_2\
        );

    \I__664\ : CascadeMux
    port map (
            O => \N__5777\,
            I => \N__5774\
        );

    \I__663\ : InMux
    port map (
            O => \N__5774\,
            I => \N__5771\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__5771\,
            I => \N__5768\
        );

    \I__661\ : Odrv4
    port map (
            O => \N__5768\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_6\
        );

    \I__660\ : InMux
    port map (
            O => \N__5765\,
            I => \N__5762\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__5762\,
            I => \N__5759\
        );

    \I__658\ : Odrv4
    port map (
            O => \N__5759\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_4\
        );

    \I__657\ : InMux
    port map (
            O => \N__5756\,
            I => \N__5753\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__5753\,
            I => \N__5750\
        );

    \I__655\ : Odrv4
    port map (
            O => \N__5750\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_4\
        );

    \I__654\ : CascadeMux
    port map (
            O => \N__5747\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4_cascade_\
        );

    \I__653\ : InMux
    port map (
            O => \N__5744\,
            I => \N__5741\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__5741\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_5\
        );

    \I__651\ : CascadeMux
    port map (
            O => \N__5738\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_\
        );

    \I__650\ : InMux
    port map (
            O => \N__5735\,
            I => \N__5732\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__5732\,
            I => \N__5729\
        );

    \I__648\ : Odrv4
    port map (
            O => \N__5729\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_5\
        );

    \I__647\ : InMux
    port map (
            O => \N__5726\,
            I => \N__5723\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__5723\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_6\
        );

    \I__645\ : InMux
    port map (
            O => \N__5720\,
            I => \N__5717\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__5717\,
            I => \N__5714\
        );

    \I__643\ : Odrv4
    port map (
            O => \N__5714\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6\
        );

    \I__642\ : InMux
    port map (
            O => \N__5711\,
            I => \N__5708\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__5708\,
            I => \N__5705\
        );

    \I__640\ : Odrv4
    port map (
            O => \N__5705\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_3\
        );

    \I__639\ : CascadeMux
    port map (
            O => \N__5702\,
            I => \DUT.fifo_rx_inst.rFifoData_awe3_cascade_\
        );

    \I__638\ : CascadeMux
    port map (
            O => \N__5699\,
            I => \DUT.fifo_rx_inst.un1_i11_i_cascade_\
        );

    \I__637\ : InMux
    port map (
            O => \N__5696\,
            I => \N__5693\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__5693\,
            I => \DUT.fifo_rx_inst.un1_rFifoCount_1_axb_2\
        );

    \I__635\ : InMux
    port map (
            O => \N__5690\,
            I => \N__5687\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__5687\,
            I => \DUT.fifo_rx_inst.un1_i11_i\
        );

    \I__633\ : CascadeMux
    port map (
            O => \N__5684\,
            I => \N__5681\
        );

    \I__632\ : InMux
    port map (
            O => \N__5681\,
            I => \N__5678\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__5678\,
            I => \DUT.fifo_rx_inst.rFifoCount_RNIK3G92Z0Z_1\
        );

    \I__630\ : CascadeMux
    port map (
            O => \N__5675\,
            I => \DUT.fifo_rx_inst.rWritePtr16_cascade_\
        );

    \I__629\ : CascadeMux
    port map (
            O => \N__5672\,
            I => \DUT.uart_inst0.g0_0_i_a3_3_cascade_\
        );

    \I__628\ : InMux
    port map (
            O => \N__5669\,
            I => \N__5666\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__5666\,
            I => \DUT.uart_inst0.g0_0_i_a3_4\
        );

    \I__626\ : InMux
    port map (
            O => \N__5663\,
            I => \N__5660\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__5660\,
            I => \N__5654\
        );

    \I__624\ : InMux
    port map (
            O => \N__5659\,
            I => \N__5651\
        );

    \I__623\ : InMux
    port map (
            O => \N__5658\,
            I => \N__5646\
        );

    \I__622\ : InMux
    port map (
            O => \N__5657\,
            I => \N__5646\
        );

    \I__621\ : Span4Mux_h
    port map (
            O => \N__5654\,
            I => \N__5639\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__5651\,
            I => \N__5634\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__5646\,
            I => \N__5634\
        );

    \I__618\ : InMux
    port map (
            O => \N__5645\,
            I => \N__5629\
        );

    \I__617\ : InMux
    port map (
            O => \N__5644\,
            I => \N__5629\
        );

    \I__616\ : InMux
    port map (
            O => \N__5643\,
            I => \N__5626\
        );

    \I__615\ : InMux
    port map (
            O => \N__5642\,
            I => \N__5623\
        );

    \I__614\ : Odrv4
    port map (
            O => \N__5639\,
            I => \DUT.uart_inst0.recv_stateZ0Z_2\
        );

    \I__613\ : Odrv12
    port map (
            O => \N__5634\,
            I => \DUT.uart_inst0.recv_stateZ0Z_2\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__5629\,
            I => \DUT.uart_inst0.recv_stateZ0Z_2\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__5626\,
            I => \DUT.uart_inst0.recv_stateZ0Z_2\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__5623\,
            I => \DUT.uart_inst0.recv_stateZ0Z_2\
        );

    \I__609\ : IoInMux
    port map (
            O => \N__5612\,
            I => \N__5609\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__5609\,
            I => \N__5606\
        );

    \I__607\ : Span4Mux_s2_v
    port map (
            O => \N__5606\,
            I => \N__5603\
        );

    \I__606\ : Span4Mux_h
    port map (
            O => \N__5603\,
            I => \N__5600\
        );

    \I__605\ : Span4Mux_v
    port map (
            O => \N__5600\,
            I => \N__5597\
        );

    \I__604\ : Span4Mux_v
    port map (
            O => \N__5597\,
            I => \N__5594\
        );

    \I__603\ : Odrv4
    port map (
            O => \N__5594\,
            I => \wPllLocked_i\
        );

    \I__602\ : InMux
    port map (
            O => \N__5591\,
            I => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0\
        );

    \I__601\ : InMux
    port map (
            O => \N__5588\,
            I => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1\
        );

    \I__600\ : InMux
    port map (
            O => \N__5585\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_4_s1\
        );

    \I__599\ : InMux
    port map (
            O => \N__5582\,
            I => \N__5579\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__5579\,
            I => \DUT.uart_inst0.m9_3\
        );

    \I__597\ : InMux
    port map (
            O => \N__5576\,
            I => \N__5573\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__5573\,
            I => \DUT.uart_inst0.m9_4\
        );

    \I__595\ : InMux
    port map (
            O => \N__5570\,
            I => \N__5567\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__5567\,
            I => \DUT.uart_inst0.N_8\
        );

    \I__593\ : CascadeMux
    port map (
            O => \N__5564\,
            I => \N__5561\
        );

    \I__592\ : InMux
    port map (
            O => \N__5561\,
            I => \N__5558\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__5558\,
            I => \DUT.uart_inst0.N_81_mux_i_i_0_0\
        );

    \I__590\ : InMux
    port map (
            O => \N__5555\,
            I => \N__5552\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__5552\,
            I => \DUT.uart_inst0.N_81_mux_i_i_a5_0_5_0\
        );

    \I__588\ : CascadeMux
    port map (
            O => \N__5549\,
            I => \DUT.uart_inst0.m4_3_cascade_\
        );

    \I__587\ : CascadeMux
    port map (
            O => \N__5546\,
            I => \N__5543\
        );

    \I__586\ : InMux
    port map (
            O => \N__5543\,
            I => \N__5540\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__5540\,
            I => \DUT.uart_inst0.N_18_mux\
        );

    \I__584\ : CascadeMux
    port map (
            O => \N__5537\,
            I => \DUT.uart_inst0.N_297_cascade_\
        );

    \I__583\ : InMux
    port map (
            O => \N__5534\,
            I => \N__5523\
        );

    \I__582\ : InMux
    port map (
            O => \N__5533\,
            I => \N__5523\
        );

    \I__581\ : InMux
    port map (
            O => \N__5532\,
            I => \N__5517\
        );

    \I__580\ : InMux
    port map (
            O => \N__5531\,
            I => \N__5517\
        );

    \I__579\ : InMux
    port map (
            O => \N__5530\,
            I => \N__5512\
        );

    \I__578\ : InMux
    port map (
            O => \N__5529\,
            I => \N__5512\
        );

    \I__577\ : CascadeMux
    port map (
            O => \N__5528\,
            I => \N__5508\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__5523\,
            I => \N__5503\
        );

    \I__575\ : InMux
    port map (
            O => \N__5522\,
            I => \N__5500\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__5517\,
            I => \N__5495\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__5512\,
            I => \N__5495\
        );

    \I__572\ : InMux
    port map (
            O => \N__5511\,
            I => \N__5492\
        );

    \I__571\ : InMux
    port map (
            O => \N__5508\,
            I => \N__5489\
        );

    \I__570\ : InMux
    port map (
            O => \N__5507\,
            I => \N__5486\
        );

    \I__569\ : InMux
    port map (
            O => \N__5506\,
            I => \N__5483\
        );

    \I__568\ : Odrv4
    port map (
            O => \N__5503\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__5500\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__566\ : Odrv4
    port map (
            O => \N__5495\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__5492\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__5489\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__5486\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__5483\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__561\ : InMux
    port map (
            O => \N__5468\,
            I => \N__5465\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__5465\,
            I => \DUT.uart_inst0.N_15_3\
        );

    \I__559\ : InMux
    port map (
            O => \N__5462\,
            I => \N__5459\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__5459\,
            I => \N__5456\
        );

    \I__557\ : Odrv4
    port map (
            O => \N__5456\,
            I => \DUT.uart_inst0.N_81_mux_i_i_a5_0_4\
        );

    \I__556\ : InMux
    port map (
            O => \N__5453\,
            I => \N__5450\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__5450\,
            I => \DUT.uart_inst0.N_81_mux_i_i_0\
        );

    \I__554\ : CascadeMux
    port map (
            O => \N__5447\,
            I => \DUT.uart_inst0.N_81_mux_i_i_a5_0_5_cascade_\
        );

    \I__553\ : InMux
    port map (
            O => \N__5444\,
            I => \N__5441\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__5441\,
            I => \DUT.uart_inst0.N_81_mux_i_i_a5_1_5\
        );

    \I__551\ : InMux
    port map (
            O => \N__5438\,
            I => \N__5435\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__5435\,
            I => \N__5432\
        );

    \I__549\ : Odrv4
    port map (
            O => \N__5432\,
            I => \DUT.uart_inst0.m8_e_2\
        );

    \I__548\ : InMux
    port map (
            O => \N__5429\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_0_s1\
        );

    \I__547\ : InMux
    port map (
            O => \N__5426\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_1_s1\
        );

    \I__546\ : InMux
    port map (
            O => \N__5423\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_2_s1\
        );

    \I__545\ : InMux
    port map (
            O => \N__5420\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_3_s1\
        );

    \I__544\ : InMux
    port map (
            O => \N__5417\,
            I => \N__5414\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__5414\,
            I => \N__5411\
        );

    \I__542\ : Odrv4
    port map (
            O => \N__5411\,
            I => \DUT.uart_inst0.m8_e_3\
        );

    \I__541\ : InMux
    port map (
            O => \N__5408\,
            I => \N__5398\
        );

    \I__540\ : CascadeMux
    port map (
            O => \N__5407\,
            I => \N__5395\
        );

    \I__539\ : InMux
    port map (
            O => \N__5406\,
            I => \N__5384\
        );

    \I__538\ : InMux
    port map (
            O => \N__5405\,
            I => \N__5384\
        );

    \I__537\ : InMux
    port map (
            O => \N__5404\,
            I => \N__5384\
        );

    \I__536\ : InMux
    port map (
            O => \N__5403\,
            I => \N__5384\
        );

    \I__535\ : InMux
    port map (
            O => \N__5402\,
            I => \N__5384\
        );

    \I__534\ : InMux
    port map (
            O => \N__5401\,
            I => \N__5381\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__5398\,
            I => \N__5378\
        );

    \I__532\ : InMux
    port map (
            O => \N__5395\,
            I => \N__5375\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__5384\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_1\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__5381\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_1\
        );

    \I__529\ : Odrv12
    port map (
            O => \N__5378\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_1\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__5375\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_1\
        );

    \I__527\ : InMux
    port map (
            O => \N__5366\,
            I => \N__5363\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__5363\,
            I => \N__5360\
        );

    \I__525\ : Odrv4
    port map (
            O => \N__5360\,
            I => \DUT.uart_inst0.g0_i_a3_6\
        );

    \I__524\ : InMux
    port map (
            O => \N__5357\,
            I => \N__5354\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__5354\,
            I => \N__5351\
        );

    \I__522\ : Odrv4
    port map (
            O => \N__5351\,
            I => \DUT.uart_inst0.recv_state_ns_0_i_a2_0_0_3\
        );

    \I__521\ : InMux
    port map (
            O => \N__5348\,
            I => \N__5339\
        );

    \I__520\ : InMux
    port map (
            O => \N__5347\,
            I => \N__5339\
        );

    \I__519\ : InMux
    port map (
            O => \N__5346\,
            I => \N__5339\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__5339\,
            I => \DUT.uart_inst0.recv_stateZ0Z_3\
        );

    \I__517\ : InMux
    port map (
            O => \N__5336\,
            I => \N__5333\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__5333\,
            I => \DUT.uart_inst0.g0_0_0\
        );

    \I__515\ : InMux
    port map (
            O => \N__5330\,
            I => \N__5327\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__5327\,
            I => \DUT.uart_inst0.g0_0_1\
        );

    \I__513\ : CascadeMux
    port map (
            O => \N__5324\,
            I => \DUT.uart_inst0.N_81_mux_i_i_a5_0_4_0_cascade_\
        );

    \I__512\ : InMux
    port map (
            O => \N__5321\,
            I => \N__5318\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__5318\,
            I => \DUT.uart_inst0.N_35_0\
        );

    \I__510\ : CascadeMux
    port map (
            O => \N__5315\,
            I => \DUT.uart_inst0.g0_0_2_cascade_\
        );

    \I__509\ : InMux
    port map (
            O => \N__5312\,
            I => \N__5307\
        );

    \I__508\ : InMux
    port map (
            O => \N__5311\,
            I => \N__5303\
        );

    \I__507\ : InMux
    port map (
            O => \N__5310\,
            I => \N__5300\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__5307\,
            I => \N__5296\
        );

    \I__505\ : InMux
    port map (
            O => \N__5306\,
            I => \N__5292\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__5303\,
            I => \N__5287\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__5300\,
            I => \N__5287\
        );

    \I__502\ : InMux
    port map (
            O => \N__5299\,
            I => \N__5284\
        );

    \I__501\ : Span4Mux_h
    port map (
            O => \N__5296\,
            I => \N__5281\
        );

    \I__500\ : InMux
    port map (
            O => \N__5295\,
            I => \N__5278\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__5292\,
            I => \N__5273\
        );

    \I__498\ : Span4Mux_v
    port map (
            O => \N__5287\,
            I => \N__5273\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__5284\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_2\
        );

    \I__496\ : Odrv4
    port map (
            O => \N__5281\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_2\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__5278\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_2\
        );

    \I__494\ : Odrv4
    port map (
            O => \N__5273\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_2\
        );

    \I__493\ : InMux
    port map (
            O => \N__5264\,
            I => \N__5261\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__5261\,
            I => \DUT.uart_inst0.g0_i_a3_0_6\
        );

    \I__491\ : CascadeMux
    port map (
            O => \N__5258\,
            I => \DUT.uart_inst0.g0_i_a3_0_7_cascade_\
        );

    \I__490\ : CascadeMux
    port map (
            O => \N__5255\,
            I => \DUT.uart_inst0.N_6_0_cascade_\
        );

    \I__489\ : CascadeMux
    port map (
            O => \N__5252\,
            I => \N__5249\
        );

    \I__488\ : InMux
    port map (
            O => \N__5249\,
            I => \N__5246\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__5246\,
            I => \N__5243\
        );

    \I__486\ : Odrv12
    port map (
            O => \N__5243\,
            I => \DUT.uart_inst0.N_40\
        );

    \I__485\ : CascadeMux
    port map (
            O => \N__5240\,
            I => \N__5237\
        );

    \I__484\ : InMux
    port map (
            O => \N__5237\,
            I => \N__5231\
        );

    \I__483\ : InMux
    port map (
            O => \N__5236\,
            I => \N__5226\
        );

    \I__482\ : InMux
    port map (
            O => \N__5235\,
            I => \N__5226\
        );

    \I__481\ : InMux
    port map (
            O => \N__5234\,
            I => \N__5223\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__5231\,
            I => \N__5220\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__5226\,
            I => \N__5217\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__5223\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_3\
        );

    \I__477\ : Odrv4
    port map (
            O => \N__5220\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_3\
        );

    \I__476\ : Odrv4
    port map (
            O => \N__5217\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_3\
        );

    \I__475\ : CascadeMux
    port map (
            O => \N__5210\,
            I => \N__5205\
        );

    \I__474\ : InMux
    port map (
            O => \N__5209\,
            I => \N__5200\
        );

    \I__473\ : InMux
    port map (
            O => \N__5208\,
            I => \N__5197\
        );

    \I__472\ : InMux
    port map (
            O => \N__5205\,
            I => \N__5192\
        );

    \I__471\ : InMux
    port map (
            O => \N__5204\,
            I => \N__5192\
        );

    \I__470\ : CascadeMux
    port map (
            O => \N__5203\,
            I => \N__5189\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__5200\,
            I => \N__5180\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__5197\,
            I => \N__5180\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__5192\,
            I => \N__5180\
        );

    \I__466\ : InMux
    port map (
            O => \N__5189\,
            I => \N__5177\
        );

    \I__465\ : InMux
    port map (
            O => \N__5188\,
            I => \N__5174\
        );

    \I__464\ : InMux
    port map (
            O => \N__5187\,
            I => \N__5171\
        );

    \I__463\ : Span4Mux_v
    port map (
            O => \N__5180\,
            I => \N__5166\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__5177\,
            I => \N__5166\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__5174\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_0\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__5171\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_0\
        );

    \I__459\ : Odrv4
    port map (
            O => \N__5166\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_0\
        );

    \I__458\ : CEMux
    port map (
            O => \N__5159\,
            I => \N__5156\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__5156\,
            I => \N__5153\
        );

    \I__456\ : Span4Mux_h
    port map (
            O => \N__5153\,
            I => \N__5150\
        );

    \I__455\ : Odrv4
    port map (
            O => \N__5150\,
            I => \DUT.uart_inst0.recv_state_RNIL139CZ0Z_2\
        );

    \I__454\ : InMux
    port map (
            O => \N__5147\,
            I => \N__5144\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__5144\,
            I => \DUT.uart_inst0.g0_0_i_a3_0_3\
        );

    \I__452\ : CascadeMux
    port map (
            O => \N__5141\,
            I => \DUT.uart_inst0.g0_0_i_a3_0_4_cascade_\
        );

    \I__451\ : InMux
    port map (
            O => \N__5138\,
            I => \N__5135\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__5135\,
            I => \DUT.uart_inst0.g0_0\
        );

    \I__449\ : CascadeMux
    port map (
            O => \N__5132\,
            I => \DUT.uart_inst0.g0_i_a3_0_5_cascade_\
        );

    \I__448\ : InMux
    port map (
            O => \N__5129\,
            I => \N__5126\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__5126\,
            I => \DUT.uart_inst0.g0_i_a3_8\
        );

    \I__446\ : CascadeMux
    port map (
            O => \N__5123\,
            I => \DUT.uart_inst0.recv_state_ns_0_i_a2_0_2_3_cascade_\
        );

    \I__445\ : CascadeMux
    port map (
            O => \N__5120\,
            I => \DUT.uart_inst0.m16_N_3L3_1_cascade_\
        );

    \I__444\ : InMux
    port map (
            O => \N__5117\,
            I => \N__5114\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__5114\,
            I => \DUT.uart_inst0.rx_bits_remaining_RNO_4Z0Z_1\
        );

    \I__442\ : CascadeMux
    port map (
            O => \N__5111\,
            I => \DUT.uart_inst0.g0_i_a3_5_cascade_\
        );

    \I__441\ : InMux
    port map (
            O => \N__5108\,
            I => \N__5105\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__5105\,
            I => \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO\
        );

    \I__439\ : CascadeMux
    port map (
            O => \N__5102\,
            I => \DUT.uart_inst0.rx_bits_remaining_RNO_1Z0Z_1_cascade_\
        );

    \I__438\ : CascadeMux
    port map (
            O => \N__5099\,
            I => \DUT.uart_inst0.m5_1_1_cascade_\
        );

    \I__437\ : InMux
    port map (
            O => \N__5096\,
            I => \N__5093\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__5093\,
            I => \DUT.uart_inst0.N_6_0_0\
        );

    \I__435\ : CascadeMux
    port map (
            O => \N__5090\,
            I => \DUT.uart_inst0.N_6_0_0_cascade_\
        );

    \I__434\ : InMux
    port map (
            O => \N__5087\,
            I => \N__5084\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__5084\,
            I => \DUT.uart_inst0.N_15_mux_0\
        );

    \I__432\ : IoInMux
    port map (
            O => \N__5081\,
            I => \N__5078\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__5078\,
            I => \N__5075\
        );

    \I__430\ : Span12Mux_s9_v
    port map (
            O => \N__5075\,
            I => \N__5072\
        );

    \I__429\ : Span12Mux_v
    port map (
            O => \N__5072\,
            I => \N__5069\
        );

    \I__428\ : Odrv12
    port map (
            O => \N__5069\,
            I => \BTN_N_c\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_11_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DUT.uart_inst0.tx_clk_divider_cry_7\,
            carryinitout => \bfn_11_19_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DUT.uart_inst0.rx_clk_divider_1_cry_7\,
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DUT.uart_inst0.rx_clk_divider_1_cry_15\,
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_11_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_22_0_\
        );

    \IN_MUX_bfv_8_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_18_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_15_0_\
        );

    \wPllLocked_i_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5612\,
            GLOBALBUFFEROUTPUT => \wPllLocked_i_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \top_pll_inst.top_pll_inst_RNISDA2\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8363\,
            GLOBALBUFFEROUTPUT => \wPllLocked_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5108\,
            lcout => \wPllLocked\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_1_1_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010101010101"
        )
    port map (
            in0 => \N__5406\,
            in1 => \N__5096\,
            in2 => \N__8362\,
            in3 => \N__5117\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.rx_bits_remaining_RNO_1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_1_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100100111"
        )
    port map (
            in0 => \N__8353\,
            in1 => \N__5087\,
            in2 => \N__5102\,
            in3 => \N__7935\,
            lcout => \DUT.uart_inst0.rx_bits_remainingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13055\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_0_3_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__5404\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5204\,
            lcout => \DUT.uart_inst0.N_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNIFF651_2_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100010"
        )
    port map (
            in0 => \N__5529\,
            in1 => \N__10141\,
            in2 => \_gnd_net_\,
            in3 => \N__5657\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.m5_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNIO2V22_0_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010100100000"
        )
    port map (
            in0 => \N__5658\,
            in1 => \N__5208\,
            in2 => \N__5099\,
            in3 => \N__5402\,
            lcout => \DUT.uart_inst0.N_6_0_0\,
            ltout => \DUT.uart_inst0.N_6_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_0_1_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110101010101"
        )
    port map (
            in0 => \N__5403\,
            in1 => \N__5417\,
            in2 => \N__5090\,
            in3 => \N__5438\,
            lcout => \DUT.uart_inst0.N_15_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_2_2_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010110"
        )
    port map (
            in0 => \N__5299\,
            in1 => \N__5405\,
            in2 => \N__5210\,
            in3 => \N__5530\,
            lcout => \DUT.uart_inst0.N_35_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_1_3_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__5295\,
            in1 => \N__5401\,
            in2 => \N__5240\,
            in3 => \N__5209\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.recv_state_ns_0_i_a2_0_2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_3_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5123\,
            in3 => \N__5659\,
            lcout => \DUT.uart_inst0.recv_state_ns_0_i_a2_0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_5_1_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6320\,
            in1 => \N__6731\,
            in2 => \_gnd_net_\,
            in3 => \N__6243\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.m16_N_3L3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_4_1_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6136\,
            in1 => \N__6562\,
            in2 => \N__5120\,
            in3 => \N__6795\,
            lcout => \DUT.uart_inst0.rx_bits_remaining_RNO_4Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_6_2_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__5511\,
            in1 => \N__6242\,
            in2 => \N__10171\,
            in3 => \N__6730\,
            lcout => \DUT.uart_inst0.m9_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_3_4_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6244\,
            in1 => \N__6321\,
            in2 => \N__6142\,
            in3 => \N__6563\,
            lcout => \DUT.uart_inst0.N_81_mux_i_i_a5_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_4_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__12060\,
            in1 => \N__6058\,
            in2 => \_gnd_net_\,
            in3 => \N__10041\,
            lcout => \DUT.uart_inst0.N_81_mux_i_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_6_2_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010001000"
        )
    port map (
            in0 => \N__8336\,
            in1 => \N__5642\,
            in2 => \N__10172\,
            in3 => \N__5507\,
            lcout => \DUT.uart_inst0.g0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_9_2_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6427\,
            in1 => \N__6491\,
            in2 => \N__5203\,
            in3 => \N__6713\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g0_i_a3_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_4_2_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__5366\,
            in1 => \N__5236\,
            in2 => \N__5111\,
            in3 => \N__5312\,
            lcout => \DUT.uart_inst0.g0_i_a3_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNI69LM2_0_0_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__6553\,
            in1 => \N__6712\,
            in2 => \N__6252\,
            in3 => \N__6314\,
            lcout => \DUT.uart_inst0.g0_0_i_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_0_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__10165\,
            in1 => \N__9976\,
            in2 => \_gnd_net_\,
            in3 => \N__7142\,
            lcout => \DUT.uart_inst0.recv_state_ns_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_2_2_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5235\,
            in1 => \N__6316\,
            in2 => \N__6566\,
            in3 => \N__6249\,
            lcout => \DUT.uart_inst0.g0_i_a3_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_7_2_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6315\,
            in1 => \N__6126\,
            in2 => \N__6796\,
            in3 => \N__6554\,
            lcout => \DUT.uart_inst0.m9_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNIS6O94_0_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__6788\,
            in1 => \_gnd_net_\,
            in2 => \N__6141\,
            in3 => \N__5147\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g0_0_i_a3_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNIL139C_2_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__5138\,
            in1 => \N__5669\,
            in2 => \N__5141\,
            in3 => \N__7937\,
            lcout => \DUT.uart_inst0.recv_state_RNIL139CZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNIBTG71_2_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110000000000"
        )
    port map (
            in0 => \N__10169\,
            in1 => \N__5644\,
            in2 => \N__5528\,
            in3 => \N__12066\,
            lcout => \DUT.uart_inst0.g0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_8_2_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5310\,
            in1 => \N__5408\,
            in2 => \_gnd_net_\,
            in3 => \N__6789\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g0_i_a3_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_3_2_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6130\,
            in1 => \N__5187\,
            in2 => \N__5132\,
            in3 => \N__6734\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g0_i_a3_0_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_2_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111101010101"
        )
    port map (
            in0 => \N__5129\,
            in1 => \N__5264\,
            in2 => \N__5258\,
            in3 => \N__7936\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_2_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010000000"
        )
    port map (
            in0 => \N__8352\,
            in1 => \N__5645\,
            in2 => \N__5255\,
            in3 => \N__5570\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13048\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_3_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101001"
        )
    port map (
            in0 => \N__5234\,
            in1 => \N__5311\,
            in2 => \N__5252\,
            in3 => \N__5534\,
            lcout => \DUT.uart_inst0.rx_bits_remainingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13043\,
            ce => \N__5159\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_0_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5533\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5188\,
            lcout => \DUT.uart_inst0.rx_bits_remainingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13043\,
            ce => \N__5159\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7418\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13037\,
            ce => \N__7487\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7374\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13037\,
            ce => \N__7487\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7326\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13037\,
            ce => \N__7487\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7809\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13037\,
            ce => \N__7487\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7754\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13037\,
            ce => \N__7487\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7703\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13037\,
            ce => \N__7487\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7652\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13037\,
            ce => \N__7487\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10491\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13037\,
            ce => \N__7487\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13088\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13032\,
            ce => \N__7205\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13277\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13032\,
            ce => \N__7205\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12497\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13032\,
            ce => \N__7205\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12421\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13032\,
            ce => \N__7205\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12381\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13032\,
            ce => \N__7205\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13130\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13032\,
            ce => \N__7205\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13209\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13032\,
            ce => \N__7205\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13319\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13032\,
            ce => \N__7205\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_7_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7422\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13027\,
            ce => \N__10441\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7376\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13027\,
            ce => \N__10441\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_7_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7327\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13027\,
            ce => \N__10441\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_7_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7758\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13027\,
            ce => \N__10441\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_7_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7707\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13027\,
            ce => \N__10441\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7655\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13027\,
            ce => \N__10441\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_7_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7810\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13021\,
            ce => \N__10437\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_0_2_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100000000"
        )
    port map (
            in0 => \N__7913\,
            in1 => \N__6334\,
            in2 => \N__6869\,
            in3 => \N__5330\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_2_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110011001100"
        )
    port map (
            in0 => \N__5321\,
            in1 => \N__5306\,
            in2 => \N__5315\,
            in3 => \N__6161\,
            lcout => \DUT.uart_inst0.rx_bits_remainingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13054\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_6_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__8358\,
            in1 => \N__5348\,
            in2 => \N__10140\,
            in3 => \N__6042\,
            lcout => \DUT.wRcvd\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13054\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_3_1_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6852\,
            in1 => \N__6428\,
            in2 => \N__6959\,
            in3 => \N__6493\,
            lcout => \DUT.uart_inst0.m8_e_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_10_2_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6993\,
            in1 => \N__6955\,
            in2 => \N__5407\,
            in3 => \N__6851\,
            lcout => \DUT.uart_inst0.g0_i_a3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_2_2_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__5531\,
            in1 => \N__10116\,
            in2 => \_gnd_net_\,
            in3 => \N__5663\,
            lcout => \DUT.uart_inst0.rx_countdown_RNO_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_5_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__10115\,
            in1 => \N__5346\,
            in2 => \_gnd_net_\,
            in3 => \N__5532\,
            lcout => \DUT.uart_inst0.N_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_3_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__5347\,
            in1 => \N__8357\,
            in2 => \N__6047\,
            in3 => \N__5357\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13054\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_3_2_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010101000"
        )
    port map (
            in0 => \N__5336\,
            in1 => \N__6697\,
            in2 => \N__6263\,
            in3 => \N__6793\,
            lcout => \DUT.uart_inst0.g0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_1_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111110111"
        )
    port map (
            in0 => \N__12059\,
            in1 => \N__9968\,
            in2 => \N__10161\,
            in3 => \N__5522\,
            lcout => \DUT.uart_inst0.N_81_mux_i_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_3_1_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6132\,
            in1 => \N__6792\,
            in2 => \N__6333\,
            in3 => \N__6561\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_81_mux_i_i_a5_0_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_1_1_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6699\,
            in1 => \N__9565\,
            in2 => \N__5324\,
            in3 => \N__6248\,
            lcout => \DUT.uart_inst0.N_81_mux_i_i_a5_0_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_1_4_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__10039\,
            in1 => \N__5462\,
            in2 => \N__6729\,
            in3 => \N__6794\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_81_mux_i_i_a5_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_4_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100010001"
        )
    port map (
            in0 => \N__5453\,
            in1 => \N__5444\,
            in2 => \N__5447\,
            in3 => \N__7917\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13052\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_4_2_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6131\,
            in1 => \N__6560\,
            in2 => \N__6254\,
            in3 => \N__6791\,
            lcout => \DUT.uart_inst0.N_13_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_2_4_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__6698\,
            in1 => \N__5960\,
            in2 => \N__10035\,
            in3 => \N__6853\,
            lcout => \DUT.uart_inst0.N_81_mux_i_i_a5_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_2_1_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__7002\,
            in1 => \_gnd_net_\,
            in2 => \N__6711\,
            in3 => \_gnd_net_\,
            lcout => \DUT.uart_inst0.m8_e_2\,
            ltout => OPEN,
            carryin => \bfn_8_15_0_\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_0_s1_c_RNIKPDT_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12747\,
            in2 => \N__6492\,
            in3 => \N__5429\,
            lcout => \DUT.uart_inst0.rx_countdown_3_s1_1\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_countdown_3_cry_0_s1\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNIMVNN_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6858\,
            in2 => \N__12807\,
            in3 => \N__5426\,
            lcout => \DUT.uart_inst0.rx_countdown_3_s1_2\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_countdown_3_cry_1_s1\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_2_s1_c_RNIO52I_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12751\,
            in2 => \N__6947\,
            in3 => \N__5423\,
            lcout => \DUT.uart_inst0.rx_countdown_3_s1_3\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_countdown_3_cry_2_s1\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_3_s1_c_RNIQBCS_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12752\,
            in2 => \N__7019\,
            in3 => \N__5420\,
            lcout => \DUT.uart_inst0.rx_countdown_3_s1_4\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_countdown_3_cry_3_s1\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_4_s1_c_RNISHMM_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6400\,
            in2 => \_gnd_net_\,
            in3 => \N__5585\,
            lcout => \DUT.uart_inst0.rx_countdown_3_s1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_1_2_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__5582\,
            in1 => \N__5576\,
            in2 => \N__5546\,
            in3 => \N__7899\,
            lcout => \DUT.uart_inst0.N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_1_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100001011"
        )
    port map (
            in0 => \N__7900\,
            in1 => \N__6182\,
            in2 => \N__5564\,
            in3 => \N__5555\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13049\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_12_2_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6479\,
            in1 => \N__6871\,
            in2 => \N__6420\,
            in3 => \N__6686\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.m4_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_5_2_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__5468\,
            in1 => \N__7030\,
            in2 => \N__5549\,
            in3 => \N__6940\,
            lcout => \DUT.uart_inst0.N_18_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_0_1_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__6480\,
            in1 => \N__7925\,
            in2 => \N__10046\,
            in3 => \N__6251\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_297_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_1_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5537\,
            in3 => \N__9541\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13044\,
            ce => \N__12000\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_11_2_LC_8_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__5506\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10146\,
            lcout => \DUT.uart_inst0.N_15_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNIPHLT1_5_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6685\,
            in1 => \N__6939\,
            in2 => \N__6424\,
            in3 => \N__6478\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g0_0_i_a3_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNI7CGS2_2_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__7031\,
            in1 => \_gnd_net_\,
            in2 => \N__5672\,
            in3 => \N__6872\,
            lcout => \DUT.uart_inst0.g0_0_i_a3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNIEQQU_5_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6396\,
            in2 => \_gnd_net_\,
            in3 => \N__6477\,
            lcout => \DUT.uart_inst0.N_13_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNI8P9F_2_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12064\,
            in2 => \_gnd_net_\,
            in3 => \N__5643\,
            lcout => \DUT.uart_inst0.m11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNISAK33_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6565\,
            in1 => \N__6140\,
            in2 => \N__6335\,
            in3 => \N__6250\,
            lcout => \DUT.uart_inst0.m10_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.wPllLocked_i_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12065\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \wPllLocked_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7148\,
            in2 => \N__7076\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_18_0_\,
            carryout => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_1_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7233\,
            in2 => \N__5684\,
            in3 => \N__5591\,
            lcout => \DUT.fifo_rx_inst.rFifoCountZ0Z_1\,
            ltout => OPEN,
            carryin => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0\,
            carryout => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1\,
            clk => \N__13038\,
            ce => 'H',
            sr => \N__10527\
        );

    \DUT.fifo_rx_inst.rFifoCount_2_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5696\,
            in2 => \_gnd_net_\,
            in3 => \N__5588\,
            lcout => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13038\,
            ce => 'H',
            sr => \N__10527\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI96D91_2_1_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5800\,
            in1 => \N__7130\,
            in2 => \N__5833\,
            in3 => \N__7271\,
            lcout => \DUT.fifo_rx_inst.rFifoData_awe3\,
            ltout => \DUT.fifo_rx_inst.rFifoData_awe3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1_1_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__12070\,
            in1 => \_gnd_net_\,
            in2 => \N__5702\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.un1_i11_i\,
            ltout => \DUT.fifo_rx_inst.un1_i11_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_0_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__5822\,
            in1 => \_gnd_net_\,
            in2 => \N__5699\,
            in3 => \N__5857\,
            lcout => \DUT.fifo_rx_inst.rWritePtrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13033\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNO_0_2_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000110"
        )
    port map (
            in0 => \N__10653\,
            in1 => \N__7273\,
            in2 => \N__7141\,
            in3 => \N__8223\,
            lcout => \DUT.fifo_rx_inst.un1_rFifoCount_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__7272\,
            in1 => \N__7229\,
            in2 => \_gnd_net_\,
            in3 => \N__7072\,
            lcout => \N_92_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_1_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000100010"
        )
    port map (
            in0 => \N__5801\,
            in1 => \N__5690\,
            in2 => \N__5834\,
            in3 => \N__5858\,
            lcout => \DUT.fifo_rx_inst.rWritePtrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13033\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNIK3G92_1_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__7131\,
            in1 => \N__10652\,
            in2 => \N__7235\,
            in3 => \N__8222\,
            lcout => \DUT.fifo_rx_inst.rFifoCount_RNIK3G92Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_8_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__5803\,
            in1 => \_gnd_net_\,
            in2 => \N__5840\,
            in3 => \N__5855\,
            lcout => \DUT.fifo_rx_inst.rFifoData_awe0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_8_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7106\,
            in2 => \_gnd_net_\,
            in3 => \N__7274\,
            lcout => \DUT.fifo_rx_inst.rWritePtr16\,
            ltout => \DUT.fifo_rx_inst.rWritePtr16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_8_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5835\,
            in2 => \N__5675\,
            in3 => \N__5802\,
            lcout => \DUT.fifo_rx_inst.rFifoData_awe1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_0_1_LC_8_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__11437\,
            in1 => \N__11606\,
            in2 => \_gnd_net_\,
            in3 => \N__11686\,
            lcout => \DUT.uart_inst0.N_8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_8_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__5856\,
            in1 => \N__5839\,
            in2 => \_gnd_net_\,
            in3 => \N__5804\,
            lcout => \DUT.fifo_rx_inst.rFifoData_awe2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_8_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__8977\,
            in1 => \N__5783\,
            in2 => \N__6017\,
            in3 => \N__8182\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rTxByte_esr_6_LC_8_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__9017\,
            in1 => \N__7610\,
            in2 => \N__5777\,
            in3 => \N__5720\,
            lcout => \rTxByteZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13022\,
            ce => \N__8877\,
            sr => \N__8844\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_8_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__5765\,
            in1 => \N__9010\,
            in2 => \N__5996\,
            in3 => \N__8197\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rTxByte_esr_4_LC_8_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__9015\,
            in1 => \N__5756\,
            in2 => \N__5747\,
            in3 => \N__7715\,
            lcout => \rTxByteZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13022\,
            ce => \N__8877\,
            sr => \N__8844\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_8_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__5744\,
            in1 => \N__9011\,
            in2 => \N__5984\,
            in3 => \N__8198\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rTxByte_esr_5_LC_8_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__9016\,
            in1 => \N__7664\,
            in2 => \N__5738\,
            in3 => \N__5735\,
            lcout => \rTxByteZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13022\,
            ce => \N__8877\,
            sr => \N__8844\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_8_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__5726\,
            in1 => \N__9009\,
            in2 => \N__5972\,
            in3 => \N__8195\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_8_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__8196\,
            in1 => \N__6005\,
            in2 => \N__9025\,
            in3 => \N__5711\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rTxByte_esr_3_LC_8_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__7766\,
            in1 => \N__5948\,
            in2 => \N__5939\,
            in3 => \N__9018\,
            lcout => \rTxByteZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13022\,
            ce => \N__8877\,
            sr => \N__8844\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_8_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__8194\,
            in1 => \N__5873\,
            in2 => \N__5936\,
            in3 => \N__9019\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rTxByte_esr_0_LC_8_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__7385\,
            in1 => \N__5927\,
            in2 => \N__5915\,
            in3 => \N__9005\,
            lcout => \rTxByteZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13016\,
            ce => \N__8879\,
            sr => \N__8852\
        );

    \rTxByte_esr_7_LC_8_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__5912\,
            in1 => \N__7556\,
            in2 => \N__7598\,
            in3 => \N__9020\,
            lcout => \rTxByteZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13016\,
            ce => \N__8879\,
            sr => \N__8852\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_8_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__5900\,
            in1 => \N__9004\,
            in2 => \N__5867\,
            in3 => \N__8193\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rTxByte_esr_2_LC_8_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000011"
        )
    port map (
            in0 => \N__5894\,
            in1 => \N__5882\,
            in2 => \N__9024\,
            in3 => \N__7280\,
            lcout => \rTxByteZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13016\,
            ce => \N__8879\,
            sr => \N__8852\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_8_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7427\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13011\,
            ce => \N__7511\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_8_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7375\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13011\,
            ce => \N__7511\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_8_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7328\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13011\,
            ce => \N__7511\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_8_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7814\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13011\,
            ce => \N__7511\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_8_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7759\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13011\,
            ce => \N__7511\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_8_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7708\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13011\,
            ce => \N__7511\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_8_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7654\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13011\,
            ce => \N__7511\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_8_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10492\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13011\,
            ce => \N__7511\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_4_4_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6954\,
            in1 => \N__6425\,
            in2 => \N__7018\,
            in3 => \N__6494\,
            lcout => \DUT.uart_inst0.N_81_mux_i_i_a5_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_4_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__6143\,
            in1 => \N__9938\,
            in2 => \N__7923\,
            in3 => \N__6998\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13053\,
            ce => \N__11980\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_4_2_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6994\,
            in2 => \_gnd_net_\,
            in3 => \N__6953\,
            lcout => \DUT.uart_inst0.G_9_i_o4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001000011"
        )
    port map (
            in0 => \N__5954\,
            in1 => \N__7895\,
            in2 => \N__6733\,
            in3 => \N__6344\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.G_21_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_2_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__6176\,
            in1 => \N__9566\,
            in2 => \N__6170\,
            in3 => \N__6068\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13053\,
            ce => \N__11980\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_1_2_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000010"
        )
    port map (
            in0 => \N__6077\,
            in1 => \N__7894\,
            in2 => \N__6732\,
            in3 => \N__6167\,
            lcout => \DUT.uart_inst0.g0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_3_s1_c_RNIMT2J1_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6125\,
            in2 => \_gnd_net_\,
            in3 => \N__6790\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.G_16_i_a3_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNIA4I1B_0_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111101010101"
        )
    port map (
            in0 => \N__6503\,
            in1 => \N__6269\,
            in2 => \N__6155\,
            in3 => \N__7893\,
            lcout => \DUT.uart_inst0.N_45\,
            ltout => \DUT.uart_inst0.N_45_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_5_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__8328\,
            in1 => \_gnd_net_\,
            in2 => \N__6152\,
            in3 => \N__6149\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13050\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_5_2_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__6124\,
            in1 => \N__6558\,
            in2 => \N__6253\,
            in3 => \N__6696\,
            lcout => \DUT.uart_inst0.N_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNI7H9R3_10_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7958\,
            in1 => \N__7829\,
            in2 => \N__7823\,
            in3 => \N__7943\,
            lcout => \DUT.uart_inst0.un2_rx_clk_divider_0\,
            ltout => \DUT.uart_inst0.un2_rx_clk_divider_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__10019\,
            in1 => \N__6325\,
            in2 => \N__6071\,
            in3 => \N__6854\,
            lcout => \DUT.uart_inst0.G_21_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_0_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111111111111"
        )
    port map (
            in0 => \N__6062\,
            in1 => \N__6046\,
            in2 => \N__8348\,
            in3 => \N__6029\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13050\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNI69LM2_0_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__6238\,
            in1 => \N__6559\,
            in2 => \N__6332\,
            in3 => \N__6695\,
            lcout => \DUT.uart_inst0.G_16_i_a3_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_5_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__6781\,
            in1 => \N__9937\,
            in2 => \N__6426\,
            in3 => \N__7920\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13045\,
            ce => \N__11989\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_7_2_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6412\,
            in2 => \_gnd_net_\,
            in3 => \N__6487\,
            lcout => \DUT.uart_inst0.g1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_0_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__6688\,
            in1 => \N__9936\,
            in2 => \_gnd_net_\,
            in3 => \N__7918\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13045\,
            ce => \N__11989\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNI2GC23_0_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001111"
        )
    port map (
            in0 => \N__6234\,
            in1 => \N__6687\,
            in2 => \N__6890\,
            in3 => \N__6780\,
            lcout => \DUT.uart_inst0.N_15_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_3_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111010111"
        )
    port map (
            in0 => \N__9564\,
            in1 => \N__9181\,
            in2 => \N__9167\,
            in3 => \N__7919\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13045\,
            ce => \N__11989\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIMQ571_1_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9180\,
            in1 => \N__9646\,
            in2 => \N__9491\,
            in3 => \N__9219\,
            lcout => \DUT.uart_inst0.un2_rx_clk_divider_a_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__9220\,
            in1 => \N__9206\,
            in2 => \_gnd_net_\,
            in3 => \N__9580\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13045\,
            ce => \N__11989\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_2_1_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__9539\,
            in1 => \N__6405\,
            in2 => \N__6575\,
            in3 => \N__6483\,
            lcout => \DUT.uart_inst0.N_81_mux_i_i_a5_1_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_4_1_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6863\,
            in1 => \N__6937\,
            in2 => \N__7034\,
            in3 => \N__6679\,
            lcout => \DUT.uart_inst0.N_81_mux_i_i_a5_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_0_3_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100001101"
        )
    port map (
            in0 => \N__6938\,
            in1 => \N__7924\,
            in2 => \N__10045\,
            in3 => \N__6564\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_300_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6509\,
            in3 => \N__9540\,
            lcout => \DUT.uart_inst0.rx_countdownZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13041\,
            ce => \N__11993\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNI237O_0_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10145\,
            in2 => \_gnd_net_\,
            in3 => \N__9969\,
            lcout => \DUT.uart_inst0.N_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNIPHLT1_2_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6862\,
            in1 => \N__6935\,
            in2 => \N__7032\,
            in3 => \N__6678\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.G_16_i_a3_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNI7CGS2_5_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6404\,
            in2 => \N__6506\,
            in3 => \N__6481\,
            lcout => \DUT.uart_inst0.G_16_i_a3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_3_2_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6482\,
            in1 => \N__6419\,
            in2 => \N__7033\,
            in3 => \N__6936\,
            lcout => \DUT.uart_inst0.N_11_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_0_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__8568\,
            in1 => \N__7043\,
            in2 => \_gnd_net_\,
            in3 => \N__8485\,
            lcout => \DUT.fifo_tx_inst.rWritePtrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13039\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_RNIN79A_2_1_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__8530\,
            in1 => \N__10663\,
            in2 => \N__8570\,
            in3 => \N__10571\,
            lcout => \DUT.fifo_tx_inst.rFifoData_awe3\,
            ltout => \DUT.fifo_tx_inst.rFifoData_awe3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_RNIJLJC_1_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7046\,
            in3 => \N__12061\,
            lcout => \DUT.fifo_tx_inst.un1_i11_i\,
            ltout => \DUT.fifo_tx_inst.un1_i11_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_1_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__8486\,
            in1 => \N__8569\,
            in2 => \N__7037\,
            in3 => \N__8531\,
            lcout => \DUT.fifo_tx_inst.rWritePtrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13039\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNI323D2_2_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__7029\,
            in1 => \N__6941\,
            in2 => \N__6889\,
            in3 => \N__6870\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNIV8RM6_0_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__6800\,
            in1 => \N__6719\,
            in2 => \N__6605\,
            in3 => \N__6602\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_11_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNIG3R3E_2_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000100000"
        )
    port map (
            in0 => \N__6596\,
            in1 => \N__6587\,
            in2 => \N__6578\,
            in3 => \N__7926\,
            lcout => \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_0_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7351\,
            lcout => \DUT.wRxByte_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13034\,
            ce => \N__7160\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_1_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7303\,
            lcout => \DUT.wRxByte_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13034\,
            ce => \N__7160\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_2_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7787\,
            lcout => \DUT.wRxByte_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13034\,
            ce => \N__7160\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_3_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7731\,
            lcout => \DUT.wRxByte_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13034\,
            ce => \N__7160\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_4_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7680\,
            lcout => \DUT.wRxByte_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13034\,
            ce => \N__7160\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_5_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7628\,
            lcout => \DUT.wRxByte_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13034\,
            ce => \N__7160\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_6_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10469\,
            lcout => \DUT.wRxByte_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13034\,
            ce => \N__7160\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_7_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10111\,
            lcout => \DUT.wRxByte_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13034\,
            ce => \N__7160\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNIPTFQ1_0_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110011001"
        )
    port map (
            in0 => \N__7138\,
            in1 => \N__10647\,
            in2 => \_gnd_net_\,
            in3 => \N__8221\,
            lcout => \DUT.fifo_rx_inst.N_87\,
            ltout => \DUT.fifo_rx_inst.N_87_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100001111"
        )
    port map (
            in0 => \N__7071\,
            in1 => \N__7139\,
            in2 => \N__7151\,
            in3 => \N__7265\,
            lcout => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_0_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100000000111"
        )
    port map (
            in0 => \N__7266\,
            in1 => \N__7140\,
            in2 => \N__7088\,
            in3 => \N__7070\,
            lcout => \DUT.fifo_rx_inst.rFifoCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13028\,
            ce => 'H',
            sr => \N__10525\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_0_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__7264\,
            in1 => \N__7228\,
            in2 => \_gnd_net_\,
            in3 => \N__7068\,
            lcout => \DUT.fifo_rx_inst.N_92\,
            ltout => \DUT.fifo_rx_inst.N_92_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rReadPtr_RNI8B9Q1_0_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__10648\,
            in1 => \_gnd_net_\,
            in2 => \N__7079\,
            in3 => \N__8163\,
            lcout => \DUT.fifo_rx_inst.CO0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rRxRead_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__7069\,
            in1 => \N__7267\,
            in2 => \_gnd_net_\,
            in3 => \N__7234\,
            lcout => \rRxReadZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13028\,
            ce => 'H',
            sr => \N__10525\
        );

    \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__8575\,
            in1 => \N__8534\,
            in2 => \_gnd_net_\,
            in3 => \N__8476\,
            lcout => \DUT.fifo_tx_inst.rFifoData_awe2\,
            ltout => \DUT.fifo_tx_inst.rFifoData_awe2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_2_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7193\,
            in3 => \N__7181\,
            lcout => \DUT.fifo_tx_inst.rFifoDataro_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13023\,
            ce => 'H',
            sr => \N__10524\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_3_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__7190\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12523\,
            lcout => \DUT.fifo_tx_inst.rFifoDataro_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13023\,
            ce => 'H',
            sr => \N__10524\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111101111111"
        )
    port map (
            in0 => \N__10901\,
            in1 => \N__7189\,
            in2 => \N__10852\,
            in3 => \N__7180\,
            lcout => \DUT.rFifoDataror_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_1_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8437\,
            in2 => \_gnd_net_\,
            in3 => \N__12861\,
            lcout => \DUT.fifo_tx_inst.rFifoDataro_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13023\,
            ce => 'H',
            sr => \N__10524\
        );

    \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_1_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__8574\,
            in1 => \N__8533\,
            in2 => \_gnd_net_\,
            in3 => \N__8475\,
            lcout => \DUT.fifo_tx_inst.rFifoData_awe0\,
            ltout => \DUT.fifo_tx_inst.rFifoData_awe0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_0_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7172\,
            in3 => \N__8450\,
            lcout => \DUT.fifo_tx_inst.rFifoDataro_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13023\,
            ce => 'H',
            sr => \N__10524\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_0_RNI0AQO1_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110111"
        )
    port map (
            in0 => \N__8161\,
            in1 => \N__7495\,
            in2 => \N__8968\,
            in3 => \N__7168\,
            lcout => \DUT.fifo_rx_inst.rTxByte_42_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_0_LC_9_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__7169\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10424\,
            lcout => \DUT.fifo_rx_inst.rFifoDataro_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13017\,
            ce => 'H',
            sr => \N__10523\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_1_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7507\,
            in2 => \_gnd_net_\,
            in3 => \N__7496\,
            lcout => \DUT.fifo_rx_inst.rFifoDataro_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13017\,
            ce => 'H',
            sr => \N__10523\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_3_LC_9_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__7469\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7585\,
            lcout => \DUT.fifo_rx_inst.rFifoDataro_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13017\,
            ce => 'H',
            sr => \N__10523\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_2_LC_9_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7459\,
            in2 => \_gnd_net_\,
            in3 => \N__7480\,
            lcout => \DUT.fifo_rx_inst.rFifoDataro_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13017\,
            ce => 'H',
            sr => \N__10523\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100111111"
        )
    port map (
            in0 => \N__7468\,
            in1 => \N__8946\,
            in2 => \N__7460\,
            in3 => \N__8162\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rTxByte_42_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_0_RNIHJV05_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111010101"
        )
    port map (
            in0 => \N__12072\,
            in1 => \N__7448\,
            in2 => \N__7442\,
            in3 => \N__8228\,
            lcout => \rFifoDatarff_0_RNIHJV05\,
            ltout => \rFifoDatarff_0_RNIHJV05_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNI250E6_0_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__7439\,
            in1 => \_gnd_net_\,
            in2 => \N__7430\,
            in3 => \_gnd_net_\,
            lcout => \N_92_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7426\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13012\,
            ce => \N__7589\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7370\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13012\,
            ce => \N__7589\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7319\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13012\,
            ce => \N__7589\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7802\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13012\,
            ce => \N__7589\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7760\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13012\,
            ce => \N__7589\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_9_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7709\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13012\,
            ce => \N__7589\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_9_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7653\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13012\,
            ce => \N__7589\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_9_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10490\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13012\,
            ce => \N__7589\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_9_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__8192\,
            in1 => \N__10451\,
            in2 => \N__9026\,
            in3 => \N__7562\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ft2232h_inst.rFifoState_1_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__11121\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11010\,
            lcout => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13051\,
            ce => 'H',
            sr => \N__10529\
        );

    \fifo_inst.ft2232h_inst.rRx_n_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111110101110000"
        )
    port map (
            in0 => \N__11011\,
            in1 => \N__11122\,
            in2 => \N__8819\,
            in3 => \N__7522\,
            lcout => \P1A3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13051\,
            ce => 'H',
            sr => \N__10529\
        );

    \fifo_inst.ft2232h_inst.rFifoState_2_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7949\,
            lcout => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13051\,
            ce => 'H',
            sr => \N__10529\
        );

    \DUT.uart_inst0.rx_clk_divider_RNI6B671_5_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9090\,
            in1 => \N__9114\,
            in2 => \N__9065\,
            in3 => \N__9141\,
            lcout => \DUT.uart_inst0.un2_rx_clk_divider_a_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_7_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__9092\,
            in1 => \N__9074\,
            in2 => \_gnd_net_\,
            in3 => \N__9591\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13046\,
            ce => \N__11976\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_5_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110011111"
        )
    port map (
            in0 => \N__9128\,
            in1 => \N__9142\,
            in2 => \N__9613\,
            in3 => \N__7921\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13046\,
            ce => \N__11976\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_6_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101110111111"
        )
    port map (
            in0 => \N__7922\,
            in1 => \N__9599\,
            in2 => \N__9119\,
            in3 => \N__9101\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13046\,
            ce => \N__11976\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_8_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000001010000"
        )
    port map (
            in0 => \N__9063\,
            in1 => \_gnd_net_\,
            in2 => \N__9612\,
            in3 => \N__9047\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13046\,
            ce => \N__11976\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_11_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__9359\,
            in1 => \N__9341\,
            in2 => \_gnd_net_\,
            in3 => \N__9590\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13046\,
            ce => \N__11976\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIB99J_10_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9357\,
            in1 => \N__9384\,
            in2 => \N__9416\,
            in3 => \N__9676\,
            lcout => \DUT.uart_inst0.un2_rx_clk_divider_a_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_9_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9414\,
            in2 => \N__9398\,
            in3 => \N__9595\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13046\,
            ce => \N__11976\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNI3ALC_17_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9276\,
            in1 => \N__9303\,
            in2 => \N__9698\,
            in3 => \N__9327\,
            lcout => \DUT.uart_inst0.un2_rx_clk_divider_a_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_13_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000001010000"
        )
    port map (
            in0 => \N__9328\,
            in1 => \_gnd_net_\,
            in2 => \N__9614\,
            in3 => \N__9314\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13042\,
            ce => \N__11978\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_14_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__9305\,
            in1 => \N__9287\,
            in2 => \_gnd_net_\,
            in3 => \N__9605\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13042\,
            ce => \N__11978\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_15_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__9606\,
            in1 => \N__9263\,
            in2 => \_gnd_net_\,
            in3 => \N__9277\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13042\,
            ce => \N__11978\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_0_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__8590\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9600\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13042\,
            ce => \N__11978\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIJI4K1_16_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__9252\,
            in1 => \N__8589\,
            in2 => \_gnd_net_\,
            in3 => \N__7964\,
            lcout => \DUT.uart_inst0.un2_rx_clk_divider_a_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_16_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__9254\,
            in1 => \N__9236\,
            in2 => \_gnd_net_\,
            in3 => \N__9607\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13042\,
            ce => \N__11978\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_10_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__9601\,
            in1 => \N__9368\,
            in2 => \_gnd_net_\,
            in3 => \N__9386\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13042\,
            ce => \N__11978\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__9734\,
            in1 => \N__9782\,
            in2 => \_gnd_net_\,
            in3 => \N__9856\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.un1_N_5_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_3_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110101111101"
        )
    port map (
            in0 => \N__7970\,
            in1 => \N__9897\,
            in2 => \N__7952\,
            in3 => \N__9752\,
            lcout => \DUT.uart_inst0.tx_bits_remainingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13040\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_5_3_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__11414\,
            in1 => \N__11834\,
            in2 => \N__11593\,
            in3 => \N__11924\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g0_i_o6_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7979\,
            in2 => \N__7982\,
            in3 => \N__11885\,
            lcout => \DUT.uart_inst0.g0_i_a6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_6_3_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__9732\,
            in1 => \N__9780\,
            in2 => \N__9901\,
            in3 => \N__9852\,
            lcout => \DUT.uart_inst0.g0_i_o6_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_4_2_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9781\,
            in1 => \N__9896\,
            in2 => \N__9857\,
            in3 => \N__9733\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_139_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_0_2_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__11415\,
            in1 => \N__11536\,
            in2 => \N__7973\,
            in3 => \N__11777\,
            lcout => \DUT.uart_inst0.g0_11_a4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNO_1_3_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__11537\,
            in1 => \N__11416\,
            in2 => \N__12073\,
            in3 => \N__11680\,
            lcout => \DUT.uart_inst0.tx_bits_remaining_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_0_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__8123\,
            in1 => \N__10180\,
            in2 => \_gnd_net_\,
            in3 => \N__9424\,
            lcout => \DUT.tx_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13035\,
            ce => 'H',
            sr => \N__10526\
        );

    \DUT.uart_inst0.tx_state_1_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__9425\,
            in1 => \N__11408\,
            in2 => \N__10184\,
            in3 => \N__10235\,
            lcout => \DUT.uart_inst0.tx_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13035\,
            ce => 'H',
            sr => \N__10526\
        );

    \DUT.uart_inst0.tx_data_0_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__10388\,
            in1 => \N__11545\,
            in2 => \N__8060\,
            in3 => \N__8389\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13030\,
            ce => \N__8002\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNINQKO8_0_0_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__9801\,
            in1 => \N__9825\,
            in2 => \N__11595\,
            in3 => \N__10232\,
            lcout => \DUT.uart_inst0.N_22_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_1_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111000000010"
        )
    port map (
            in0 => \N__10355\,
            in1 => \N__11548\,
            in2 => \N__8396\,
            in3 => \N__8051\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13030\,
            ce => \N__8002\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_2_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010111000000"
        )
    port map (
            in0 => \N__8387\,
            in1 => \N__8045\,
            in2 => \N__11596\,
            in3 => \N__8099\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13030\,
            ce => \N__8002\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_3_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__8069\,
            in1 => \N__11546\,
            in2 => \N__8039\,
            in3 => \N__8390\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13030\,
            ce => \N__8002\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_4_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010111000000"
        )
    port map (
            in0 => \N__8388\,
            in1 => \N__8030\,
            in2 => \N__11597\,
            in3 => \N__10328\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13030\,
            ce => \N__8002\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_5_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011100010"
        )
    port map (
            in0 => \N__10934\,
            in1 => \N__11547\,
            in2 => \N__8021\,
            in3 => \N__8391\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13030\,
            ce => \N__8002\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_6_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011001010"
        )
    port map (
            in0 => \N__10748\,
            in1 => \N__8012\,
            in2 => \N__11598\,
            in3 => \N__8395\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13030\,
            ce => \N__8002\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_7_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000100010"
        )
    port map (
            in0 => \N__10280\,
            in1 => \N__11576\,
            in2 => \N__8423\,
            in3 => \N__8411\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13025\,
            ce => \N__8003\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_1_5_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__11412\,
            in1 => \_gnd_net_\,
            in2 => \N__11603\,
            in3 => \N__11664\,
            lcout => \DUT.uart_inst0.N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_3_2_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__11665\,
            in1 => \N__11566\,
            in2 => \_gnd_net_\,
            in3 => \N__11413\,
            lcout => \DUT.uart_inst0.N_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNICU6U_1_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111111"
        )
    port map (
            in0 => \N__11410\,
            in1 => \_gnd_net_\,
            in2 => \N__11601\,
            in3 => \N__11662\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_79_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNI5PJS2_1_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101011111"
        )
    port map (
            in0 => \N__12063\,
            in1 => \_gnd_net_\,
            in2 => \N__8126\,
            in3 => \N__12227\,
            lcout => \DUT.uart_inst0.N_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNO_0_0_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101111"
        )
    port map (
            in0 => \N__11411\,
            in1 => \_gnd_net_\,
            in2 => \N__11602\,
            in3 => \N__11663\,
            lcout => \DUT.uart_inst0.tx_state_ns_i_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNI3R8C_1_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__12062\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11409\,
            lcout => \DUT.rTransmitc_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNIBTN81_0_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__11565\,
            in1 => \N__9872\,
            in2 => \_gnd_net_\,
            in3 => \N__11661\,
            lcout => \DUT.uart_inst0.N_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__8090\,
            in1 => \N__10826\,
            in2 => \N__12461\,
            in3 => \N__10903\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__10830\,
            in1 => \N__12095\,
            in2 => \N__8114\,
            in3 => \N__8111\,
            lcout => \DUT.rFifoDatarx_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12499\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13019\,
            ce => \N__13189\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__10904\,
            in1 => \N__12410\,
            in2 => \N__10853\,
            in3 => \N__8456\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__12086\,
            in1 => \N__8084\,
            in2 => \N__8072\,
            in3 => \N__10831\,
            lcout => \DUT.rFifoDatarx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12438\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13019\,
            ce => \N__13189\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_0_RNI86BE_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111011101"
        )
    port map (
            in0 => \N__8449\,
            in1 => \N__10825\,
            in2 => \N__8438\,
            in3 => \N__10902\,
            lcout => \DUT.rFifoDataror_1\,
            ltout => \DUT.rFifoDataror_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_0_RNIKCMS_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8414\,
            in3 => \N__8407\,
            lcout => \DUT.rFifoDataror_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.rTransmit_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__8492\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11605\,
            lcout => \DUT.rTransmitZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13014\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rReadPtr_1_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__8246\,
            in1 => \_gnd_net_\,
            in2 => \N__9003\,
            in3 => \N__8237\,
            lcout => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13014\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rReadPtr_1_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100100001100"
        )
    port map (
            in0 => \N__10598\,
            in1 => \N__10851\,
            in2 => \N__9038\,
            in3 => \N__10915\,
            lcout => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13014\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rReadPtr_0_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__10914\,
            in1 => \N__9034\,
            in2 => \_gnd_net_\,
            in3 => \N__10597\,
            lcout => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13014\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rReadPtr_RNI4NC92_1_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__8332\,
            in1 => \N__8964\,
            in2 => \_gnd_net_\,
            in3 => \N__8245\,
            lcout => \DUT.fifo_rx_inst.un1_i11_2_i\,
            ltout => \DUT.fifo_rx_inst.un1_i11_2_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rReadPtr_0_LC_10_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000110"
        )
    port map (
            in0 => \N__8176\,
            in1 => \N__10654\,
            in2 => \N__8231\,
            in3 => \N__8227\,
            lcout => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13014\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_RNIN79A_0_1_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__8576\,
            in1 => \N__8532\,
            in2 => \_gnd_net_\,
            in3 => \N__8474\,
            lcout => \DUT.fifo_tx_inst.rFifoData_awe1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNI8CH01_1_LC_10_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__11604\,
            in1 => \N__11438\,
            in2 => \N__12074\,
            in3 => \N__11660\,
            lcout => \DUT.uart_inst0.N_65_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__10555\,
            in1 => \N__10658\,
            in2 => \N__10736\,
            in3 => \N__8501\,
            lcout => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNIME2J_0_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010111"
        )
    port map (
            in0 => \N__11636\,
            in1 => \N__10682\,
            in2 => \N__10734\,
            in3 => \N__10553\,
            lcout => \DUT.fifo_tx_inst.N_83\,
            ltout => \DUT.fifo_tx_inst.N_83_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNIDGST_0_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10655\,
            in2 => \N__8504\,
            in3 => \N__11637\,
            lcout => \DUT.fifo_tx_inst.N_88\,
            ltout => \DUT.fifo_tx_inst.N_88_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_0_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100000000111"
        )
    port map (
            in0 => \N__10659\,
            in1 => \N__10557\,
            in2 => \N__8495\,
            in3 => \N__10730\,
            lcout => \DUT.rFifoCount_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13008\,
            ce => 'H',
            sr => \N__10522\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNIBPFM_1_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \N__10684\,
            in1 => \N__10594\,
            in2 => \_gnd_net_\,
            in3 => \N__10657\,
            lcout => \DUT.fifo_tx_inst.rFifoCount_RNIBPFMZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.rTransmit_RNO_0_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101011"
        )
    port map (
            in0 => \N__9830\,
            in1 => \N__10683\,
            in2 => \N__10735\,
            in3 => \N__10556\,
            lcout => \DUT.rTransmitc\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNIMBD3_2_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__10554\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10656\,
            lcout => \DUT.fifo_tx_inst.rWritePtr16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rReadPtr_RNILV421_0_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100110011"
        )
    port map (
            in0 => \N__10595\,
            in1 => \N__12071\,
            in2 => \N__10916\,
            in3 => \N__10850\,
            lcout => \DUT.fifo_tx_inst.un1_i11_2_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rTxByte_esr_1_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__8976\,
            in1 => \N__8909\,
            in2 => \N__8897\,
            in3 => \N__8888\,
            lcout => \rTxByteZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13005\,
            ce => \N__8878\,
            sr => \N__8851\
        );

    \fifo_inst.ft2232h_inst.rFifoState_4_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__8612\,
            in1 => \N__8637\,
            in2 => \_gnd_net_\,
            in3 => \N__8761\,
            lcout => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13047\,
            ce => 'H',
            sr => \N__10528\
        );

    \fifo_inst.ft2232h_inst.rFifoState_0_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__8638\,
            in1 => \N__8815\,
            in2 => \N__8617\,
            in3 => \N__10982\,
            lcout => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13047\,
            ce => 'H',
            sr => \N__10528\
        );

    \fifo_inst.ft2232h_inst.rTx_n_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__8639\,
            in1 => \N__8762\,
            in2 => \N__8618\,
            in3 => \N__8775\,
            lcout => \P1A4_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13047\,
            ce => 'H',
            sr => \N__10528\
        );

    \fifo_inst.ft2232h_inst.rFifoState_3_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__11120\,
            in1 => \N__11066\,
            in2 => \_gnd_net_\,
            in3 => \N__11009\,
            lcout => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13047\,
            ce => 'H',
            sr => \N__10528\
        );

    \fifo_inst.ft2232h_inst.rTxBusReady_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101110000"
        )
    port map (
            in0 => \N__8613\,
            in1 => \N__8635\,
            in2 => \N__8679\,
            in3 => \N__9911\,
            lcout => \rTxBusReady\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13047\,
            ce => 'H',
            sr => \N__10528\
        );

    \fifo_inst.ft2232h_inst.rTxRdEn_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8608\,
            in2 => \_gnd_net_\,
            in3 => \N__8636\,
            lcout => \fifo_inst.ft2232h_inst.rTxRdEnZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13047\,
            ce => 'H',
            sr => \N__10528\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8591\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9227\,
            in2 => \N__12842\,
            in3 => \N__9194\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_0\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9647\,
            in2 => \N__12846\,
            in3 => \N__9191\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_1\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_2_THRU_LUT4_0_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9188\,
            in2 => \N__12843\,
            in3 => \N__9149\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_2\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9490\,
            in2 => \N__12847\,
            in3 => \N__9146\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_3\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_4_THRU_LUT4_0_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9143\,
            in2 => \N__12844\,
            in3 => \N__9122\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_4\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_5_THRU_LUT4_0_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9118\,
            in2 => \N__12848\,
            in3 => \N__9095\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_5\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9091\,
            in2 => \N__12845\,
            in3 => \N__9068\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_6\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9064\,
            in2 => \N__12817\,
            in3 => \N__9041\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_11_14_0_\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9415\,
            in2 => \N__12814\,
            in3 => \N__9389\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_8\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_LUT4_0_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9385\,
            in2 => \N__12818\,
            in3 => \N__9362\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_9\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_LUT4_0_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9358\,
            in2 => \N__12811\,
            in3 => \N__9335\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_10\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_LUT4_0_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9677\,
            in2 => \N__12815\,
            in3 => \N__9332\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_11\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_LUT4_0_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9329\,
            in2 => \N__12812\,
            in3 => \N__9308\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_12\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_LUT4_0_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9304\,
            in2 => \N__12816\,
            in3 => \N__9281\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_13\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_LUT4_0_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9278\,
            in2 => \N__12813\,
            in3 => \N__9257\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_14\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_LUT4_0_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9253\,
            in2 => \N__12763\,
            in3 => \N__9230\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_17_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__9609\,
            in1 => \N__9697\,
            in2 => \_gnd_net_\,
            in3 => \N__9701\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13036\,
            ce => \N__11979\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_12_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100001000100"
        )
    port map (
            in0 => \N__9683\,
            in1 => \N__9608\,
            in2 => \_gnd_net_\,
            in3 => \N__9675\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13036\,
            ce => \N__11979\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_2_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__9610\,
            in1 => \N__9656\,
            in2 => \_gnd_net_\,
            in3 => \N__9645\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13036\,
            ce => \N__11979\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_4_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100001000100"
        )
    port map (
            in0 => \N__9623\,
            in1 => \N__9611\,
            in2 => \_gnd_net_\,
            in3 => \N__9486\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13036\,
            ce => \N__11979\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_RNO_1_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__11407\,
            in1 => \N__9431\,
            in2 => \N__11600\,
            in3 => \N__10234\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_98_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__9448\,
            in1 => \N__9806\,
            in2 => \N__9464\,
            in3 => \N__10211\,
            lcout => \P1A7_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13031\,
            ce => \N__11985\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_RNO_2_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9873\,
            in2 => \_gnd_net_\,
            in3 => \N__10246\,
            lcout => \DUT.uart_inst0.N_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNISP995_0_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9874\,
            in1 => \N__11150\,
            in2 => \N__11594\,
            in3 => \N__12221\,
            lcout => \DUT.uart_inst0.N_99\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNISP995_0_0_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__12222\,
            in1 => \N__9875\,
            in2 => \N__11599\,
            in3 => \N__11222\,
            lcout => \DUT.uart_inst0.N_100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNIHH651_0_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__10170\,
            in1 => \N__10040\,
            in2 => \_gnd_net_\,
            in3 => \N__9977\,
            lcout => \DUT.uart_inst0.N_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ft2232h_inst.rFifoState_RNIRPB71_0_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__11061\,
            in1 => \N__11108\,
            in2 => \_gnd_net_\,
            in3 => \N__11015\,
            lcout => \fifo_inst.ft2232h_inst.rFifoStatec_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_3_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9843\,
            in1 => \N__9716\,
            in2 => \N__9902\,
            in3 => \N__9769\,
            lcout => \DUT.uart_inst0.N_139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_2_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001001"
        )
    port map (
            in0 => \N__9772\,
            in1 => \N__9844\,
            in2 => \N__9731\,
            in3 => \N__9748\,
            lcout => \DUT.uart_inst0.tx_bits_remainingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13026\,
            ce => 'H',
            sr => \N__10265\
        );

    \DUT.uart_inst0.tx_countdown_RNI3MLP6_1_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__11221\,
            in1 => \N__11149\,
            in2 => \_gnd_net_\,
            in3 => \N__12199\,
            lcout => \DUT.uart_inst0.N_85\,
            ltout => \DUT.uart_inst0.N_85_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNINQKO8_0_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__11541\,
            in1 => \N__9829\,
            in2 => \N__9809\,
            in3 => \N__9802\,
            lcout => \DUT.uart_inst0.N_22\,
            ltout => \DUT.uart_inst0.N_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_0_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9785\,
            in3 => \N__9770\,
            lcout => \DUT.uart_inst0.tx_bits_remainingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13026\,
            ce => 'H',
            sr => \N__10265\
        );

    \DUT.uart_inst0.tx_bits_remaining_1_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010100101"
        )
    port map (
            in0 => \N__9771\,
            in1 => \_gnd_net_\,
            in2 => \N__9730\,
            in3 => \N__9747\,
            lcout => \DUT.uart_inst0.tx_bits_remainingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13026\,
            ce => 'H',
            sr => \N__10265\
        );

    \DUT.uart_inst0.tx_out_RNO_0_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011100100"
        )
    port map (
            in0 => \N__11564\,
            in1 => \N__11406\,
            in2 => \N__10250\,
            in3 => \N__10233\,
            lcout => \DUT.uart_inst0.N_89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11240\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_1_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11252\,
            in2 => \N__12759\,
            in3 => \N__10205\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_1\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_0\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_1\,
            clk => \N__13020\,
            ce => 'H',
            sr => \N__11268\
        );

    \DUT.uart_inst0.tx_clk_divider_2_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12350\,
            in2 => \N__12741\,
            in3 => \N__10202\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_2\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_1\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_2\,
            clk => \N__13020\,
            ce => 'H',
            sr => \N__11268\
        );

    \DUT.uart_inst0.tx_clk_divider_3_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12311\,
            in2 => \N__12760\,
            in3 => \N__10199\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_3\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_2\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_3\,
            clk => \N__13020\,
            ce => 'H',
            sr => \N__11268\
        );

    \DUT.uart_inst0.tx_clk_divider_4_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12338\,
            in2 => \N__12742\,
            in3 => \N__10196\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_4\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_3\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_4\,
            clk => \N__13020\,
            ce => 'H',
            sr => \N__11268\
        );

    \DUT.uart_inst0.tx_clk_divider_5_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12325\,
            in2 => \N__12761\,
            in3 => \N__10193\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_5\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_4\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_5\,
            clk => \N__13020\,
            ce => 'H',
            sr => \N__11268\
        );

    \DUT.uart_inst0.tx_clk_divider_6_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12260\,
            in2 => \N__12743\,
            in3 => \N__10190\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_6\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_5\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_6\,
            clk => \N__13020\,
            ce => 'H',
            sr => \N__11268\
        );

    \DUT.uart_inst0.tx_clk_divider_7_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12287\,
            in2 => \N__12762\,
            in3 => \N__10187\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_7\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_6\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_7\,
            clk => \N__13020\,
            ce => 'H',
            sr => \N__11268\
        );

    \DUT.uart_inst0.tx_clk_divider_8_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11288\,
            in2 => \N__12758\,
            in3 => \N__10310\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_11_19_0_\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_8\,
            clk => \N__13015\,
            ce => 'H',
            sr => \N__11272\
        );

    \DUT.uart_inst0.tx_clk_divider_9_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12702\,
            in2 => \N__11333\,
            in3 => \N__10307\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_9\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_8\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_9\,
            clk => \N__13015\,
            ce => 'H',
            sr => \N__11272\
        );

    \DUT.uart_inst0.tx_clk_divider_10_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11318\,
            in2 => \N__12756\,
            in3 => \N__10304\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_10\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_9\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_10\,
            clk => \N__13015\,
            ce => 'H',
            sr => \N__11272\
        );

    \DUT.uart_inst0.tx_clk_divider_11_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12695\,
            in2 => \N__11306\,
            in3 => \N__10301\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_11\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_10\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_11\,
            clk => \N__13015\,
            ce => 'H',
            sr => \N__11272\
        );

    \DUT.uart_inst0.tx_clk_divider_12_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12299\,
            in2 => \N__12757\,
            in3 => \N__10298\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_12\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_11\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_12\,
            clk => \N__13015\,
            ce => 'H',
            sr => \N__11272\
        );

    \DUT.uart_inst0.tx_clk_divider_13_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12274\,
            in2 => \_gnd_net_\,
            in3 => \N__10295\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13015\,
            ce => 'H',
            sr => \N__11272\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__10907\,
            in1 => \N__13283\,
            in2 => \N__10855\,
            in3 => \N__10271\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__10292\,
            in1 => \N__12533\,
            in2 => \N__10283\,
            in3 => \N__10841\,
            lcout => \DUT.rFifoDatarx_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13320\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13009\,
            ce => \N__13190\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__10376\,
            in1 => \N__10832\,
            in2 => \N__13067\,
            in3 => \N__10905\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__10839\,
            in1 => \N__12107\,
            in2 => \N__10403\,
            in3 => \N__10400\,
            lcout => \DUT.rFifoDatarxZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13098\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13009\,
            ce => \N__13190\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__10906\,
            in1 => \N__12506\,
            in2 => \N__10854\,
            in3 => \N__13235\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__12101\,
            in1 => \N__10370\,
            in2 => \N__10358\,
            in3 => \N__10840\,
            lcout => \DUT.rFifoDatarx_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__10316\,
            in1 => \N__10842\,
            in2 => \N__12368\,
            in3 => \N__10908\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__10847\,
            in1 => \N__12569\,
            in2 => \N__10343\,
            in3 => \N__10340\,
            lcout => \DUT.rFifoDatarx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12390\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13006\,
            ce => \N__13187\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__10909\,
            in1 => \N__13115\,
            in2 => \N__10856\,
            in3 => \N__10922\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_11_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__12557\,
            in1 => \N__10949\,
            in2 => \N__10937\,
            in3 => \N__10848\,
            lcout => \DUT.rFifoDatarx_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13140\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13006\,
            ce => \N__13187\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__13196\,
            in1 => \N__10846\,
            in2 => \N__12359\,
            in3 => \N__10910\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_11_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__10849\,
            in1 => \N__12545\,
            in2 => \N__10763\,
            in3 => \N__10760\,
            lcout => \DUT.rFifoDatarx_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10729\,
            in2 => \N__10703\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_22_0_\,
            carryout => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_1_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10685\,
            in2 => \N__10694\,
            in3 => \N__10667\,
            lcout => \DUT.rFifoCount_1\,
            ltout => OPEN,
            carryin => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0\,
            carryout => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1\,
            clk => \N__13003\,
            ce => 'H',
            sr => \N__10521\
        );

    \DUT.fifo_tx_inst.rFifoCount_2_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001111011100001"
        )
    port map (
            in0 => \N__10664\,
            in1 => \N__10596\,
            in2 => \N__10567\,
            in3 => \N__10574\,
            lcout => \DUT.rFifoCount_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13003\,
            ce => 'H',
            sr => \N__10521\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10496\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13001\,
            ce => \N__10442\,
            sr => \_gnd_net_\
        );

    \fifo_inst.ft2232h_inst.rFifoState_RNO_0_0_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11123\,
            in1 => \N__11065\,
            in2 => \_gnd_net_\,
            in3 => \N__11005\,
            lcout => \fifo_inst.ft2232h_inst.N_101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_7_3_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000100"
        )
    port map (
            in0 => \N__11882\,
            in1 => \N__11719\,
            in2 => \_gnd_net_\,
            in3 => \N__11765\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_4_3_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__11609\,
            in1 => \N__11431\,
            in2 => \N__10976\,
            in3 => \N__11687\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g0_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__12170\,
            in1 => \N__11879\,
            in2 => \N__10973\,
            in3 => \N__12223\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g0_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_3_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100000101"
        )
    port map (
            in0 => \N__10958\,
            in1 => \N__10970\,
            in2 => \N__10961\,
            in3 => \N__12116\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13029\,
            ce => \N__11975\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_2_3_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__11880\,
            in1 => \N__11724\,
            in2 => \_gnd_net_\,
            in3 => \N__11768\,
            lcout => \DUT.uart_inst0.g0_i_a6_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_0_4_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__11767\,
            in1 => \N__11881\,
            in2 => \N__11728\,
            in3 => \N__12169\,
            lcout => \DUT.uart_inst0.g0_i_o2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_2_5_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11878\,
            in2 => \_gnd_net_\,
            in3 => \N__11766\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g0_i_o2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_0_5_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__11723\,
            in1 => \N__11919\,
            in2 => \N__10952\,
            in3 => \N__12168\,
            lcout => \DUT.uart_inst0.g0_i_o2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNI67HK1_5_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__11910\,
            in1 => \N__11868\,
            in2 => \N__11829\,
            in3 => \N__11717\,
            lcout => \DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0\,
            ltout => \DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNIJKPE2_1_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11764\,
            in2 => \N__11225\,
            in3 => \N__12154\,
            lcout => \DUT.uart_inst0.N_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_4_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000010010"
        )
    port map (
            in0 => \N__12225\,
            in1 => \N__11342\,
            in2 => \N__11920\,
            in3 => \N__11210\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13024\,
            ce => \N__11977\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_5_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100100001100"
        )
    port map (
            in0 => \N__11204\,
            in1 => \N__11821\,
            in2 => \N__11198\,
            in3 => \N__12226\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13024\,
            ce => \N__11977\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_2_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110111110101"
        )
    port map (
            in0 => \N__11693\,
            in1 => \N__11183\,
            in2 => \N__11171\,
            in3 => \N__11786\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13024\,
            ce => \N__11977\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNIUUGK1_2_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__11718\,
            in1 => \N__11763\,
            in2 => \N__11883\,
            in3 => \N__12153\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_state_ns_i_i_o2_a0_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNIJKPE2_5_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__11911\,
            in1 => \_gnd_net_\,
            in2 => \N__11153\,
            in3 => \N__11822\,
            lcout => \DUT.uart_inst0.N_71_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_1_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100100001010"
        )
    port map (
            in0 => \N__11773\,
            in1 => \N__12155\,
            in2 => \N__11138\,
            in3 => \N__12224\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13024\,
            ce => \N__11977\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_0_0_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__11608\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11684\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g0_i_a3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_0_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011000000110"
        )
    port map (
            in0 => \N__12217\,
            in1 => \N__12167\,
            in2 => \N__12077\,
            in3 => \N__11433\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13018\,
            ce => \N__11981\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_5_2_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__11918\,
            in1 => \N__11884\,
            in2 => \N__11833\,
            in3 => \N__12156\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g0_11_a3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_2_2_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010110001"
        )
    port map (
            in0 => \N__12216\,
            in1 => \N__11795\,
            in2 => \N__11789\,
            in3 => \N__12166\,
            lcout => \DUT.uart_inst0.N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_1_2_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111000001111"
        )
    port map (
            in0 => \N__11772\,
            in1 => \N__12157\,
            in2 => \N__11729\,
            in3 => \N__12215\,
            lcout => \DUT.uart_inst0.N_6_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_1_4_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__11685\,
            in1 => \N__11607\,
            in2 => \_gnd_net_\,
            in3 => \N__11432\,
            lcout => \DUT.uart_inst0.N_11_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_8_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11329\,
            in1 => \N__11317\,
            in2 => \N__11305\,
            in3 => \N__11287\,
            lcout => \DUT.uart_inst0.un1_tx_clk_divider_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_0_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__11239\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12636\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13013\,
            ce => 'H',
            sr => \N__11276\
        );

    \DUT.uart_inst0.tx_clk_divider_RNIBPK2_0_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11251\,
            in2 => \_gnd_net_\,
            in3 => \N__11238\,
            lcout => \DUT.uart_inst0.un1_tx_clk_divider_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_RNI2V95_2_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12349\,
            in1 => \N__12337\,
            in2 => \N__12326\,
            in3 => \N__12310\,
            lcout => \DUT.uart_inst0.un1_tx_clk_divider_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_13_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12298\,
            in1 => \N__12286\,
            in2 => \N__12275\,
            in3 => \N__12259\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.un1_tx_clk_divider_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_RNITC2S1_0_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12248\,
            in1 => \N__12242\,
            in2 => \N__12236\,
            in3 => \N__12233\,
            lcout => \DUT.uart_inst0.un1_tx_clk_divider_0\,
            ltout => \DUT.uart_inst0.un1_tx_clk_divider_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_3_3_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__12158\,
            in1 => \_gnd_net_\,
            in2 => \N__12119\,
            in3 => \_gnd_net_\,
            lcout => \DUT.uart_inst0.N_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13106\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13007\,
            ce => \N__12527\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13276\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13007\,
            ce => \N__12527\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12500\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13007\,
            ce => \N__12527\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12446\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13007\,
            ce => \N__12527\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12398\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13007\,
            ce => \N__12527\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13148\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13007\,
            ce => \N__12527\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13229\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13007\,
            ce => \N__12527\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13322\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13007\,
            ce => \N__12527\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13275\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13004\,
            ce => \N__12879\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12498\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13004\,
            ce => \N__12879\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12445\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13004\,
            ce => \N__12879\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12397\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13004\,
            ce => \N__12879\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13228\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13004\,
            ce => \N__12879\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13321\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13004\,
            ce => \N__12879\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_12_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13274\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13002\,
            ce => \N__13188\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13216\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13002\,
            ce => \N__13188\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13147\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13000\,
            ce => \N__12884\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13105\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13010\,
            ce => \N__12883\,
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
