-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Mar 30 2020 12:32:26

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    ioFifoData : out std_logic_vector(7 downto 0);
    P1A9 : out std_logic;
    P1A1 : in std_logic;
    P1A8 : out std_logic;
    oRx_n : out std_logic;
    P1A7 : out std_logic;
    P1A3 : out std_logic;
    iTxE_n : in std_logic;
    iRxF_n : in std_logic;
    iClk : in std_logic;
    P1A2 : out std_logic;
    BTN_N : in std_logic;
    BTN1 : in std_logic;
    oTx_n : out std_logic;
    P1A4 : out std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__14220\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14205\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14196\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14187\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14169\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14160\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14151\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14142\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14134\ : std_logic;
signal \N__14133\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14123\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14106\ : std_logic;
signal \N__14105\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14097\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14079\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14069\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14061\ : std_logic;
signal \N__14060\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14052\ : std_logic;
signal \N__14051\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14043\ : std_logic;
signal \N__14042\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14034\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14016\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__14012\ : std_logic;
signal \N__14009\ : std_logic;
signal \N__14006\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14004\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13982\ : std_logic;
signal \N__13979\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13971\ : std_logic;
signal \N__13968\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13962\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13926\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13920\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13914\ : std_logic;
signal \N__13913\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13911\ : std_logic;
signal \N__13908\ : std_logic;
signal \N__13907\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13899\ : std_logic;
signal \N__13898\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13892\ : std_logic;
signal \N__13887\ : std_logic;
signal \N__13884\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13872\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13870\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13863\ : std_logic;
signal \N__13860\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13854\ : std_logic;
signal \N__13853\ : std_logic;
signal \N__13850\ : std_logic;
signal \N__13847\ : std_logic;
signal \N__13844\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13838\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13829\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13826\ : std_logic;
signal \N__13823\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13817\ : std_logic;
signal \N__13814\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13805\ : std_logic;
signal \N__13796\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13769\ : std_logic;
signal \N__13766\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13763\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13746\ : std_logic;
signal \N__13743\ : std_logic;
signal \N__13740\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13730\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13724\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13667\ : std_logic;
signal \N__13664\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13657\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13653\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13617\ : std_logic;
signal \N__13614\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13610\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13598\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13587\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13578\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13573\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13567\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13552\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13518\ : std_logic;
signal \N__13515\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13498\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13495\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13491\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13489\ : std_logic;
signal \N__13488\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13483\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13481\ : std_logic;
signal \N__13480\ : std_logic;
signal \N__13479\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13476\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13473\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13471\ : std_logic;
signal \N__13470\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13464\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13462\ : std_logic;
signal \N__13461\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13459\ : std_logic;
signal \N__13458\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13453\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13446\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13444\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13441\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13438\ : std_logic;
signal \N__13437\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13435\ : std_logic;
signal \N__13434\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13292\ : std_logic;
signal \N__13291\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13285\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13282\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13245\ : std_logic;
signal \N__13242\ : std_logic;
signal \N__13239\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13191\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13146\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13138\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13083\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13022\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12959\ : std_logic;
signal \N__12956\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12939\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12922\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12886\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12877\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12847\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12838\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12820\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12768\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12757\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12748\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12730\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12724\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12721\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12714\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12710\ : std_logic;
signal \N__12707\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12585\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12388\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12382\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12326\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12293\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12254\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12219\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12211\ : std_logic;
signal \N__12208\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12189\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12182\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12176\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10629\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10434\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10380\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10177\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8829\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7902\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7893\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7551\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7499\ : std_logic;
signal \N__7496\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7350\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7212\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6432\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6315\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6312\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6231\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5364\ : std_logic;
signal \N__5361\ : std_logic;
signal \BTN_N_c\ : std_logic;
signal \wTxRdData_3\ : std_logic;
signal \wTxRdData_5\ : std_logic;
signal \wTxRdData_2\ : std_logic;
signal \wTxRdData_6\ : std_logic;
signal \wTxRdData_7\ : std_logic;
signal \wTxRdData_0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \wTxRdData_4\ : std_logic;
signal \wTxRdData_1\ : std_logic;
signal \GNDG0\ : std_logic;
signal \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_3_cascade_\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_11\ : std_logic;
signal \bfn_10_16_0_\ : std_logic;
signal \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0\ : std_logic;
signal \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_awe3_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.un1_i11_i_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.un1_i11_i\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_0\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_1\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_3\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_2\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_3\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_4\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_5\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_7\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_6\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_7\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_8\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO\ : std_logic;
signal \bfn_11_12_0_\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_9\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_8\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_10\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_9\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_11\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_10\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_12\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_11\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_12\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_13\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_14\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_15\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_16\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.recv_state_ns_0_0_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_50\ : std_logic;
signal \DUT.uart_inst0.recv_state_srsts_1_3_cascade_\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_3\ : std_logic;
signal \DUT.fifo_rx_inst.N_88_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoCount_RNIK3G92Z0Z_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoCountZ0Z_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1Z0Z_0_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.N_97_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0\ : std_logic;
signal \DUT.fifo_rx_inst.N_97\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoCountZ0Z_0\ : std_logic;
signal \DUT.wRcvd\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoCountZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ1Z_1\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_9_cascade_\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_15_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_17\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_12\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_13\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_14\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_15\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_16\ : std_logic;
signal \DUT.uart_inst0.N_46_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_0\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_RNI8KQG9Z0Z_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_8_i_o2_2_2_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_42_cascade_\ : std_logic;
signal \bfn_12_14_0_\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_0\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_1\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_2\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_3\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_4\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_5\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_6\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_7\ : std_logic;
signal \bfn_12_15_0_\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_8\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_9\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_10\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_11\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_12\ : std_logic;
signal \DUT.uart_inst0.N_12_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_7_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remainingZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.m5_0_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_6_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remainingZ0Z_2\ : std_logic;
signal \DUT.fifo_rx_inst.un1_i11_2_i\ : std_logic;
signal \DUT.fifo_rx_inst.un1_i11_2_i_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.N_88\ : std_logic;
signal \DUT.fifo_rx_inst.rWritePtrZ0Z_0\ : std_logic;
signal \DUT.fifo_rx_inst.rWritePtrZ0Z_1\ : std_logic;
signal \DUT.fifo_rx_inst.N_85\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remainingZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.m5_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_6_0\ : std_logic;
signal \wPllLocked_i\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_5\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_6\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_6\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_0_c_RNOZ0\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_RNICSMA4Z0Z_1\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_1\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_0\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_1\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ1Z_3\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_RNIEUMA4Z0Z_3\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_2\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_3\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_4\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_5\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_RNIFVMA4Z0Z_4\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_15\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_14\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_RNIDTMA4Z0Z_2\ : std_logic;
signal \DUT.uart_inst0.N_47\ : std_logic;
signal \DUT.uart_inst0.N_68\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_2\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_3\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_4\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa_0_a2_0_a2_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_8_i_o2_2_2\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_12\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_7\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_13\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_6\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_8_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_9_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_3_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_11\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_10\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_9\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_8\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_7_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_10_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_1_sqmuxa_1_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_1_sqmuxa_1_i\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.g0_0_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remainingZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.N_62_4\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.recv_state_srsts_1_2_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_42\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.m5_0_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDataro_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDataro_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_6\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remaining_RNI5UON8Z0Z_3_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_109_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIKK41CZ0_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_109\ : std_logic;
signal \DUT.uart_inst0.tx_state_ns_i_i_a3_1_0\ : std_logic;
signal \DUT.uart_inst0.N_82\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_3_cry_0_c_RNOZ0\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_3\ : std_logic;
signal \bfn_14_14_0_\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_3_cry_0\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_RNI5L692Z0Z_2\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_3_cry_1\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_3_cry_2\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_RNI7N692Z0Z_4\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_3_cry_3\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_3_axb_5\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_3_cry_4\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_RNI4K692Z0Z_1\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_10\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ1Z_3\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_8\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_9\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_RNI6M692Z0Z_3\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \DUT.uart_inst0.un1_tx_bits_remaining_cry_0\ : std_logic;
signal \DUT.uart_inst0.un1_tx_bits_remaining_cry_1\ : std_logic;
signal \DUT.uart_inst0.un1_tx_bits_remaining_cry_2\ : std_logic;
signal \P1A3_c\ : std_logic;
signal \N_100_i\ : std_logic;
signal \DUT.fifo_rx_inst.rTxByte_52_1\ : std_logic;
signal \DUT.fifo_rx_inst.rTxByte_52_0_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1Z0Z_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_6\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_awe1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_5\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_5\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_6\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_5\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \P1A1_c\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_4\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_3\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_3_cascade_\ : std_logic;
signal \P1A7_c\ : std_logic;
signal \DUT.uart_inst0.N_112\ : std_logic;
signal \DUT.uart_inst0.tx_out_6_iv_0_a3_1_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_out_6_iv_0_a3_1_sx_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_113\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_7_i_a3_0_sx_3_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_116\ : std_logic;
signal \DUT.uart_inst0.N_76_i\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_3_2\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_3_4\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_3_1\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_3_3\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_3_0\ : std_logic;
signal \DUT.uart_inst0.N_77_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_3_5\ : std_logic;
signal \DUT.uart_inst0.tx_state_RNI9DTT5Z0Z_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIMJ5ECZ0\ : std_logic;
signal \DUT.uart_inst0.N_99_cascade_\ : std_logic;
signal \DUT.uart_inst0.un1_tx_bits_remaining_cry_0_c_RNOZ0\ : std_logic;
signal \DUT.tx_state_1\ : std_logic;
signal \DUT.uart_inst0.N_77\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remaining_RNO_0Z0Z_3\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remaining_RNIAIE4LZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remainingZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remainingZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.N_124\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remainingZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remaining_RNIBJE4LZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remainingZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.N_96\ : std_logic;
signal \DUT.uart_inst0.N_99\ : std_logic;
signal \DUT.uart_inst0.un1_tx_bits_remaining_axb_3\ : std_logic;
signal \P1A4_c\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDataro_3\ : std_logic;
signal \fifo_inst.ft2232h_inst.rFifoStateZ0Z_1\ : std_logic;
signal \fifo_inst.ft2232h_inst.N_103\ : std_logic;
signal \fifo_inst.ft2232h_inst.rFifoStateZ0Z_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDataro_2\ : std_logic;
signal \fifo_inst.ft2232h_inst.rFifoStateZ0Z_0\ : std_logic;
signal \iTxE_n_c\ : std_logic;
signal \iRxF_n_c\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_0\ : std_logic;
signal \DUT.fifo_rx_inst.rReadPtrZ0Z_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1\ : std_logic;
signal \DUT.fifo_rx_inst.rReadPtrZ0Z_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2\ : std_logic;
signal \N_100_i_0\ : std_logic;
signal \rFifoDatarff_0_RNIHJV05\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_awe3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_0\ : std_logic;
signal \DUT.wRxByte_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_1\ : std_logic;
signal \DUT.wRxByte_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_2\ : std_logic;
signal \DUT.wRxByte_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_3\ : std_logic;
signal \DUT.wRxByte_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_4\ : std_logic;
signal \DUT.wRxByte_5\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_5\ : std_logic;
signal \DUT.wRxByte_6\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_6\ : std_logic;
signal \DUT.wRxByte_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_awe2\ : std_logic;
signal \DUT.wRxByte_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_awe0\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddr_0_2\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_1_1_cascade_\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIZ0Z_1\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddr_0_1\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIZ0Z_1_cascade_\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_1\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_7\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_6\ : std_logic;
signal \DUT.tx_state_0\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.N_71_i\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_\ : std_logic;
signal \DUT.rFifoDatarx_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_\ : std_logic;
signal \DUT.rFifoDatarx_6\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_6\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_6\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_4\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddr_0_7\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddr_0_4\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddr_0_6\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_1_1\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_2\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1_c_RNI5GZ0Z02\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_4\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_3_c_RNI7KZ0Z22\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_3\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_4\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_5_c_RNI9OZ0Z42\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_5\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_6_c_RNIAQZ0Z52\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_6\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_7\ : std_logic;
signal \fifo_inst.ft2232h_inst.rFifoState_RNIG8PKZ0Z_4\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_7\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_6\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un15_rRamRdAddr_5\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un15_rRamRdAddr_cascade_\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddr_0_0\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddr_rst_cascade_\ : std_logic;
signal \bfn_17_12_0_\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_3\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIJ4MZ0Z4\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_4\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_7\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_7\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_8\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_3\ : std_logic;
signal \DUT.rFifoDatarx_3\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_7\ : std_logic;
signal \DUT.rFifoDatarx_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_5\ : std_logic;
signal \DUT.rFifoDatarx_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1_cascade_\ : std_logic;
signal \DUT.rFifoDatarx_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoDataro_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoDataror_1_0_cascade_\ : std_logic;
signal \DUT.rFifoDataror_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_0\ : std_logic;
signal \DUT.rFifoDatarxZ0Z_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_3\ : std_logic;
signal \rTxByteZ0Z_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_6\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoDataro_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_awe2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_awe2_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoDataro_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_awe3_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.un1_i11_i\ : std_logic;
signal \DUT.fifo_tx_inst.un1_i11_i_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rWritePtrZ0Z_1\ : std_logic;
signal \DUT.fifo_tx_inst.rWritePtrZ0Z_0\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddr_rst_7\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddr_0_8\ : std_logic;
signal \fifo_inst.rTxRdEn_RNIS0VN\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddr_rst_4\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddr_0_5\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_5\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un18_rRamWrAddr_4\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un18_rRamWrAddr\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_2\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI6IZ0Z12\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddr_0_3\ : std_logic;
signal \fifo_inst.rTxRdEn_fast\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI20CZ0Z4_cascade_\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un15_rRamRdAddr\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_3\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_0\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_3_cascade_\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_8\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un15_rRamRdAddr_4\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNII2LZ0Z4\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_6\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNIJQZ0Z47\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_7\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIK6NZ0Z4\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_4\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_5\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_2\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_4_cascade_\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un18_rRamWrAddr_5\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_1\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_1_cascade_\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_0\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIZ0\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIZ0_cascade_\ : std_logic;
signal \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7\ : std_logic;
signal \DUT.fifo_tx_inst.N_101_cascade_\ : std_logic;
signal \wPllLocked\ : std_logic;
signal \DUT.fifo_tx_inst.un1_i11_2_i_cascade_\ : std_logic;
signal \wPllLocked_g\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNIIOZ0Z37\ : std_logic;
signal \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_6\ : std_logic;
signal \DUT.fifo_tx_inst.N_101\ : std_logic;
signal \DUT.fifo_tx_inst.un1_i11_2_i\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0\ : std_logic;
signal \rTxByteZ0Z_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_0\ : std_logic;
signal \rTxByteZ0Z_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_1\ : std_logic;
signal \DUT.fifo_tx_inst.rReadPtrZ0Z_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rReadPtrZ0Z_1\ : std_logic;
signal \DUT.rFifoDatarx_2\ : std_logic;
signal \rTxByteZ0Z_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_2\ : std_logic;
signal \rTxByteZ0Z_6\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_6\ : std_logic;
signal \rTxByteZ0Z_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_7\ : std_logic;
signal \rTxByteZ0Z_3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_3\ : std_logic;
signal \DUT.fifo_tx_inst.N_105\ : std_logic;
signal \DUT.N_93_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.N_98_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.N_86\ : std_logic;
signal \DUT.N_93\ : std_logic;
signal \DUT.rTransmitZ0\ : std_logic;
signal \rRxReadZ0\ : std_logic;
signal \DUT.fifo_tx_inst.N_98\ : std_logic;
signal \fifo_inst.ft2232h_inst.rFifoStateZ0Z_3\ : std_logic;
signal \rTxByteZ0Z_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_awe1\ : std_logic;
signal \fifo_inst.ft2232h_inst.rFifoStatec_0\ : std_logic;
signal \fifo_inst.ft2232h_inst.rFifoStateZ0Z_4\ : std_logic;
signal \fifo_inst.wTxRdEn\ : std_logic;
signal \rTxBusReady\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoCountZ0Z_0\ : std_logic;
signal \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0\ : std_logic;
signal \bfn_20_17_0_\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoCount_RNIBPFMZ0Z_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoCountZ0Z_1\ : std_logic;
signal \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0\ : std_logic;
signal \DUT.fifo_tx_inst.un1_rFifoCount_1_axb_2\ : std_logic;
signal \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoCountZ0Z_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_awe3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoDataro_3\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_48mhz_0 : std_logic;
signal \wPllLocked_i_g\ : std_logic;

signal \iClk_wire\ : std_logic;
signal \P1A8_wire\ : std_logic;
signal \ioFifoData_wire\ : std_logic_vector(7 downto 0);
signal \P1A2_wire\ : std_logic;
signal \P1A4_wire\ : std_logic;
signal \oRx_n_wire\ : std_logic;
signal \iRxF_n_wire\ : std_logic;
signal \P1A3_wire\ : std_logic;
signal \P1A7_wire\ : std_logic;
signal \BTN_N_wire\ : std_logic;
signal \oTx_n_wire\ : std_logic;
signal \iTxE_n_wire\ : std_logic;
signal \P1A1_wire\ : std_logic;
signal \P1A9_wire\ : std_logic;
signal \fifo_inst.tx_fifo_inst.ram512x8_inst_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \fifo_inst.tx_fifo_inst.ram512x8_inst_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \fifo_inst.tx_fifo_inst.ram512x8_inst_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \fifo_inst.tx_fifo_inst.ram512x8_inst_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \fifo_inst.tx_fifo_inst.ram512x8_inst_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \top_pll_inst.top_pll_inst_pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \iClk_wire\ <= iClk;
    P1A8 <= \P1A8_wire\;
    ioFifoData <= \ioFifoData_wire\;
    P1A2 <= \P1A2_wire\;
    P1A4 <= \P1A4_wire\;
    oRx_n <= \oRx_n_wire\;
    \iRxF_n_wire\ <= iRxF_n;
    P1A3 <= \P1A3_wire\;
    P1A7 <= \P1A7_wire\;
    \BTN_N_wire\ <= BTN_N;
    oTx_n <= \oTx_n_wire\;
    \iTxE_n_wire\ <= iTxE_n;
    \P1A1_wire\ <= P1A1;
    P1A9 <= \P1A9_wire\;
    \wTxRdData_7\ <= \fifo_inst.tx_fifo_inst.ram512x8_inst_physical_RDATA_wire\(14);
    \wTxRdData_6\ <= \fifo_inst.tx_fifo_inst.ram512x8_inst_physical_RDATA_wire\(12);
    \wTxRdData_5\ <= \fifo_inst.tx_fifo_inst.ram512x8_inst_physical_RDATA_wire\(10);
    \wTxRdData_4\ <= \fifo_inst.tx_fifo_inst.ram512x8_inst_physical_RDATA_wire\(8);
    \wTxRdData_3\ <= \fifo_inst.tx_fifo_inst.ram512x8_inst_physical_RDATA_wire\(6);
    \wTxRdData_2\ <= \fifo_inst.tx_fifo_inst.ram512x8_inst_physical_RDATA_wire\(4);
    \wTxRdData_1\ <= \fifo_inst.tx_fifo_inst.ram512x8_inst_physical_RDATA_wire\(2);
    \wTxRdData_0\ <= \fifo_inst.tx_fifo_inst.ram512x8_inst_physical_RDATA_wire\(0);
    \fifo_inst.tx_fifo_inst.ram512x8_inst_physical_RADDR_wire\ <= '0'&'0'&\N__11445\&\N__10890\&\N__10857\&\N__11667\&\N__10728\&\N__11520\&\N__10773\&\N__10335\&\N__11499\;
    \fifo_inst.tx_fifo_inst.ram512x8_inst_physical_WADDR_wire\ <= '0'&'0'&\N__10965\&\N__11871\&\N__11403\&\N__11829\&\N__11841\&\N__8658\&\N__11799\&\N__11709\&\N__11760\;
    \fifo_inst.tx_fifo_inst.ram512x8_inst_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \fifo_inst.tx_fifo_inst.ram512x8_inst_physical_WDATA_wire\ <= '0'&'0'&'0'&\N__8388\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__12167\;
    \top_pll_inst.top_pll_inst_pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \fifo_inst.tx_fifo_inst.ram512x8_inst_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \fifo_inst.tx_fifo_inst.ram512x8_inst_physical_RDATA_wire\,
            RADDR => \fifo_inst.tx_fifo_inst.ram512x8_inst_physical_RADDR_wire\,
            WADDR => \fifo_inst.tx_fifo_inst.ram512x8_inst_physical_WADDR_wire\,
            MASK => \fifo_inst.tx_fifo_inst.ram512x8_inst_physical_MASK_wire\,
            WDATA => \fifo_inst.tx_fifo_inst.ram512x8_inst_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__13500\,
            RE => \N__13853\,
            WCLKE => 'H',
            WCLK => \N__13499\,
            WE => \N__12168\
        );

    \top_pll_inst.top_pll_inst_pll\ : PLL40
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "0111111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            PLLOUTGLOBAL => clk_48mhz_0,
            SDI => \GNDG0\,
            BYPASS => \GNDG0\,
            RESETB => \N__5433\,
            PLLOUTCORE => OPEN,
            LOCK => \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO\,
            SDO => OPEN,
            SCLK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            EXTFEEDBACK => \GNDG0\,
            DYNAMICDELAY => \top_pll_inst.top_pll_inst_pll_DYNAMICDELAY_wire\,
            PLLIN => \N__14220\
        );

    \top_pll_inst.top_pll_inst_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \VCCG0\,
            DIN => '0',
            DOUT => \N__14220\,
            PACKAGEPIN => \iClk_wire\
        );

    \P1A8_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14206\,
            DIN => \N__14205\,
            DOUT => \N__14204\,
            PACKAGEPIN => \P1A8_wire\
        );

    \P1A8_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__14206\,
            PADOUT => \N__14205\,
            PADIN => \N__14204\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14197\,
            DIN => \N__14196\,
            DOUT => \N__14195\,
            PACKAGEPIN => \ioFifoData_wire\(1)
        );

    \ioFifoData_obuft_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__14197\,
            PADOUT => \N__14196\,
            PADIN => \N__14195\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__13765\,
            DIN0 => OPEN,
            DOUT0 => \N__5502\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14188\,
            DIN => \N__14187\,
            DOUT => \N__14186\,
            PACKAGEPIN => \ioFifoData_wire\(4)
        );

    \ioFifoData_obuft_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__14188\,
            PADOUT => \N__14187\,
            PADIN => \N__14186\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__13749\,
            DIN0 => OPEN,
            DOUT0 => \N__5514\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A2_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14179\,
            DIN => \N__14178\,
            DOUT => \N__14177\,
            PACKAGEPIN => \P1A2_wire\
        );

    \P1A2_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__14179\,
            PADOUT => \N__14178\,
            PADIN => \N__14177\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A4_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14170\,
            DIN => \N__14169\,
            DOUT => \N__14168\,
            PACKAGEPIN => \P1A4_wire\
        );

    \P1A4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14170\,
            PADOUT => \N__14169\,
            PADIN => \N__14168\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9030\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14161\,
            DIN => \N__14160\,
            DOUT => \N__14159\,
            PACKAGEPIN => \ioFifoData_wire\(0)
        );

    \ioFifoData_obuft_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__14161\,
            PADOUT => \N__14160\,
            PADIN => \N__14159\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__13770\,
            DIN0 => OPEN,
            DOUT0 => \N__5454\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \oRx_n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14152\,
            DIN => \N__14151\,
            DOUT => \N__14150\,
            PACKAGEPIN => \oRx_n_wire\
        );

    \oRx_n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14152\,
            PADOUT => \N__14151\,
            PADIN => \N__14150\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7667\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14143\,
            DIN => \N__14142\,
            DOUT => \N__14141\,
            PACKAGEPIN => \ioFifoData_wire\(7)
        );

    \ioFifoData_obuft_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__14143\,
            PADOUT => \N__14142\,
            PADIN => \N__14141\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__13763\,
            DIN0 => OPEN,
            DOUT0 => \N__5469\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \iRxF_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14134\,
            DIN => \N__14133\,
            DOUT => \N__14132\,
            PACKAGEPIN => \iRxF_n_wire\
        );

    \iRxF_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__14134\,
            PADOUT => \N__14133\,
            PADIN => \N__14132\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \iRxF_n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14125\,
            DIN => \N__14124\,
            DOUT => \N__14123\,
            PACKAGEPIN => \P1A3_wire\
        );

    \P1A3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14125\,
            PADOUT => \N__14124\,
            PADIN => \N__14123\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7674\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A7_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14116\,
            DIN => \N__14115\,
            DOUT => \N__14114\,
            PACKAGEPIN => \P1A7_wire\
        );

    \P1A7_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14116\,
            PADOUT => \N__14115\,
            PADIN => \N__14114\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8640\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BTN_N_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14107\,
            DIN => \N__14106\,
            DOUT => \N__14105\,
            PACKAGEPIN => \BTN_N_wire\
        );

    \BTN_N_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__14107\,
            PADOUT => \N__14106\,
            PADIN => \N__14105\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \BTN_N_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14098\,
            DIN => \N__14097\,
            DOUT => \N__14096\,
            PACKAGEPIN => \ioFifoData_wire\(3)
        );

    \ioFifoData_obuft_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__14098\,
            PADOUT => \N__14097\,
            PADIN => \N__14096\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__13729\,
            DIN0 => OPEN,
            DOUT0 => \N__5418\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14089\,
            DIN => \N__14088\,
            DOUT => \N__14087\,
            PACKAGEPIN => \ioFifoData_wire\(6)
        );

    \ioFifoData_obuft_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__14089\,
            PADOUT => \N__14088\,
            PADIN => \N__14087\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__13762\,
            DIN0 => OPEN,
            DOUT0 => \N__5370\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14080\,
            DIN => \N__14079\,
            DOUT => \N__14078\,
            PACKAGEPIN => \ioFifoData_wire\(5)
        );

    \ioFifoData_obuft_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__14080\,
            PADOUT => \N__14079\,
            PADIN => \N__14078\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__13764\,
            DIN0 => OPEN,
            DOUT0 => \N__5400\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \oTx_n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14071\,
            DIN => \N__14070\,
            DOUT => \N__14069\,
            PACKAGEPIN => \oTx_n_wire\
        );

    \oTx_n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__14071\,
            PADOUT => \N__14070\,
            PADIN => \N__14069\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9029\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \iTxE_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14062\,
            DIN => \N__14061\,
            DOUT => \N__14060\,
            PACKAGEPIN => \iTxE_n_wire\
        );

    \iTxE_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__14062\,
            PADOUT => \N__14061\,
            PADIN => \N__14060\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \iTxE_n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14053\,
            DIN => \N__14052\,
            DOUT => \N__14051\,
            PACKAGEPIN => \ioFifoData_wire\(2)
        );

    \ioFifoData_obuft_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__14053\,
            PADOUT => \N__14052\,
            PADIN => \N__14051\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__13769\,
            DIN0 => OPEN,
            DOUT0 => \N__5388\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14044\,
            DIN => \N__14043\,
            DOUT => \N__14042\,
            PACKAGEPIN => \P1A1_wire\
        );

    \P1A1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__14044\,
            PADOUT => \N__14043\,
            PADIN => \N__14042\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \P1A1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A9_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__14035\,
            DIN => \N__14034\,
            DOUT => \N__14033\,
            PACKAGEPIN => \P1A9_wire\
        );

    \P1A9_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__14035\,
            PADOUT => \N__14034\,
            PADIN => \N__14033\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__3332\ : InMux
    port map (
            O => \N__14016\,
            I => \N__14013\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__14013\,
            I => \N__14009\
        );

    \I__3330\ : InMux
    port map (
            O => \N__14012\,
            I => \N__14006\
        );

    \I__3329\ : Span4Mux_v
    port map (
            O => \N__14009\,
            I => \N__14001\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__14006\,
            I => \N__13998\
        );

    \I__3327\ : InMux
    port map (
            O => \N__14005\,
            I => \N__13995\
        );

    \I__3326\ : InMux
    port map (
            O => \N__14004\,
            I => \N__13992\
        );

    \I__3325\ : Span4Mux_h
    port map (
            O => \N__14001\,
            I => \N__13987\
        );

    \I__3324\ : Span4Mux_v
    port map (
            O => \N__13998\,
            I => \N__13987\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__13995\,
            I => \N__13982\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__13992\,
            I => \N__13982\
        );

    \I__3321\ : Span4Mux_v
    port map (
            O => \N__13987\,
            I => \N__13979\
        );

    \I__3320\ : Span4Mux_h
    port map (
            O => \N__13982\,
            I => \N__13976\
        );

    \I__3319\ : Odrv4
    port map (
            O => \N__13979\,
            I => \rTxByteZ0Z_5\
        );

    \I__3318\ : Odrv4
    port map (
            O => \N__13976\,
            I => \rTxByteZ0Z_5\
        );

    \I__3317\ : InMux
    port map (
            O => \N__13971\,
            I => \N__13968\
        );

    \I__3316\ : LocalMux
    port map (
            O => \N__13968\,
            I => \N__13965\
        );

    \I__3315\ : Odrv4
    port map (
            O => \N__13965\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_5\
        );

    \I__3314\ : CEMux
    port map (
            O => \N__13962\,
            I => \N__13958\
        );

    \I__3313\ : CEMux
    port map (
            O => \N__13961\,
            I => \N__13955\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__13958\,
            I => \N__13949\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__13955\,
            I => \N__13949\
        );

    \I__3310\ : CEMux
    port map (
            O => \N__13954\,
            I => \N__13946\
        );

    \I__3309\ : Span4Mux_h
    port map (
            O => \N__13949\,
            I => \N__13942\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__13946\,
            I => \N__13939\
        );

    \I__3307\ : InMux
    port map (
            O => \N__13945\,
            I => \N__13936\
        );

    \I__3306\ : Odrv4
    port map (
            O => \N__13942\,
            I => \DUT.fifo_tx_inst.rFifoData_awe1\
        );

    \I__3305\ : Odrv4
    port map (
            O => \N__13939\,
            I => \DUT.fifo_tx_inst.rFifoData_awe1\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__13936\,
            I => \DUT.fifo_tx_inst.rFifoData_awe1\
        );

    \I__3303\ : InMux
    port map (
            O => \N__13929\,
            I => \N__13926\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__13926\,
            I => \N__13923\
        );

    \I__3301\ : Odrv12
    port map (
            O => \N__13923\,
            I => \fifo_inst.ft2232h_inst.rFifoStatec_0\
        );

    \I__3300\ : InMux
    port map (
            O => \N__13920\,
            I => \N__13914\
        );

    \I__3299\ : InMux
    port map (
            O => \N__13919\,
            I => \N__13914\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__13914\,
            I => \N__13908\
        );

    \I__3297\ : InMux
    port map (
            O => \N__13913\,
            I => \N__13904\
        );

    \I__3296\ : InMux
    port map (
            O => \N__13912\,
            I => \N__13899\
        );

    \I__3295\ : InMux
    port map (
            O => \N__13911\,
            I => \N__13899\
        );

    \I__3294\ : Span4Mux_v
    port map (
            O => \N__13908\,
            I => \N__13895\
        );

    \I__3293\ : InMux
    port map (
            O => \N__13907\,
            I => \N__13892\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__13904\,
            I => \N__13887\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__13899\,
            I => \N__13887\
        );

    \I__3290\ : InMux
    port map (
            O => \N__13898\,
            I => \N__13884\
        );

    \I__3289\ : Span4Mux_h
    port map (
            O => \N__13895\,
            I => \N__13877\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__13892\,
            I => \N__13877\
        );

    \I__3287\ : Span4Mux_h
    port map (
            O => \N__13887\,
            I => \N__13877\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__13884\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_4\
        );

    \I__3285\ : Odrv4
    port map (
            O => \N__13877\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_4\
        );

    \I__3284\ : CascadeMux
    port map (
            O => \N__13872\,
            I => \N__13867\
        );

    \I__3283\ : CascadeMux
    port map (
            O => \N__13871\,
            I => \N__13864\
        );

    \I__3282\ : CascadeMux
    port map (
            O => \N__13870\,
            I => \N__13860\
        );

    \I__3281\ : InMux
    port map (
            O => \N__13867\,
            I => \N__13855\
        );

    \I__3280\ : InMux
    port map (
            O => \N__13864\,
            I => \N__13855\
        );

    \I__3279\ : InMux
    port map (
            O => \N__13863\,
            I => \N__13850\
        );

    \I__3278\ : InMux
    port map (
            O => \N__13860\,
            I => \N__13847\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__13855\,
            I => \N__13844\
        );

    \I__3276\ : InMux
    port map (
            O => \N__13854\,
            I => \N__13840\
        );

    \I__3275\ : SRMux
    port map (
            O => \N__13853\,
            I => \N__13835\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__13850\,
            I => \N__13830\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__13847\,
            I => \N__13830\
        );

    \I__3272\ : Span4Mux_h
    port map (
            O => \N__13844\,
            I => \N__13823\
        );

    \I__3271\ : InMux
    port map (
            O => \N__13843\,
            I => \N__13820\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__13840\,
            I => \N__13817\
        );

    \I__3269\ : CascadeMux
    port map (
            O => \N__13839\,
            I => \N__13814\
        );

    \I__3268\ : CascadeMux
    port map (
            O => \N__13838\,
            I => \N__13811\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__13835\,
            I => \N__13808\
        );

    \I__3266\ : Span4Mux_v
    port map (
            O => \N__13830\,
            I => \N__13805\
        );

    \I__3265\ : InMux
    port map (
            O => \N__13829\,
            I => \N__13796\
        );

    \I__3264\ : InMux
    port map (
            O => \N__13828\,
            I => \N__13796\
        );

    \I__3263\ : InMux
    port map (
            O => \N__13827\,
            I => \N__13796\
        );

    \I__3262\ : InMux
    port map (
            O => \N__13826\,
            I => \N__13796\
        );

    \I__3261\ : Span4Mux_v
    port map (
            O => \N__13823\,
            I => \N__13791\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__13820\,
            I => \N__13791\
        );

    \I__3259\ : Span4Mux_h
    port map (
            O => \N__13817\,
            I => \N__13788\
        );

    \I__3258\ : InMux
    port map (
            O => \N__13814\,
            I => \N__13783\
        );

    \I__3257\ : InMux
    port map (
            O => \N__13811\,
            I => \N__13783\
        );

    \I__3256\ : Odrv4
    port map (
            O => \N__13808\,
            I => \fifo_inst.wTxRdEn\
        );

    \I__3255\ : Odrv4
    port map (
            O => \N__13805\,
            I => \fifo_inst.wTxRdEn\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__13796\,
            I => \fifo_inst.wTxRdEn\
        );

    \I__3253\ : Odrv4
    port map (
            O => \N__13791\,
            I => \fifo_inst.wTxRdEn\
        );

    \I__3252\ : Odrv4
    port map (
            O => \N__13788\,
            I => \fifo_inst.wTxRdEn\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__13783\,
            I => \fifo_inst.wTxRdEn\
        );

    \I__3250\ : IoInMux
    port map (
            O => \N__13770\,
            I => \N__13766\
        );

    \I__3249\ : IoInMux
    port map (
            O => \N__13769\,
            I => \N__13759\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__13766\,
            I => \N__13756\
        );

    \I__3247\ : IoInMux
    port map (
            O => \N__13765\,
            I => \N__13753\
        );

    \I__3246\ : IoInMux
    port map (
            O => \N__13764\,
            I => \N__13750\
        );

    \I__3245\ : IoInMux
    port map (
            O => \N__13763\,
            I => \N__13746\
        );

    \I__3244\ : IoInMux
    port map (
            O => \N__13762\,
            I => \N__13743\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__13759\,
            I => \N__13740\
        );

    \I__3242\ : IoSpan4Mux
    port map (
            O => \N__13756\,
            I => \N__13733\
        );

    \I__3241\ : LocalMux
    port map (
            O => \N__13753\,
            I => \N__13733\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__13750\,
            I => \N__13733\
        );

    \I__3239\ : IoInMux
    port map (
            O => \N__13749\,
            I => \N__13730\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__13746\,
            I => \N__13724\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__13743\,
            I => \N__13724\
        );

    \I__3236\ : IoSpan4Mux
    port map (
            O => \N__13740\,
            I => \N__13719\
        );

    \I__3235\ : IoSpan4Mux
    port map (
            O => \N__13733\,
            I => \N__13719\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__13730\,
            I => \N__13716\
        );

    \I__3233\ : IoInMux
    port map (
            O => \N__13729\,
            I => \N__13713\
        );

    \I__3232\ : Span4Mux_s3_v
    port map (
            O => \N__13724\,
            I => \N__13710\
        );

    \I__3231\ : Span4Mux_s2_v
    port map (
            O => \N__13719\,
            I => \N__13705\
        );

    \I__3230\ : Span4Mux_s2_v
    port map (
            O => \N__13716\,
            I => \N__13705\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__13713\,
            I => \N__13702\
        );

    \I__3228\ : Span4Mux_v
    port map (
            O => \N__13710\,
            I => \N__13699\
        );

    \I__3227\ : Span4Mux_v
    port map (
            O => \N__13705\,
            I => \N__13696\
        );

    \I__3226\ : Span12Mux_s2_v
    port map (
            O => \N__13702\,
            I => \N__13693\
        );

    \I__3225\ : Span4Mux_v
    port map (
            O => \N__13699\,
            I => \N__13690\
        );

    \I__3224\ : Span4Mux_v
    port map (
            O => \N__13696\,
            I => \N__13687\
        );

    \I__3223\ : Span12Mux_v
    port map (
            O => \N__13693\,
            I => \N__13683\
        );

    \I__3222\ : Span4Mux_v
    port map (
            O => \N__13690\,
            I => \N__13678\
        );

    \I__3221\ : Span4Mux_v
    port map (
            O => \N__13687\,
            I => \N__13678\
        );

    \I__3220\ : InMux
    port map (
            O => \N__13686\,
            I => \N__13675\
        );

    \I__3219\ : Odrv12
    port map (
            O => \N__13683\,
            I => \rTxBusReady\
        );

    \I__3218\ : Odrv4
    port map (
            O => \N__13678\,
            I => \rTxBusReady\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__13675\,
            I => \rTxBusReady\
        );

    \I__3216\ : InMux
    port map (
            O => \N__13668\,
            I => \N__13664\
        );

    \I__3215\ : CascadeMux
    port map (
            O => \N__13667\,
            I => \N__13661\
        );

    \I__3214\ : LocalMux
    port map (
            O => \N__13664\,
            I => \N__13658\
        );

    \I__3213\ : InMux
    port map (
            O => \N__13661\,
            I => \N__13653\
        );

    \I__3212\ : Span4Mux_h
    port map (
            O => \N__13658\,
            I => \N__13650\
        );

    \I__3211\ : InMux
    port map (
            O => \N__13657\,
            I => \N__13645\
        );

    \I__3210\ : InMux
    port map (
            O => \N__13656\,
            I => \N__13645\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__13653\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_0\
        );

    \I__3208\ : Odrv4
    port map (
            O => \N__13650\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_0\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__13645\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_0\
        );

    \I__3206\ : CascadeMux
    port map (
            O => \N__13638\,
            I => \N__13635\
        );

    \I__3205\ : InMux
    port map (
            O => \N__13635\,
            I => \N__13632\
        );

    \I__3204\ : LocalMux
    port map (
            O => \N__13632\,
            I => \N__13629\
        );

    \I__3203\ : Odrv4
    port map (
            O => \N__13629\,
            I => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0\
        );

    \I__3202\ : CascadeMux
    port map (
            O => \N__13626\,
            I => \N__13623\
        );

    \I__3201\ : InMux
    port map (
            O => \N__13623\,
            I => \N__13620\
        );

    \I__3200\ : LocalMux
    port map (
            O => \N__13620\,
            I => \N__13617\
        );

    \I__3199\ : Odrv4
    port map (
            O => \N__13617\,
            I => \DUT.fifo_tx_inst.rFifoCount_RNIBPFMZ0Z_1\
        );

    \I__3198\ : CascadeMux
    port map (
            O => \N__13614\,
            I => \N__13611\
        );

    \I__3197\ : InMux
    port map (
            O => \N__13611\,
            I => \N__13604\
        );

    \I__3196\ : InMux
    port map (
            O => \N__13610\,
            I => \N__13604\
        );

    \I__3195\ : InMux
    port map (
            O => \N__13609\,
            I => \N__13601\
        );

    \I__3194\ : LocalMux
    port map (
            O => \N__13604\,
            I => \N__13598\
        );

    \I__3193\ : LocalMux
    port map (
            O => \N__13601\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_1\
        );

    \I__3192\ : Odrv4
    port map (
            O => \N__13598\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_1\
        );

    \I__3191\ : InMux
    port map (
            O => \N__13593\,
            I => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0\
        );

    \I__3190\ : InMux
    port map (
            O => \N__13590\,
            I => \N__13587\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__13587\,
            I => \N__13584\
        );

    \I__3188\ : Odrv12
    port map (
            O => \N__13584\,
            I => \DUT.fifo_tx_inst.un1_rFifoCount_1_axb_2\
        );

    \I__3187\ : InMux
    port map (
            O => \N__13581\,
            I => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1\
        );

    \I__3186\ : InMux
    port map (
            O => \N__13578\,
            I => \N__13574\
        );

    \I__3185\ : CascadeMux
    port map (
            O => \N__13577\,
            I => \N__13570\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__13574\,
            I => \N__13564\
        );

    \I__3183\ : InMux
    port map (
            O => \N__13573\,
            I => \N__13561\
        );

    \I__3182\ : InMux
    port map (
            O => \N__13570\,
            I => \N__13552\
        );

    \I__3181\ : InMux
    port map (
            O => \N__13569\,
            I => \N__13552\
        );

    \I__3180\ : InMux
    port map (
            O => \N__13568\,
            I => \N__13552\
        );

    \I__3179\ : InMux
    port map (
            O => \N__13567\,
            I => \N__13552\
        );

    \I__3178\ : Span4Mux_h
    port map (
            O => \N__13564\,
            I => \N__13549\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__13561\,
            I => \N__13544\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__13552\,
            I => \N__13544\
        );

    \I__3175\ : Odrv4
    port map (
            O => \N__13549\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_2\
        );

    \I__3174\ : Odrv4
    port map (
            O => \N__13544\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_2\
        );

    \I__3173\ : InMux
    port map (
            O => \N__13539\,
            I => \N__13535\
        );

    \I__3172\ : CEMux
    port map (
            O => \N__13538\,
            I => \N__13532\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__13535\,
            I => \N__13529\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__13532\,
            I => \N__13526\
        );

    \I__3169\ : Span4Mux_h
    port map (
            O => \N__13529\,
            I => \N__13523\
        );

    \I__3168\ : Odrv4
    port map (
            O => \N__13526\,
            I => \DUT.fifo_tx_inst.rFifoData_awe3\
        );

    \I__3167\ : Odrv4
    port map (
            O => \N__13523\,
            I => \DUT.fifo_tx_inst.rFifoData_awe3\
        );

    \I__3166\ : InMux
    port map (
            O => \N__13518\,
            I => \N__13515\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__13515\,
            I => \N__13511\
        );

    \I__3164\ : InMux
    port map (
            O => \N__13514\,
            I => \N__13508\
        );

    \I__3163\ : Span4Mux_h
    port map (
            O => \N__13511\,
            I => \N__13505\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__13508\,
            I => \DUT.fifo_tx_inst.rFifoDataro_3\
        );

    \I__3161\ : Odrv4
    port map (
            O => \N__13505\,
            I => \DUT.fifo_tx_inst.rFifoDataro_3\
        );

    \I__3160\ : ClkMux
    port map (
            O => \N__13500\,
            I => \N__13296\
        );

    \I__3159\ : ClkMux
    port map (
            O => \N__13499\,
            I => \N__13296\
        );

    \I__3158\ : ClkMux
    port map (
            O => \N__13498\,
            I => \N__13296\
        );

    \I__3157\ : ClkMux
    port map (
            O => \N__13497\,
            I => \N__13296\
        );

    \I__3156\ : ClkMux
    port map (
            O => \N__13496\,
            I => \N__13296\
        );

    \I__3155\ : ClkMux
    port map (
            O => \N__13495\,
            I => \N__13296\
        );

    \I__3154\ : ClkMux
    port map (
            O => \N__13494\,
            I => \N__13296\
        );

    \I__3153\ : ClkMux
    port map (
            O => \N__13493\,
            I => \N__13296\
        );

    \I__3152\ : ClkMux
    port map (
            O => \N__13492\,
            I => \N__13296\
        );

    \I__3151\ : ClkMux
    port map (
            O => \N__13491\,
            I => \N__13296\
        );

    \I__3150\ : ClkMux
    port map (
            O => \N__13490\,
            I => \N__13296\
        );

    \I__3149\ : ClkMux
    port map (
            O => \N__13489\,
            I => \N__13296\
        );

    \I__3148\ : ClkMux
    port map (
            O => \N__13488\,
            I => \N__13296\
        );

    \I__3147\ : ClkMux
    port map (
            O => \N__13487\,
            I => \N__13296\
        );

    \I__3146\ : ClkMux
    port map (
            O => \N__13486\,
            I => \N__13296\
        );

    \I__3145\ : ClkMux
    port map (
            O => \N__13485\,
            I => \N__13296\
        );

    \I__3144\ : ClkMux
    port map (
            O => \N__13484\,
            I => \N__13296\
        );

    \I__3143\ : ClkMux
    port map (
            O => \N__13483\,
            I => \N__13296\
        );

    \I__3142\ : ClkMux
    port map (
            O => \N__13482\,
            I => \N__13296\
        );

    \I__3141\ : ClkMux
    port map (
            O => \N__13481\,
            I => \N__13296\
        );

    \I__3140\ : ClkMux
    port map (
            O => \N__13480\,
            I => \N__13296\
        );

    \I__3139\ : ClkMux
    port map (
            O => \N__13479\,
            I => \N__13296\
        );

    \I__3138\ : ClkMux
    port map (
            O => \N__13478\,
            I => \N__13296\
        );

    \I__3137\ : ClkMux
    port map (
            O => \N__13477\,
            I => \N__13296\
        );

    \I__3136\ : ClkMux
    port map (
            O => \N__13476\,
            I => \N__13296\
        );

    \I__3135\ : ClkMux
    port map (
            O => \N__13475\,
            I => \N__13296\
        );

    \I__3134\ : ClkMux
    port map (
            O => \N__13474\,
            I => \N__13296\
        );

    \I__3133\ : ClkMux
    port map (
            O => \N__13473\,
            I => \N__13296\
        );

    \I__3132\ : ClkMux
    port map (
            O => \N__13472\,
            I => \N__13296\
        );

    \I__3131\ : ClkMux
    port map (
            O => \N__13471\,
            I => \N__13296\
        );

    \I__3130\ : ClkMux
    port map (
            O => \N__13470\,
            I => \N__13296\
        );

    \I__3129\ : ClkMux
    port map (
            O => \N__13469\,
            I => \N__13296\
        );

    \I__3128\ : ClkMux
    port map (
            O => \N__13468\,
            I => \N__13296\
        );

    \I__3127\ : ClkMux
    port map (
            O => \N__13467\,
            I => \N__13296\
        );

    \I__3126\ : ClkMux
    port map (
            O => \N__13466\,
            I => \N__13296\
        );

    \I__3125\ : ClkMux
    port map (
            O => \N__13465\,
            I => \N__13296\
        );

    \I__3124\ : ClkMux
    port map (
            O => \N__13464\,
            I => \N__13296\
        );

    \I__3123\ : ClkMux
    port map (
            O => \N__13463\,
            I => \N__13296\
        );

    \I__3122\ : ClkMux
    port map (
            O => \N__13462\,
            I => \N__13296\
        );

    \I__3121\ : ClkMux
    port map (
            O => \N__13461\,
            I => \N__13296\
        );

    \I__3120\ : ClkMux
    port map (
            O => \N__13460\,
            I => \N__13296\
        );

    \I__3119\ : ClkMux
    port map (
            O => \N__13459\,
            I => \N__13296\
        );

    \I__3118\ : ClkMux
    port map (
            O => \N__13458\,
            I => \N__13296\
        );

    \I__3117\ : ClkMux
    port map (
            O => \N__13457\,
            I => \N__13296\
        );

    \I__3116\ : ClkMux
    port map (
            O => \N__13456\,
            I => \N__13296\
        );

    \I__3115\ : ClkMux
    port map (
            O => \N__13455\,
            I => \N__13296\
        );

    \I__3114\ : ClkMux
    port map (
            O => \N__13454\,
            I => \N__13296\
        );

    \I__3113\ : ClkMux
    port map (
            O => \N__13453\,
            I => \N__13296\
        );

    \I__3112\ : ClkMux
    port map (
            O => \N__13452\,
            I => \N__13296\
        );

    \I__3111\ : ClkMux
    port map (
            O => \N__13451\,
            I => \N__13296\
        );

    \I__3110\ : ClkMux
    port map (
            O => \N__13450\,
            I => \N__13296\
        );

    \I__3109\ : ClkMux
    port map (
            O => \N__13449\,
            I => \N__13296\
        );

    \I__3108\ : ClkMux
    port map (
            O => \N__13448\,
            I => \N__13296\
        );

    \I__3107\ : ClkMux
    port map (
            O => \N__13447\,
            I => \N__13296\
        );

    \I__3106\ : ClkMux
    port map (
            O => \N__13446\,
            I => \N__13296\
        );

    \I__3105\ : ClkMux
    port map (
            O => \N__13445\,
            I => \N__13296\
        );

    \I__3104\ : ClkMux
    port map (
            O => \N__13444\,
            I => \N__13296\
        );

    \I__3103\ : ClkMux
    port map (
            O => \N__13443\,
            I => \N__13296\
        );

    \I__3102\ : ClkMux
    port map (
            O => \N__13442\,
            I => \N__13296\
        );

    \I__3101\ : ClkMux
    port map (
            O => \N__13441\,
            I => \N__13296\
        );

    \I__3100\ : ClkMux
    port map (
            O => \N__13440\,
            I => \N__13296\
        );

    \I__3099\ : ClkMux
    port map (
            O => \N__13439\,
            I => \N__13296\
        );

    \I__3098\ : ClkMux
    port map (
            O => \N__13438\,
            I => \N__13296\
        );

    \I__3097\ : ClkMux
    port map (
            O => \N__13437\,
            I => \N__13296\
        );

    \I__3096\ : ClkMux
    port map (
            O => \N__13436\,
            I => \N__13296\
        );

    \I__3095\ : ClkMux
    port map (
            O => \N__13435\,
            I => \N__13296\
        );

    \I__3094\ : ClkMux
    port map (
            O => \N__13434\,
            I => \N__13296\
        );

    \I__3093\ : ClkMux
    port map (
            O => \N__13433\,
            I => \N__13296\
        );

    \I__3092\ : GlobalMux
    port map (
            O => \N__13296\,
            I => clk_48mhz_0
        );

    \I__3091\ : SRMux
    port map (
            O => \N__13293\,
            I => \N__13245\
        );

    \I__3090\ : SRMux
    port map (
            O => \N__13292\,
            I => \N__13245\
        );

    \I__3089\ : SRMux
    port map (
            O => \N__13291\,
            I => \N__13245\
        );

    \I__3088\ : SRMux
    port map (
            O => \N__13290\,
            I => \N__13245\
        );

    \I__3087\ : SRMux
    port map (
            O => \N__13289\,
            I => \N__13245\
        );

    \I__3086\ : SRMux
    port map (
            O => \N__13288\,
            I => \N__13245\
        );

    \I__3085\ : SRMux
    port map (
            O => \N__13287\,
            I => \N__13245\
        );

    \I__3084\ : SRMux
    port map (
            O => \N__13286\,
            I => \N__13245\
        );

    \I__3083\ : SRMux
    port map (
            O => \N__13285\,
            I => \N__13245\
        );

    \I__3082\ : SRMux
    port map (
            O => \N__13284\,
            I => \N__13245\
        );

    \I__3081\ : SRMux
    port map (
            O => \N__13283\,
            I => \N__13245\
        );

    \I__3080\ : SRMux
    port map (
            O => \N__13282\,
            I => \N__13245\
        );

    \I__3079\ : SRMux
    port map (
            O => \N__13281\,
            I => \N__13245\
        );

    \I__3078\ : SRMux
    port map (
            O => \N__13280\,
            I => \N__13245\
        );

    \I__3077\ : SRMux
    port map (
            O => \N__13279\,
            I => \N__13245\
        );

    \I__3076\ : SRMux
    port map (
            O => \N__13278\,
            I => \N__13245\
        );

    \I__3075\ : GlobalMux
    port map (
            O => \N__13245\,
            I => \N__13242\
        );

    \I__3074\ : gio2CtrlBuf
    port map (
            O => \N__13242\,
            I => \wPllLocked_i_g\
        );

    \I__3073\ : InMux
    port map (
            O => \N__13239\,
            I => \N__13235\
        );

    \I__3072\ : InMux
    port map (
            O => \N__13238\,
            I => \N__13232\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__13235\,
            I => \N__13228\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__13232\,
            I => \N__13225\
        );

    \I__3069\ : InMux
    port map (
            O => \N__13231\,
            I => \N__13222\
        );

    \I__3068\ : Span4Mux_v
    port map (
            O => \N__13228\,
            I => \N__13214\
        );

    \I__3067\ : Span4Mux_v
    port map (
            O => \N__13225\,
            I => \N__13214\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__13222\,
            I => \N__13214\
        );

    \I__3065\ : InMux
    port map (
            O => \N__13221\,
            I => \N__13211\
        );

    \I__3064\ : Span4Mux_h
    port map (
            O => \N__13214\,
            I => \N__13208\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__13211\,
            I => \N__13205\
        );

    \I__3062\ : Span4Mux_v
    port map (
            O => \N__13208\,
            I => \N__13202\
        );

    \I__3061\ : Span4Mux_v
    port map (
            O => \N__13205\,
            I => \N__13199\
        );

    \I__3060\ : Odrv4
    port map (
            O => \N__13202\,
            I => \rTxByteZ0Z_3\
        );

    \I__3059\ : Odrv4
    port map (
            O => \N__13199\,
            I => \rTxByteZ0Z_3\
        );

    \I__3058\ : InMux
    port map (
            O => \N__13194\,
            I => \N__13191\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__13191\,
            I => \N__13188\
        );

    \I__3056\ : Odrv4
    port map (
            O => \N__13188\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_3\
        );

    \I__3055\ : CEMux
    port map (
            O => \N__13185\,
            I => \N__13182\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__13182\,
            I => \N__13178\
        );

    \I__3053\ : CEMux
    port map (
            O => \N__13181\,
            I => \N__13175\
        );

    \I__3052\ : Span4Mux_h
    port map (
            O => \N__13178\,
            I => \N__13168\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__13175\,
            I => \N__13168\
        );

    \I__3050\ : CEMux
    port map (
            O => \N__13174\,
            I => \N__13165\
        );

    \I__3049\ : InMux
    port map (
            O => \N__13173\,
            I => \N__13162\
        );

    \I__3048\ : Span4Mux_h
    port map (
            O => \N__13168\,
            I => \N__13159\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__13165\,
            I => \N__13156\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__13162\,
            I => \N__13153\
        );

    \I__3045\ : Odrv4
    port map (
            O => \N__13159\,
            I => \DUT.fifo_tx_inst.N_105\
        );

    \I__3044\ : Odrv12
    port map (
            O => \N__13156\,
            I => \DUT.fifo_tx_inst.N_105\
        );

    \I__3043\ : Odrv4
    port map (
            O => \N__13153\,
            I => \DUT.fifo_tx_inst.N_105\
        );

    \I__3042\ : CascadeMux
    port map (
            O => \N__13146\,
            I => \DUT.N_93_cascade_\
        );

    \I__3041\ : CascadeMux
    port map (
            O => \N__13143\,
            I => \DUT.fifo_tx_inst.N_98_cascade_\
        );

    \I__3040\ : InMux
    port map (
            O => \N__13140\,
            I => \N__13131\
        );

    \I__3039\ : InMux
    port map (
            O => \N__13139\,
            I => \N__13131\
        );

    \I__3038\ : InMux
    port map (
            O => \N__13138\,
            I => \N__13124\
        );

    \I__3037\ : InMux
    port map (
            O => \N__13137\,
            I => \N__13124\
        );

    \I__3036\ : InMux
    port map (
            O => \N__13136\,
            I => \N__13124\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__13131\,
            I => \DUT.fifo_tx_inst.N_86\
        );

    \I__3034\ : LocalMux
    port map (
            O => \N__13124\,
            I => \DUT.fifo_tx_inst.N_86\
        );

    \I__3033\ : InMux
    port map (
            O => \N__13119\,
            I => \N__13116\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__13116\,
            I => \N__13111\
        );

    \I__3031\ : InMux
    port map (
            O => \N__13115\,
            I => \N__13104\
        );

    \I__3030\ : InMux
    port map (
            O => \N__13114\,
            I => \N__13104\
        );

    \I__3029\ : Span12Mux_v
    port map (
            O => \N__13111\,
            I => \N__13101\
        );

    \I__3028\ : InMux
    port map (
            O => \N__13110\,
            I => \N__13098\
        );

    \I__3027\ : InMux
    port map (
            O => \N__13109\,
            I => \N__13095\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__13104\,
            I => \N__13092\
        );

    \I__3025\ : Odrv12
    port map (
            O => \N__13101\,
            I => \DUT.N_93\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__13098\,
            I => \DUT.N_93\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__13095\,
            I => \DUT.N_93\
        );

    \I__3022\ : Odrv12
    port map (
            O => \N__13092\,
            I => \DUT.N_93\
        );

    \I__3021\ : InMux
    port map (
            O => \N__13083\,
            I => \N__13073\
        );

    \I__3020\ : InMux
    port map (
            O => \N__13082\,
            I => \N__13073\
        );

    \I__3019\ : InMux
    port map (
            O => \N__13081\,
            I => \N__13066\
        );

    \I__3018\ : InMux
    port map (
            O => \N__13080\,
            I => \N__13066\
        );

    \I__3017\ : InMux
    port map (
            O => \N__13079\,
            I => \N__13066\
        );

    \I__3016\ : CascadeMux
    port map (
            O => \N__13078\,
            I => \N__13062\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__13073\,
            I => \N__13059\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__13066\,
            I => \N__13056\
        );

    \I__3013\ : CascadeMux
    port map (
            O => \N__13065\,
            I => \N__13053\
        );

    \I__3012\ : InMux
    port map (
            O => \N__13062\,
            I => \N__13049\
        );

    \I__3011\ : Span4Mux_v
    port map (
            O => \N__13059\,
            I => \N__13044\
        );

    \I__3010\ : Span4Mux_v
    port map (
            O => \N__13056\,
            I => \N__13044\
        );

    \I__3009\ : InMux
    port map (
            O => \N__13053\,
            I => \N__13041\
        );

    \I__3008\ : InMux
    port map (
            O => \N__13052\,
            I => \N__13038\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__13049\,
            I => \N__13029\
        );

    \I__3006\ : Span4Mux_h
    port map (
            O => \N__13044\,
            I => \N__13029\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__13041\,
            I => \N__13029\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__13038\,
            I => \N__13029\
        );

    \I__3003\ : Odrv4
    port map (
            O => \N__13029\,
            I => \DUT.rTransmitZ0\
        );

    \I__3002\ : InMux
    port map (
            O => \N__13026\,
            I => \N__13023\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__13023\,
            I => \N__13012\
        );

    \I__3000\ : InMux
    port map (
            O => \N__13022\,
            I => \N__13009\
        );

    \I__2999\ : InMux
    port map (
            O => \N__13021\,
            I => \N__13000\
        );

    \I__2998\ : InMux
    port map (
            O => \N__13020\,
            I => \N__13000\
        );

    \I__2997\ : InMux
    port map (
            O => \N__13019\,
            I => \N__13000\
        );

    \I__2996\ : InMux
    port map (
            O => \N__13018\,
            I => \N__13000\
        );

    \I__2995\ : InMux
    port map (
            O => \N__13017\,
            I => \N__12997\
        );

    \I__2994\ : InMux
    port map (
            O => \N__13016\,
            I => \N__12992\
        );

    \I__2993\ : InMux
    port map (
            O => \N__13015\,
            I => \N__12992\
        );

    \I__2992\ : Span4Mux_v
    port map (
            O => \N__13012\,
            I => \N__12983\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__13009\,
            I => \N__12983\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__13000\,
            I => \N__12983\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__12997\,
            I => \N__12983\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__12992\,
            I => \N__12980\
        );

    \I__2987\ : Span4Mux_h
    port map (
            O => \N__12983\,
            I => \N__12977\
        );

    \I__2986\ : Odrv12
    port map (
            O => \N__12980\,
            I => \rRxReadZ0\
        );

    \I__2985\ : Odrv4
    port map (
            O => \N__12977\,
            I => \rRxReadZ0\
        );

    \I__2984\ : InMux
    port map (
            O => \N__12972\,
            I => \N__12969\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__12969\,
            I => \DUT.fifo_tx_inst.N_98\
        );

    \I__2982\ : InMux
    port map (
            O => \N__12966\,
            I => \N__12963\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__12963\,
            I => \N__12960\
        );

    \I__2980\ : Span4Mux_h
    port map (
            O => \N__12960\,
            I => \N__12956\
        );

    \I__2979\ : InMux
    port map (
            O => \N__12959\,
            I => \N__12953\
        );

    \I__2978\ : Span4Mux_h
    port map (
            O => \N__12956\,
            I => \N__12950\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__12953\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_3\
        );

    \I__2976\ : Odrv4
    port map (
            O => \N__12950\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_3\
        );

    \I__2975\ : InMux
    port map (
            O => \N__12945\,
            I => \N__12942\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__12942\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_0\
        );

    \I__2973\ : InMux
    port map (
            O => \N__12939\,
            I => \N__12936\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__12936\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0\
        );

    \I__2971\ : InMux
    port map (
            O => \N__12933\,
            I => \N__12930\
        );

    \I__2970\ : LocalMux
    port map (
            O => \N__12930\,
            I => \N__12925\
        );

    \I__2969\ : InMux
    port map (
            O => \N__12929\,
            I => \N__12922\
        );

    \I__2968\ : InMux
    port map (
            O => \N__12928\,
            I => \N__12919\
        );

    \I__2967\ : Span4Mux_v
    port map (
            O => \N__12925\,
            I => \N__12911\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__12922\,
            I => \N__12911\
        );

    \I__2965\ : LocalMux
    port map (
            O => \N__12919\,
            I => \N__12911\
        );

    \I__2964\ : InMux
    port map (
            O => \N__12918\,
            I => \N__12908\
        );

    \I__2963\ : Span4Mux_h
    port map (
            O => \N__12911\,
            I => \N__12905\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__12908\,
            I => \N__12902\
        );

    \I__2961\ : Odrv4
    port map (
            O => \N__12905\,
            I => \rTxByteZ0Z_0\
        );

    \I__2960\ : Odrv4
    port map (
            O => \N__12902\,
            I => \rTxByteZ0Z_0\
        );

    \I__2959\ : InMux
    port map (
            O => \N__12897\,
            I => \N__12894\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__12894\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_0\
        );

    \I__2957\ : InMux
    port map (
            O => \N__12891\,
            I => \N__12888\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__12888\,
            I => \N__12883\
        );

    \I__2955\ : InMux
    port map (
            O => \N__12887\,
            I => \N__12880\
        );

    \I__2954\ : InMux
    port map (
            O => \N__12886\,
            I => \N__12877\
        );

    \I__2953\ : Span4Mux_v
    port map (
            O => \N__12883\,
            I => \N__12869\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__12880\,
            I => \N__12869\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__12877\,
            I => \N__12869\
        );

    \I__2950\ : InMux
    port map (
            O => \N__12876\,
            I => \N__12866\
        );

    \I__2949\ : Span4Mux_h
    port map (
            O => \N__12869\,
            I => \N__12863\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__12866\,
            I => \N__12860\
        );

    \I__2947\ : Odrv4
    port map (
            O => \N__12863\,
            I => \rTxByteZ0Z_1\
        );

    \I__2946\ : Odrv4
    port map (
            O => \N__12860\,
            I => \rTxByteZ0Z_1\
        );

    \I__2945\ : InMux
    port map (
            O => \N__12855\,
            I => \N__12852\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__12852\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_1\
        );

    \I__2943\ : InMux
    port map (
            O => \N__12849\,
            I => \N__12840\
        );

    \I__2942\ : InMux
    port map (
            O => \N__12848\,
            I => \N__12840\
        );

    \I__2941\ : InMux
    port map (
            O => \N__12847\,
            I => \N__12829\
        );

    \I__2940\ : InMux
    port map (
            O => \N__12846\,
            I => \N__12829\
        );

    \I__2939\ : InMux
    port map (
            O => \N__12845\,
            I => \N__12826\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__12840\,
            I => \N__12823\
        );

    \I__2937\ : InMux
    port map (
            O => \N__12839\,
            I => \N__12820\
        );

    \I__2936\ : InMux
    port map (
            O => \N__12838\,
            I => \N__12817\
        );

    \I__2935\ : InMux
    port map (
            O => \N__12837\,
            I => \N__12810\
        );

    \I__2934\ : InMux
    port map (
            O => \N__12836\,
            I => \N__12810\
        );

    \I__2933\ : InMux
    port map (
            O => \N__12835\,
            I => \N__12810\
        );

    \I__2932\ : InMux
    port map (
            O => \N__12834\,
            I => \N__12807\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__12829\,
            I => \N__12800\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__12826\,
            I => \N__12800\
        );

    \I__2929\ : Span4Mux_v
    port map (
            O => \N__12823\,
            I => \N__12800\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__12820\,
            I => \N__12795\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__12817\,
            I => \N__12795\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__12810\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__12807\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__2924\ : Odrv4
    port map (
            O => \N__12800\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__2923\ : Odrv4
    port map (
            O => \N__12795\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__2922\ : InMux
    port map (
            O => \N__12786\,
            I => \N__12783\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__12783\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_2\
        );

    \I__2920\ : InMux
    port map (
            O => \N__12780\,
            I => \N__12777\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__12777\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_2\
        );

    \I__2918\ : InMux
    port map (
            O => \N__12774\,
            I => \N__12771\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__12771\,
            I => \N__12768\
        );

    \I__2916\ : Span4Mux_h
    port map (
            O => \N__12768\,
            I => \N__12765\
        );

    \I__2915\ : Odrv4
    port map (
            O => \N__12765\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_2\
        );

    \I__2914\ : CascadeMux
    port map (
            O => \N__12762\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_\
        );

    \I__2913\ : CascadeMux
    port map (
            O => \N__12759\,
            I => \N__12753\
        );

    \I__2912\ : CascadeMux
    port map (
            O => \N__12758\,
            I => \N__12750\
        );

    \I__2911\ : InMux
    port map (
            O => \N__12757\,
            I => \N__12736\
        );

    \I__2910\ : InMux
    port map (
            O => \N__12756\,
            I => \N__12736\
        );

    \I__2909\ : InMux
    port map (
            O => \N__12753\,
            I => \N__12736\
        );

    \I__2908\ : InMux
    port map (
            O => \N__12750\,
            I => \N__12736\
        );

    \I__2907\ : CascadeMux
    port map (
            O => \N__12749\,
            I => \N__12731\
        );

    \I__2906\ : CascadeMux
    port map (
            O => \N__12748\,
            I => \N__12727\
        );

    \I__2905\ : CascadeMux
    port map (
            O => \N__12747\,
            I => \N__12717\
        );

    \I__2904\ : CascadeMux
    port map (
            O => \N__12746\,
            I => \N__12714\
        );

    \I__2903\ : CascadeMux
    port map (
            O => \N__12745\,
            I => \N__12710\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__12736\,
            I => \N__12707\
        );

    \I__2901\ : InMux
    port map (
            O => \N__12735\,
            I => \N__12700\
        );

    \I__2900\ : InMux
    port map (
            O => \N__12734\,
            I => \N__12700\
        );

    \I__2899\ : InMux
    port map (
            O => \N__12731\,
            I => \N__12700\
        );

    \I__2898\ : InMux
    port map (
            O => \N__12730\,
            I => \N__12697\
        );

    \I__2897\ : InMux
    port map (
            O => \N__12727\,
            I => \N__12694\
        );

    \I__2896\ : InMux
    port map (
            O => \N__12726\,
            I => \N__12687\
        );

    \I__2895\ : InMux
    port map (
            O => \N__12725\,
            I => \N__12687\
        );

    \I__2894\ : InMux
    port map (
            O => \N__12724\,
            I => \N__12687\
        );

    \I__2893\ : InMux
    port map (
            O => \N__12723\,
            I => \N__12674\
        );

    \I__2892\ : InMux
    port map (
            O => \N__12722\,
            I => \N__12674\
        );

    \I__2891\ : InMux
    port map (
            O => \N__12721\,
            I => \N__12674\
        );

    \I__2890\ : InMux
    port map (
            O => \N__12720\,
            I => \N__12674\
        );

    \I__2889\ : InMux
    port map (
            O => \N__12717\,
            I => \N__12674\
        );

    \I__2888\ : InMux
    port map (
            O => \N__12714\,
            I => \N__12674\
        );

    \I__2887\ : InMux
    port map (
            O => \N__12713\,
            I => \N__12669\
        );

    \I__2886\ : InMux
    port map (
            O => \N__12710\,
            I => \N__12669\
        );

    \I__2885\ : Span4Mux_h
    port map (
            O => \N__12707\,
            I => \N__12666\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__12700\,
            I => \N__12663\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__12697\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__12694\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__12687\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__12674\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__12669\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__2878\ : Odrv4
    port map (
            O => \N__12666\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__2877\ : Odrv4
    port map (
            O => \N__12663\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__2876\ : InMux
    port map (
            O => \N__12648\,
            I => \N__12645\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__12645\,
            I => \N__12642\
        );

    \I__2874\ : Span4Mux_h
    port map (
            O => \N__12642\,
            I => \N__12639\
        );

    \I__2873\ : Odrv4
    port map (
            O => \N__12639\,
            I => \DUT.rFifoDatarx_2\
        );

    \I__2872\ : InMux
    port map (
            O => \N__12636\,
            I => \N__12632\
        );

    \I__2871\ : InMux
    port map (
            O => \N__12635\,
            I => \N__12628\
        );

    \I__2870\ : LocalMux
    port map (
            O => \N__12632\,
            I => \N__12625\
        );

    \I__2869\ : InMux
    port map (
            O => \N__12631\,
            I => \N__12622\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__12628\,
            I => \N__12619\
        );

    \I__2867\ : Span4Mux_v
    port map (
            O => \N__12625\,
            I => \N__12614\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__12622\,
            I => \N__12614\
        );

    \I__2865\ : Span4Mux_h
    port map (
            O => \N__12619\,
            I => \N__12610\
        );

    \I__2864\ : Span4Mux_h
    port map (
            O => \N__12614\,
            I => \N__12607\
        );

    \I__2863\ : InMux
    port map (
            O => \N__12613\,
            I => \N__12604\
        );

    \I__2862\ : Odrv4
    port map (
            O => \N__12610\,
            I => \rTxByteZ0Z_2\
        );

    \I__2861\ : Odrv4
    port map (
            O => \N__12607\,
            I => \rTxByteZ0Z_2\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__12604\,
            I => \rTxByteZ0Z_2\
        );

    \I__2859\ : CascadeMux
    port map (
            O => \N__12597\,
            I => \N__12594\
        );

    \I__2858\ : InMux
    port map (
            O => \N__12594\,
            I => \N__12591\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__12591\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_2\
        );

    \I__2856\ : InMux
    port map (
            O => \N__12588\,
            I => \N__12585\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__12585\,
            I => \N__12579\
        );

    \I__2854\ : InMux
    port map (
            O => \N__12584\,
            I => \N__12576\
        );

    \I__2853\ : InMux
    port map (
            O => \N__12583\,
            I => \N__12573\
        );

    \I__2852\ : InMux
    port map (
            O => \N__12582\,
            I => \N__12570\
        );

    \I__2851\ : Span4Mux_h
    port map (
            O => \N__12579\,
            I => \N__12567\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__12576\,
            I => \N__12562\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__12573\,
            I => \N__12562\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__12570\,
            I => \N__12559\
        );

    \I__2847\ : Span4Mux_v
    port map (
            O => \N__12567\,
            I => \N__12556\
        );

    \I__2846\ : Span4Mux_h
    port map (
            O => \N__12562\,
            I => \N__12553\
        );

    \I__2845\ : Span4Mux_h
    port map (
            O => \N__12559\,
            I => \N__12550\
        );

    \I__2844\ : Odrv4
    port map (
            O => \N__12556\,
            I => \rTxByteZ0Z_6\
        );

    \I__2843\ : Odrv4
    port map (
            O => \N__12553\,
            I => \rTxByteZ0Z_6\
        );

    \I__2842\ : Odrv4
    port map (
            O => \N__12550\,
            I => \rTxByteZ0Z_6\
        );

    \I__2841\ : InMux
    port map (
            O => \N__12543\,
            I => \N__12540\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__12540\,
            I => \N__12537\
        );

    \I__2839\ : Span4Mux_v
    port map (
            O => \N__12537\,
            I => \N__12534\
        );

    \I__2838\ : Odrv4
    port map (
            O => \N__12534\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_6\
        );

    \I__2837\ : InMux
    port map (
            O => \N__12531\,
            I => \N__12526\
        );

    \I__2836\ : InMux
    port map (
            O => \N__12530\,
            I => \N__12523\
        );

    \I__2835\ : InMux
    port map (
            O => \N__12529\,
            I => \N__12519\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__12526\,
            I => \N__12514\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__12523\,
            I => \N__12514\
        );

    \I__2832\ : InMux
    port map (
            O => \N__12522\,
            I => \N__12511\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__12519\,
            I => \N__12508\
        );

    \I__2830\ : Span4Mux_v
    port map (
            O => \N__12514\,
            I => \N__12505\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__12511\,
            I => \N__12502\
        );

    \I__2828\ : Span4Mux_h
    port map (
            O => \N__12508\,
            I => \N__12499\
        );

    \I__2827\ : Odrv4
    port map (
            O => \N__12505\,
            I => \rTxByteZ0Z_7\
        );

    \I__2826\ : Odrv4
    port map (
            O => \N__12502\,
            I => \rTxByteZ0Z_7\
        );

    \I__2825\ : Odrv4
    port map (
            O => \N__12499\,
            I => \rTxByteZ0Z_7\
        );

    \I__2824\ : InMux
    port map (
            O => \N__12492\,
            I => \N__12489\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__12489\,
            I => \N__12486\
        );

    \I__2822\ : Odrv4
    port map (
            O => \N__12486\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_7\
        );

    \I__2821\ : CascadeMux
    port map (
            O => \N__12483\,
            I => \DUT.fifo_tx_inst.N_101_cascade_\
        );

    \I__2820\ : CascadeMux
    port map (
            O => \N__12480\,
            I => \N__12473\
        );

    \I__2819\ : CascadeMux
    port map (
            O => \N__12479\,
            I => \N__12470\
        );

    \I__2818\ : CascadeMux
    port map (
            O => \N__12478\,
            I => \N__12467\
        );

    \I__2817\ : CascadeMux
    port map (
            O => \N__12477\,
            I => \N__12464\
        );

    \I__2816\ : CascadeMux
    port map (
            O => \N__12476\,
            I => \N__12457\
        );

    \I__2815\ : InMux
    port map (
            O => \N__12473\,
            I => \N__12450\
        );

    \I__2814\ : InMux
    port map (
            O => \N__12470\,
            I => \N__12437\
        );

    \I__2813\ : InMux
    port map (
            O => \N__12467\,
            I => \N__12437\
        );

    \I__2812\ : InMux
    port map (
            O => \N__12464\,
            I => \N__12437\
        );

    \I__2811\ : InMux
    port map (
            O => \N__12463\,
            I => \N__12437\
        );

    \I__2810\ : InMux
    port map (
            O => \N__12462\,
            I => \N__12437\
        );

    \I__2809\ : InMux
    port map (
            O => \N__12461\,
            I => \N__12437\
        );

    \I__2808\ : InMux
    port map (
            O => \N__12460\,
            I => \N__12432\
        );

    \I__2807\ : InMux
    port map (
            O => \N__12457\,
            I => \N__12429\
        );

    \I__2806\ : CascadeMux
    port map (
            O => \N__12456\,
            I => \N__12425\
        );

    \I__2805\ : CascadeMux
    port map (
            O => \N__12455\,
            I => \N__12421\
        );

    \I__2804\ : IoInMux
    port map (
            O => \N__12454\,
            I => \N__12414\
        );

    \I__2803\ : InMux
    port map (
            O => \N__12453\,
            I => \N__12411\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__12450\,
            I => \N__12408\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__12437\,
            I => \N__12405\
        );

    \I__2800\ : InMux
    port map (
            O => \N__12436\,
            I => \N__12402\
        );

    \I__2799\ : InMux
    port map (
            O => \N__12435\,
            I => \N__12399\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__12432\,
            I => \N__12394\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__12429\,
            I => \N__12394\
        );

    \I__2796\ : InMux
    port map (
            O => \N__12428\,
            I => \N__12391\
        );

    \I__2795\ : InMux
    port map (
            O => \N__12425\,
            I => \N__12388\
        );

    \I__2794\ : InMux
    port map (
            O => \N__12424\,
            I => \N__12385\
        );

    \I__2793\ : InMux
    port map (
            O => \N__12421\,
            I => \N__12382\
        );

    \I__2792\ : CascadeMux
    port map (
            O => \N__12420\,
            I => \N__12378\
        );

    \I__2791\ : CascadeMux
    port map (
            O => \N__12419\,
            I => \N__12375\
        );

    \I__2790\ : CascadeMux
    port map (
            O => \N__12418\,
            I => \N__12372\
        );

    \I__2789\ : CascadeMux
    port map (
            O => \N__12417\,
            I => \N__12369\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__12414\,
            I => \N__12363\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__12411\,
            I => \N__12360\
        );

    \I__2786\ : Span4Mux_v
    port map (
            O => \N__12408\,
            I => \N__12351\
        );

    \I__2785\ : Span4Mux_v
    port map (
            O => \N__12405\,
            I => \N__12351\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__12402\,
            I => \N__12351\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__12399\,
            I => \N__12351\
        );

    \I__2782\ : Span4Mux_h
    port map (
            O => \N__12394\,
            I => \N__12340\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__12391\,
            I => \N__12340\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__12388\,
            I => \N__12340\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__12385\,
            I => \N__12340\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__12382\,
            I => \N__12340\
        );

    \I__2777\ : InMux
    port map (
            O => \N__12381\,
            I => \N__12337\
        );

    \I__2776\ : InMux
    port map (
            O => \N__12378\,
            I => \N__12330\
        );

    \I__2775\ : InMux
    port map (
            O => \N__12375\,
            I => \N__12330\
        );

    \I__2774\ : InMux
    port map (
            O => \N__12372\,
            I => \N__12330\
        );

    \I__2773\ : InMux
    port map (
            O => \N__12369\,
            I => \N__12327\
        );

    \I__2772\ : CascadeMux
    port map (
            O => \N__12368\,
            I => \N__12321\
        );

    \I__2771\ : InMux
    port map (
            O => \N__12367\,
            I => \N__12317\
        );

    \I__2770\ : InMux
    port map (
            O => \N__12366\,
            I => \N__12314\
        );

    \I__2769\ : Span4Mux_s1_v
    port map (
            O => \N__12363\,
            I => \N__12309\
        );

    \I__2768\ : Span4Mux_v
    port map (
            O => \N__12360\,
            I => \N__12304\
        );

    \I__2767\ : Span4Mux_v
    port map (
            O => \N__12351\,
            I => \N__12304\
        );

    \I__2766\ : Span4Mux_v
    port map (
            O => \N__12340\,
            I => \N__12299\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__12337\,
            I => \N__12299\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__12330\,
            I => \N__12293\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__12327\,
            I => \N__12290\
        );

    \I__2762\ : InMux
    port map (
            O => \N__12326\,
            I => \N__12283\
        );

    \I__2761\ : InMux
    port map (
            O => \N__12325\,
            I => \N__12283\
        );

    \I__2760\ : InMux
    port map (
            O => \N__12324\,
            I => \N__12283\
        );

    \I__2759\ : InMux
    port map (
            O => \N__12321\,
            I => \N__12278\
        );

    \I__2758\ : InMux
    port map (
            O => \N__12320\,
            I => \N__12278\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__12317\,
            I => \N__12273\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__12314\,
            I => \N__12273\
        );

    \I__2755\ : InMux
    port map (
            O => \N__12313\,
            I => \N__12268\
        );

    \I__2754\ : InMux
    port map (
            O => \N__12312\,
            I => \N__12268\
        );

    \I__2753\ : Sp12to4
    port map (
            O => \N__12309\,
            I => \N__12265\
        );

    \I__2752\ : Span4Mux_h
    port map (
            O => \N__12304\,
            I => \N__12262\
        );

    \I__2751\ : Span4Mux_h
    port map (
            O => \N__12299\,
            I => \N__12259\
        );

    \I__2750\ : InMux
    port map (
            O => \N__12298\,
            I => \N__12254\
        );

    \I__2749\ : InMux
    port map (
            O => \N__12297\,
            I => \N__12254\
        );

    \I__2748\ : InMux
    port map (
            O => \N__12296\,
            I => \N__12251\
        );

    \I__2747\ : Span4Mux_v
    port map (
            O => \N__12293\,
            I => \N__12246\
        );

    \I__2746\ : Span4Mux_v
    port map (
            O => \N__12290\,
            I => \N__12246\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__12283\,
            I => \N__12241\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__12278\,
            I => \N__12241\
        );

    \I__2743\ : Sp12to4
    port map (
            O => \N__12273\,
            I => \N__12236\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__12268\,
            I => \N__12236\
        );

    \I__2741\ : Span12Mux_h
    port map (
            O => \N__12265\,
            I => \N__12233\
        );

    \I__2740\ : Sp12to4
    port map (
            O => \N__12262\,
            I => \N__12224\
        );

    \I__2739\ : Sp12to4
    port map (
            O => \N__12259\,
            I => \N__12224\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__12254\,
            I => \N__12224\
        );

    \I__2737\ : LocalMux
    port map (
            O => \N__12251\,
            I => \N__12224\
        );

    \I__2736\ : Span4Mux_h
    port map (
            O => \N__12246\,
            I => \N__12219\
        );

    \I__2735\ : Span4Mux_v
    port map (
            O => \N__12241\,
            I => \N__12219\
        );

    \I__2734\ : Span12Mux_v
    port map (
            O => \N__12236\,
            I => \N__12216\
        );

    \I__2733\ : Span12Mux_v
    port map (
            O => \N__12233\,
            I => \N__12211\
        );

    \I__2732\ : Span12Mux_h
    port map (
            O => \N__12224\,
            I => \N__12211\
        );

    \I__2731\ : Sp12to4
    port map (
            O => \N__12219\,
            I => \N__12208\
        );

    \I__2730\ : Span12Mux_h
    port map (
            O => \N__12216\,
            I => \N__12203\
        );

    \I__2729\ : Span12Mux_v
    port map (
            O => \N__12211\,
            I => \N__12203\
        );

    \I__2728\ : Span12Mux_h
    port map (
            O => \N__12208\,
            I => \N__12200\
        );

    \I__2727\ : Odrv12
    port map (
            O => \N__12203\,
            I => \wPllLocked\
        );

    \I__2726\ : Odrv12
    port map (
            O => \N__12200\,
            I => \wPllLocked\
        );

    \I__2725\ : CascadeMux
    port map (
            O => \N__12195\,
            I => \DUT.fifo_tx_inst.un1_i11_2_i_cascade_\
        );

    \I__2724\ : CascadeMux
    port map (
            O => \N__12192\,
            I => \N__12172\
        );

    \I__2723\ : InMux
    port map (
            O => \N__12191\,
            I => \N__12156\
        );

    \I__2722\ : InMux
    port map (
            O => \N__12190\,
            I => \N__12153\
        );

    \I__2721\ : InMux
    port map (
            O => \N__12189\,
            I => \N__12150\
        );

    \I__2720\ : InMux
    port map (
            O => \N__12188\,
            I => \N__12147\
        );

    \I__2719\ : InMux
    port map (
            O => \N__12187\,
            I => \N__12144\
        );

    \I__2718\ : InMux
    port map (
            O => \N__12186\,
            I => \N__12141\
        );

    \I__2717\ : InMux
    port map (
            O => \N__12185\,
            I => \N__12130\
        );

    \I__2716\ : InMux
    port map (
            O => \N__12184\,
            I => \N__12130\
        );

    \I__2715\ : InMux
    port map (
            O => \N__12183\,
            I => \N__12130\
        );

    \I__2714\ : InMux
    port map (
            O => \N__12182\,
            I => \N__12130\
        );

    \I__2713\ : InMux
    port map (
            O => \N__12181\,
            I => \N__12130\
        );

    \I__2712\ : InMux
    port map (
            O => \N__12180\,
            I => \N__12125\
        );

    \I__2711\ : InMux
    port map (
            O => \N__12179\,
            I => \N__12125\
        );

    \I__2710\ : InMux
    port map (
            O => \N__12178\,
            I => \N__12118\
        );

    \I__2709\ : InMux
    port map (
            O => \N__12177\,
            I => \N__12118\
        );

    \I__2708\ : InMux
    port map (
            O => \N__12176\,
            I => \N__12118\
        );

    \I__2707\ : InMux
    port map (
            O => \N__12175\,
            I => \N__12115\
        );

    \I__2706\ : InMux
    port map (
            O => \N__12172\,
            I => \N__12112\
        );

    \I__2705\ : InMux
    port map (
            O => \N__12171\,
            I => \N__12105\
        );

    \I__2704\ : InMux
    port map (
            O => \N__12170\,
            I => \N__12105\
        );

    \I__2703\ : InMux
    port map (
            O => \N__12169\,
            I => \N__12105\
        );

    \I__2702\ : SRMux
    port map (
            O => \N__12168\,
            I => \N__12102\
        );

    \I__2701\ : InMux
    port map (
            O => \N__12167\,
            I => \N__12099\
        );

    \I__2700\ : InMux
    port map (
            O => \N__12166\,
            I => \N__12096\
        );

    \I__2699\ : InMux
    port map (
            O => \N__12165\,
            I => \N__12093\
        );

    \I__2698\ : InMux
    port map (
            O => \N__12164\,
            I => \N__12090\
        );

    \I__2697\ : InMux
    port map (
            O => \N__12163\,
            I => \N__12085\
        );

    \I__2696\ : InMux
    port map (
            O => \N__12162\,
            I => \N__12085\
        );

    \I__2695\ : InMux
    port map (
            O => \N__12161\,
            I => \N__12082\
        );

    \I__2694\ : InMux
    port map (
            O => \N__12160\,
            I => \N__12077\
        );

    \I__2693\ : InMux
    port map (
            O => \N__12159\,
            I => \N__12077\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__12156\,
            I => \N__12074\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__12153\,
            I => \N__12071\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__12150\,
            I => \N__12068\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__12147\,
            I => \N__12065\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__12144\,
            I => \N__12062\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__12141\,
            I => \N__12059\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__12130\,
            I => \N__12056\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__12125\,
            I => \N__12053\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__12118\,
            I => \N__12050\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__12115\,
            I => \N__12047\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__12112\,
            I => \N__12044\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__12105\,
            I => \N__12041\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__12102\,
            I => \N__12038\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__12099\,
            I => \N__12035\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__12096\,
            I => \N__12032\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__12093\,
            I => \N__12029\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__12090\,
            I => \N__12026\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__12085\,
            I => \N__12023\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__12082\,
            I => \N__12018\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__12077\,
            I => \N__12015\
        );

    \I__2672\ : Glb2LocalMux
    port map (
            O => \N__12074\,
            I => \N__11946\
        );

    \I__2671\ : Glb2LocalMux
    port map (
            O => \N__12071\,
            I => \N__11946\
        );

    \I__2670\ : Glb2LocalMux
    port map (
            O => \N__12068\,
            I => \N__11946\
        );

    \I__2669\ : Glb2LocalMux
    port map (
            O => \N__12065\,
            I => \N__11946\
        );

    \I__2668\ : Glb2LocalMux
    port map (
            O => \N__12062\,
            I => \N__11946\
        );

    \I__2667\ : Glb2LocalMux
    port map (
            O => \N__12059\,
            I => \N__11946\
        );

    \I__2666\ : Glb2LocalMux
    port map (
            O => \N__12056\,
            I => \N__11946\
        );

    \I__2665\ : Glb2LocalMux
    port map (
            O => \N__12053\,
            I => \N__11946\
        );

    \I__2664\ : Glb2LocalMux
    port map (
            O => \N__12050\,
            I => \N__11946\
        );

    \I__2663\ : Glb2LocalMux
    port map (
            O => \N__12047\,
            I => \N__11946\
        );

    \I__2662\ : Glb2LocalMux
    port map (
            O => \N__12044\,
            I => \N__11946\
        );

    \I__2661\ : Glb2LocalMux
    port map (
            O => \N__12041\,
            I => \N__11946\
        );

    \I__2660\ : Glb2LocalMux
    port map (
            O => \N__12038\,
            I => \N__11946\
        );

    \I__2659\ : Glb2LocalMux
    port map (
            O => \N__12035\,
            I => \N__11946\
        );

    \I__2658\ : Glb2LocalMux
    port map (
            O => \N__12032\,
            I => \N__11946\
        );

    \I__2657\ : Glb2LocalMux
    port map (
            O => \N__12029\,
            I => \N__11946\
        );

    \I__2656\ : Glb2LocalMux
    port map (
            O => \N__12026\,
            I => \N__11946\
        );

    \I__2655\ : Glb2LocalMux
    port map (
            O => \N__12023\,
            I => \N__11946\
        );

    \I__2654\ : CEMux
    port map (
            O => \N__12022\,
            I => \N__11946\
        );

    \I__2653\ : CEMux
    port map (
            O => \N__12021\,
            I => \N__11946\
        );

    \I__2652\ : Glb2LocalMux
    port map (
            O => \N__12018\,
            I => \N__11946\
        );

    \I__2651\ : Glb2LocalMux
    port map (
            O => \N__12015\,
            I => \N__11946\
        );

    \I__2650\ : CEMux
    port map (
            O => \N__12014\,
            I => \N__11946\
        );

    \I__2649\ : CEMux
    port map (
            O => \N__12013\,
            I => \N__11946\
        );

    \I__2648\ : CEMux
    port map (
            O => \N__12012\,
            I => \N__11946\
        );

    \I__2647\ : CEMux
    port map (
            O => \N__12011\,
            I => \N__11946\
        );

    \I__2646\ : CEMux
    port map (
            O => \N__12010\,
            I => \N__11946\
        );

    \I__2645\ : CEMux
    port map (
            O => \N__12009\,
            I => \N__11946\
        );

    \I__2644\ : CEMux
    port map (
            O => \N__12008\,
            I => \N__11946\
        );

    \I__2643\ : CEMux
    port map (
            O => \N__12007\,
            I => \N__11946\
        );

    \I__2642\ : GlobalMux
    port map (
            O => \N__11946\,
            I => \N__11943\
        );

    \I__2641\ : gio2CtrlBuf
    port map (
            O => \N__11943\,
            I => \wPllLocked_g\
        );

    \I__2640\ : InMux
    port map (
            O => \N__11940\,
            I => \N__11936\
        );

    \I__2639\ : InMux
    port map (
            O => \N__11939\,
            I => \N__11933\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__11936\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNIIOZ0Z37\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__11933\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNIIOZ0Z37\
        );

    \I__2636\ : InMux
    port map (
            O => \N__11928\,
            I => \N__11925\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__11925\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_6\
        );

    \I__2634\ : InMux
    port map (
            O => \N__11922\,
            I => \N__11919\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__11919\,
            I => \DUT.fifo_tx_inst.N_101\
        );

    \I__2632\ : InMux
    port map (
            O => \N__11916\,
            I => \N__11913\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__11913\,
            I => \DUT.fifo_tx_inst.un1_i11_2_i\
        );

    \I__2630\ : InMux
    port map (
            O => \N__11910\,
            I => \N__11907\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__11907\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_1\
        );

    \I__2628\ : CascadeMux
    port map (
            O => \N__11904\,
            I => \N__11901\
        );

    \I__2627\ : InMux
    port map (
            O => \N__11901\,
            I => \N__11898\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__11898\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_3\
        );

    \I__2625\ : InMux
    port map (
            O => \N__11895\,
            I => \N__11892\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__11892\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_7\
        );

    \I__2623\ : InMux
    port map (
            O => \N__11889\,
            I => \N__11886\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__11886\,
            I => \N__11883\
        );

    \I__2621\ : Span4Mux_v
    port map (
            O => \N__11883\,
            I => \N__11879\
        );

    \I__2620\ : InMux
    port map (
            O => \N__11882\,
            I => \N__11876\
        );

    \I__2619\ : Odrv4
    port map (
            O => \N__11879\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNIJQZ0Z47\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__11876\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNIJQZ0Z47\
        );

    \I__2617\ : CascadeMux
    port map (
            O => \N__11871\,
            I => \N__11868\
        );

    \I__2616\ : InMux
    port map (
            O => \N__11868\,
            I => \N__11865\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__11865\,
            I => \N__11861\
        );

    \I__2614\ : InMux
    port map (
            O => \N__11864\,
            I => \N__11858\
        );

    \I__2613\ : Odrv4
    port map (
            O => \N__11861\,
            I => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_7\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__11858\,
            I => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_7\
        );

    \I__2611\ : InMux
    port map (
            O => \N__11853\,
            I => \N__11849\
        );

    \I__2610\ : InMux
    port map (
            O => \N__11852\,
            I => \N__11846\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__11849\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIK6NZ0Z4\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__11846\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIK6NZ0Z4\
        );

    \I__2607\ : CascadeMux
    port map (
            O => \N__11841\,
            I => \N__11838\
        );

    \I__2606\ : InMux
    port map (
            O => \N__11838\,
            I => \N__11835\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__11835\,
            I => \N__11832\
        );

    \I__2604\ : Odrv4
    port map (
            O => \N__11832\,
            I => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_4\
        );

    \I__2603\ : CascadeMux
    port map (
            O => \N__11829\,
            I => \N__11826\
        );

    \I__2602\ : InMux
    port map (
            O => \N__11826\,
            I => \N__11823\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__11823\,
            I => \N__11819\
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__11822\,
            I => \N__11815\
        );

    \I__2599\ : Span4Mux_v
    port map (
            O => \N__11819\,
            I => \N__11812\
        );

    \I__2598\ : InMux
    port map (
            O => \N__11818\,
            I => \N__11809\
        );

    \I__2597\ : InMux
    port map (
            O => \N__11815\,
            I => \N__11806\
        );

    \I__2596\ : Odrv4
    port map (
            O => \N__11812\,
            I => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_5\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__11809\,
            I => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_5\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__11806\,
            I => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_5\
        );

    \I__2593\ : CascadeMux
    port map (
            O => \N__11799\,
            I => \N__11796\
        );

    \I__2592\ : InMux
    port map (
            O => \N__11796\,
            I => \N__11792\
        );

    \I__2591\ : InMux
    port map (
            O => \N__11795\,
            I => \N__11789\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__11792\,
            I => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_2\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__11789\,
            I => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_2\
        );

    \I__2588\ : CascadeMux
    port map (
            O => \N__11784\,
            I => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_4_cascade_\
        );

    \I__2587\ : InMux
    port map (
            O => \N__11781\,
            I => \N__11778\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__11778\,
            I => \fifo_inst.tx_fifo_inst.un18_rRamWrAddr_5\
        );

    \I__2585\ : CascadeMux
    port map (
            O => \N__11775\,
            I => \N__11772\
        );

    \I__2584\ : InMux
    port map (
            O => \N__11772\,
            I => \N__11769\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__11769\,
            I => \N__11766\
        );

    \I__2582\ : Odrv4
    port map (
            O => \N__11766\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_1\
        );

    \I__2581\ : CascadeMux
    port map (
            O => \N__11763\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_1_cascade_\
        );

    \I__2580\ : CascadeMux
    port map (
            O => \N__11760\,
            I => \N__11757\
        );

    \I__2579\ : InMux
    port map (
            O => \N__11757\,
            I => \N__11754\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__11754\,
            I => \N__11750\
        );

    \I__2577\ : InMux
    port map (
            O => \N__11753\,
            I => \N__11746\
        );

    \I__2576\ : Span4Mux_v
    port map (
            O => \N__11750\,
            I => \N__11741\
        );

    \I__2575\ : InMux
    port map (
            O => \N__11749\,
            I => \N__11738\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__11746\,
            I => \N__11735\
        );

    \I__2573\ : InMux
    port map (
            O => \N__11745\,
            I => \N__11732\
        );

    \I__2572\ : InMux
    port map (
            O => \N__11744\,
            I => \N__11729\
        );

    \I__2571\ : Odrv4
    port map (
            O => \N__11741\,
            I => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_0\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__11738\,
            I => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_0\
        );

    \I__2569\ : Odrv4
    port map (
            O => \N__11735\,
            I => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_0\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__11732\,
            I => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_0\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__11729\,
            I => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_0\
        );

    \I__2566\ : InMux
    port map (
            O => \N__11718\,
            I => \N__11715\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__11715\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIZ0\
        );

    \I__2564\ : CascadeMux
    port map (
            O => \N__11712\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIZ0_cascade_\
        );

    \I__2563\ : CascadeMux
    port map (
            O => \N__11709\,
            I => \N__11706\
        );

    \I__2562\ : InMux
    port map (
            O => \N__11706\,
            I => \N__11703\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__11703\,
            I => \N__11699\
        );

    \I__2560\ : InMux
    port map (
            O => \N__11702\,
            I => \N__11696\
        );

    \I__2559\ : Odrv4
    port map (
            O => \N__11699\,
            I => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_1\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__11696\,
            I => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_1\
        );

    \I__2557\ : InMux
    port map (
            O => \N__11691\,
            I => \N__11688\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__11688\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7\
        );

    \I__2555\ : InMux
    port map (
            O => \N__11685\,
            I => \N__11681\
        );

    \I__2554\ : InMux
    port map (
            O => \N__11684\,
            I => \N__11678\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__11681\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddr_rst_4\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__11678\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddr_rst_4\
        );

    \I__2551\ : InMux
    port map (
            O => \N__11673\,
            I => \N__11670\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__11670\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddr_0_5\
        );

    \I__2549\ : CascadeMux
    port map (
            O => \N__11667\,
            I => \N__11664\
        );

    \I__2548\ : InMux
    port map (
            O => \N__11664\,
            I => \N__11661\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__11661\,
            I => \N__11656\
        );

    \I__2546\ : InMux
    port map (
            O => \N__11660\,
            I => \N__11653\
        );

    \I__2545\ : CascadeMux
    port map (
            O => \N__11659\,
            I => \N__11650\
        );

    \I__2544\ : Span4Mux_v
    port map (
            O => \N__11656\,
            I => \N__11645\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__11653\,
            I => \N__11645\
        );

    \I__2542\ : InMux
    port map (
            O => \N__11650\,
            I => \N__11642\
        );

    \I__2541\ : Odrv4
    port map (
            O => \N__11645\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_5\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__11642\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_5\
        );

    \I__2539\ : InMux
    port map (
            O => \N__11637\,
            I => \N__11634\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__11634\,
            I => \N__11631\
        );

    \I__2537\ : Odrv4
    port map (
            O => \N__11631\,
            I => \fifo_inst.tx_fifo_inst.un18_rRamWrAddr_4\
        );

    \I__2536\ : InMux
    port map (
            O => \N__11628\,
            I => \N__11624\
        );

    \I__2535\ : InMux
    port map (
            O => \N__11627\,
            I => \N__11621\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__11624\,
            I => \N__11617\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__11621\,
            I => \N__11614\
        );

    \I__2532\ : InMux
    port map (
            O => \N__11620\,
            I => \N__11611\
        );

    \I__2531\ : Odrv12
    port map (
            O => \N__11617\,
            I => \fifo_inst.tx_fifo_inst.un18_rRamWrAddr\
        );

    \I__2530\ : Odrv4
    port map (
            O => \N__11614\,
            I => \fifo_inst.tx_fifo_inst.un18_rRamWrAddr\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__11611\,
            I => \fifo_inst.tx_fifo_inst.un18_rRamWrAddr\
        );

    \I__2528\ : InMux
    port map (
            O => \N__11604\,
            I => \N__11601\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__11601\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_2\
        );

    \I__2526\ : InMux
    port map (
            O => \N__11598\,
            I => \N__11594\
        );

    \I__2525\ : InMux
    port map (
            O => \N__11597\,
            I => \N__11591\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__11594\,
            I => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI6IZ0Z12\
        );

    \I__2523\ : LocalMux
    port map (
            O => \N__11591\,
            I => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI6IZ0Z12\
        );

    \I__2522\ : InMux
    port map (
            O => \N__11586\,
            I => \N__11583\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__11583\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddr_0_3\
        );

    \I__2520\ : InMux
    port map (
            O => \N__11580\,
            I => \N__11570\
        );

    \I__2519\ : InMux
    port map (
            O => \N__11579\,
            I => \N__11570\
        );

    \I__2518\ : InMux
    port map (
            O => \N__11578\,
            I => \N__11567\
        );

    \I__2517\ : InMux
    port map (
            O => \N__11577\,
            I => \N__11564\
        );

    \I__2516\ : InMux
    port map (
            O => \N__11576\,
            I => \N__11559\
        );

    \I__2515\ : InMux
    port map (
            O => \N__11575\,
            I => \N__11559\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__11570\,
            I => \N__11556\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__11567\,
            I => \fifo_inst.rTxRdEn_fast\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__11564\,
            I => \fifo_inst.rTxRdEn_fast\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__11559\,
            I => \fifo_inst.rTxRdEn_fast\
        );

    \I__2510\ : Odrv4
    port map (
            O => \N__11556\,
            I => \fifo_inst.rTxRdEn_fast\
        );

    \I__2509\ : CascadeMux
    port map (
            O => \N__11547\,
            I => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI20CZ0Z4_cascade_\
        );

    \I__2508\ : CascadeMux
    port map (
            O => \N__11544\,
            I => \N__11540\
        );

    \I__2507\ : InMux
    port map (
            O => \N__11543\,
            I => \N__11537\
        );

    \I__2506\ : InMux
    port map (
            O => \N__11540\,
            I => \N__11533\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__11537\,
            I => \N__11530\
        );

    \I__2504\ : InMux
    port map (
            O => \N__11536\,
            I => \N__11527\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__11533\,
            I => \fifo_inst.tx_fifo_inst.un15_rRamRdAddr\
        );

    \I__2502\ : Odrv4
    port map (
            O => \N__11530\,
            I => \fifo_inst.tx_fifo_inst.un15_rRamRdAddr\
        );

    \I__2501\ : LocalMux
    port map (
            O => \N__11527\,
            I => \fifo_inst.tx_fifo_inst.un15_rRamRdAddr\
        );

    \I__2500\ : CascadeMux
    port map (
            O => \N__11520\,
            I => \N__11517\
        );

    \I__2499\ : InMux
    port map (
            O => \N__11517\,
            I => \N__11513\
        );

    \I__2498\ : CascadeMux
    port map (
            O => \N__11516\,
            I => \N__11510\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__11513\,
            I => \N__11507\
        );

    \I__2496\ : InMux
    port map (
            O => \N__11510\,
            I => \N__11504\
        );

    \I__2495\ : Odrv4
    port map (
            O => \N__11507\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_3\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__11504\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_3\
        );

    \I__2493\ : CascadeMux
    port map (
            O => \N__11499\,
            I => \N__11496\
        );

    \I__2492\ : InMux
    port map (
            O => \N__11496\,
            I => \N__11491\
        );

    \I__2491\ : CascadeMux
    port map (
            O => \N__11495\,
            I => \N__11488\
        );

    \I__2490\ : InMux
    port map (
            O => \N__11494\,
            I => \N__11483\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__11491\,
            I => \N__11480\
        );

    \I__2488\ : InMux
    port map (
            O => \N__11488\,
            I => \N__11477\
        );

    \I__2487\ : InMux
    port map (
            O => \N__11487\,
            I => \N__11473\
        );

    \I__2486\ : InMux
    port map (
            O => \N__11486\,
            I => \N__11470\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__11483\,
            I => \N__11467\
        );

    \I__2484\ : Span4Mux_h
    port map (
            O => \N__11480\,
            I => \N__11462\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__11477\,
            I => \N__11462\
        );

    \I__2482\ : InMux
    port map (
            O => \N__11476\,
            I => \N__11459\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__11473\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_0\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__11470\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_0\
        );

    \I__2479\ : Odrv4
    port map (
            O => \N__11467\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_0\
        );

    \I__2478\ : Odrv4
    port map (
            O => \N__11462\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_0\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__11459\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_0\
        );

    \I__2476\ : CascadeMux
    port map (
            O => \N__11448\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_3_cascade_\
        );

    \I__2475\ : CascadeMux
    port map (
            O => \N__11445\,
            I => \N__11440\
        );

    \I__2474\ : InMux
    port map (
            O => \N__11444\,
            I => \N__11437\
        );

    \I__2473\ : InMux
    port map (
            O => \N__11443\,
            I => \N__11434\
        );

    \I__2472\ : InMux
    port map (
            O => \N__11440\,
            I => \N__11431\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__11437\,
            I => \N__11428\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__11434\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_8\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__11431\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_8\
        );

    \I__2468\ : Odrv4
    port map (
            O => \N__11428\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_8\
        );

    \I__2467\ : CascadeMux
    port map (
            O => \N__11421\,
            I => \N__11418\
        );

    \I__2466\ : InMux
    port map (
            O => \N__11418\,
            I => \N__11415\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__11415\,
            I => \fifo_inst.tx_fifo_inst.un15_rRamRdAddr_4\
        );

    \I__2464\ : InMux
    port map (
            O => \N__11412\,
            I => \N__11406\
        );

    \I__2463\ : InMux
    port map (
            O => \N__11411\,
            I => \N__11406\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__11406\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNII2LZ0Z4\
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__11403\,
            I => \N__11399\
        );

    \I__2460\ : CascadeMux
    port map (
            O => \N__11402\,
            I => \N__11396\
        );

    \I__2459\ : InMux
    port map (
            O => \N__11399\,
            I => \N__11393\
        );

    \I__2458\ : InMux
    port map (
            O => \N__11396\,
            I => \N__11390\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__11393\,
            I => \N__11387\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__11390\,
            I => \N__11384\
        );

    \I__2455\ : Odrv4
    port map (
            O => \N__11387\,
            I => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_6\
        );

    \I__2454\ : Odrv4
    port map (
            O => \N__11384\,
            I => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_6\
        );

    \I__2453\ : CascadeMux
    port map (
            O => \N__11379\,
            I => \DUT.fifo_tx_inst.rFifoData_awe3_cascade_\
        );

    \I__2452\ : CascadeMux
    port map (
            O => \N__11376\,
            I => \N__11373\
        );

    \I__2451\ : InMux
    port map (
            O => \N__11373\,
            I => \N__11370\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__11370\,
            I => \DUT.fifo_tx_inst.un1_i11_i\
        );

    \I__2449\ : CascadeMux
    port map (
            O => \N__11367\,
            I => \DUT.fifo_tx_inst.un1_i11_i_cascade_\
        );

    \I__2448\ : InMux
    port map (
            O => \N__11364\,
            I => \N__11357\
        );

    \I__2447\ : InMux
    port map (
            O => \N__11363\,
            I => \N__11354\
        );

    \I__2446\ : InMux
    port map (
            O => \N__11362\,
            I => \N__11347\
        );

    \I__2445\ : InMux
    port map (
            O => \N__11361\,
            I => \N__11347\
        );

    \I__2444\ : InMux
    port map (
            O => \N__11360\,
            I => \N__11347\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__11357\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_1\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__11354\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_1\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__11347\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_1\
        );

    \I__2440\ : CascadeMux
    port map (
            O => \N__11340\,
            I => \N__11332\
        );

    \I__2439\ : CascadeMux
    port map (
            O => \N__11339\,
            I => \N__11329\
        );

    \I__2438\ : InMux
    port map (
            O => \N__11338\,
            I => \N__11324\
        );

    \I__2437\ : InMux
    port map (
            O => \N__11337\,
            I => \N__11324\
        );

    \I__2436\ : InMux
    port map (
            O => \N__11336\,
            I => \N__11315\
        );

    \I__2435\ : InMux
    port map (
            O => \N__11335\,
            I => \N__11315\
        );

    \I__2434\ : InMux
    port map (
            O => \N__11332\,
            I => \N__11315\
        );

    \I__2433\ : InMux
    port map (
            O => \N__11329\,
            I => \N__11315\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__11324\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_0\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__11315\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_0\
        );

    \I__2430\ : InMux
    port map (
            O => \N__11310\,
            I => \N__11306\
        );

    \I__2429\ : InMux
    port map (
            O => \N__11309\,
            I => \N__11303\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__11306\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddr_rst_7\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__11303\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddr_rst_7\
        );

    \I__2426\ : InMux
    port map (
            O => \N__11298\,
            I => \N__11295\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__11295\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddr_0_8\
        );

    \I__2424\ : CEMux
    port map (
            O => \N__11292\,
            I => \N__11289\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__11289\,
            I => \N__11284\
        );

    \I__2422\ : CEMux
    port map (
            O => \N__11288\,
            I => \N__11281\
        );

    \I__2421\ : CEMux
    port map (
            O => \N__11287\,
            I => \N__11278\
        );

    \I__2420\ : Span4Mux_v
    port map (
            O => \N__11284\,
            I => \N__11275\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__11281\,
            I => \N__11272\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__11278\,
            I => \N__11269\
        );

    \I__2417\ : Span4Mux_h
    port map (
            O => \N__11275\,
            I => \N__11266\
        );

    \I__2416\ : Sp12to4
    port map (
            O => \N__11272\,
            I => \N__11261\
        );

    \I__2415\ : Sp12to4
    port map (
            O => \N__11269\,
            I => \N__11261\
        );

    \I__2414\ : Odrv4
    port map (
            O => \N__11266\,
            I => \fifo_inst.rTxRdEn_RNIS0VN\
        );

    \I__2413\ : Odrv12
    port map (
            O => \N__11261\,
            I => \fifo_inst.rTxRdEn_RNIS0VN\
        );

    \I__2412\ : InMux
    port map (
            O => \N__11256\,
            I => \N__11253\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__11253\,
            I => \N__11250\
        );

    \I__2410\ : Odrv4
    port map (
            O => \N__11250\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_3\
        );

    \I__2409\ : InMux
    port map (
            O => \N__11247\,
            I => \N__11244\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__11244\,
            I => \N__11238\
        );

    \I__2407\ : InMux
    port map (
            O => \N__11243\,
            I => \N__11235\
        );

    \I__2406\ : InMux
    port map (
            O => \N__11242\,
            I => \N__11232\
        );

    \I__2405\ : InMux
    port map (
            O => \N__11241\,
            I => \N__11229\
        );

    \I__2404\ : Span4Mux_h
    port map (
            O => \N__11238\,
            I => \N__11226\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__11235\,
            I => \N__11223\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__11232\,
            I => \N__11218\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__11229\,
            I => \N__11218\
        );

    \I__2400\ : Sp12to4
    port map (
            O => \N__11226\,
            I => \N__11215\
        );

    \I__2399\ : Span4Mux_h
    port map (
            O => \N__11223\,
            I => \N__11212\
        );

    \I__2398\ : Span4Mux_h
    port map (
            O => \N__11218\,
            I => \N__11209\
        );

    \I__2397\ : Odrv12
    port map (
            O => \N__11215\,
            I => \rTxByteZ0Z_4\
        );

    \I__2396\ : Odrv4
    port map (
            O => \N__11212\,
            I => \rTxByteZ0Z_4\
        );

    \I__2395\ : Odrv4
    port map (
            O => \N__11209\,
            I => \rTxByteZ0Z_4\
        );

    \I__2394\ : InMux
    port map (
            O => \N__11202\,
            I => \N__11199\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__11199\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_4\
        );

    \I__2392\ : InMux
    port map (
            O => \N__11196\,
            I => \N__11193\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__11193\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_1\
        );

    \I__2390\ : InMux
    port map (
            O => \N__11190\,
            I => \N__11187\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__11187\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_6\
        );

    \I__2388\ : CascadeMux
    port map (
            O => \N__11184\,
            I => \N__11181\
        );

    \I__2387\ : InMux
    port map (
            O => \N__11181\,
            I => \N__11178\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__11178\,
            I => \N__11175\
        );

    \I__2385\ : Odrv4
    port map (
            O => \N__11175\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_7\
        );

    \I__2384\ : InMux
    port map (
            O => \N__11172\,
            I => \N__11168\
        );

    \I__2383\ : InMux
    port map (
            O => \N__11171\,
            I => \N__11165\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__11168\,
            I => \N__11162\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__11165\,
            I => \DUT.fifo_tx_inst.rFifoDataro_1\
        );

    \I__2380\ : Odrv4
    port map (
            O => \N__11162\,
            I => \DUT.fifo_tx_inst.rFifoDataro_1\
        );

    \I__2379\ : CEMux
    port map (
            O => \N__11157\,
            I => \N__11153\
        );

    \I__2378\ : CEMux
    port map (
            O => \N__11156\,
            I => \N__11150\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__11153\,
            I => \N__11147\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__11150\,
            I => \N__11144\
        );

    \I__2375\ : Odrv4
    port map (
            O => \N__11147\,
            I => \DUT.fifo_tx_inst.rFifoData_awe2\
        );

    \I__2374\ : Odrv4
    port map (
            O => \N__11144\,
            I => \DUT.fifo_tx_inst.rFifoData_awe2\
        );

    \I__2373\ : CascadeMux
    port map (
            O => \N__11139\,
            I => \DUT.fifo_tx_inst.rFifoData_awe2_cascade_\
        );

    \I__2372\ : InMux
    port map (
            O => \N__11136\,
            I => \N__11132\
        );

    \I__2371\ : InMux
    port map (
            O => \N__11135\,
            I => \N__11129\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__11132\,
            I => \N__11126\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__11129\,
            I => \DUT.fifo_tx_inst.rFifoDataro_2\
        );

    \I__2368\ : Odrv4
    port map (
            O => \N__11126\,
            I => \DUT.fifo_tx_inst.rFifoDataro_2\
        );

    \I__2367\ : CascadeMux
    port map (
            O => \N__11121\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_\
        );

    \I__2366\ : InMux
    port map (
            O => \N__11118\,
            I => \N__11115\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__11115\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_5\
        );

    \I__2364\ : CascadeMux
    port map (
            O => \N__11112\,
            I => \N__11109\
        );

    \I__2363\ : InMux
    port map (
            O => \N__11109\,
            I => \N__11106\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__11106\,
            I => \DUT.rFifoDatarx_5\
        );

    \I__2361\ : InMux
    port map (
            O => \N__11103\,
            I => \N__11100\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__11100\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_1\
        );

    \I__2359\ : CascadeMux
    port map (
            O => \N__11097\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1_cascade_\
        );

    \I__2358\ : CascadeMux
    port map (
            O => \N__11094\,
            I => \N__11091\
        );

    \I__2357\ : InMux
    port map (
            O => \N__11091\,
            I => \N__11088\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__11088\,
            I => \N__11085\
        );

    \I__2355\ : Odrv4
    port map (
            O => \N__11085\,
            I => \DUT.rFifoDatarx_1\
        );

    \I__2354\ : InMux
    port map (
            O => \N__11082\,
            I => \N__11079\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__11079\,
            I => \N__11075\
        );

    \I__2352\ : InMux
    port map (
            O => \N__11078\,
            I => \N__11072\
        );

    \I__2351\ : Span4Mux_h
    port map (
            O => \N__11075\,
            I => \N__11069\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__11072\,
            I => \DUT.fifo_tx_inst.rFifoDataro_0\
        );

    \I__2349\ : Odrv4
    port map (
            O => \N__11069\,
            I => \DUT.fifo_tx_inst.rFifoDataro_0\
        );

    \I__2348\ : CascadeMux
    port map (
            O => \N__11064\,
            I => \DUT.fifo_tx_inst.rFifoDataror_1_0_cascade_\
        );

    \I__2347\ : CascadeMux
    port map (
            O => \N__11061\,
            I => \N__11056\
        );

    \I__2346\ : InMux
    port map (
            O => \N__11060\,
            I => \N__11042\
        );

    \I__2345\ : InMux
    port map (
            O => \N__11059\,
            I => \N__11042\
        );

    \I__2344\ : InMux
    port map (
            O => \N__11056\,
            I => \N__11042\
        );

    \I__2343\ : InMux
    port map (
            O => \N__11055\,
            I => \N__11042\
        );

    \I__2342\ : InMux
    port map (
            O => \N__11054\,
            I => \N__11033\
        );

    \I__2341\ : InMux
    port map (
            O => \N__11053\,
            I => \N__11033\
        );

    \I__2340\ : InMux
    port map (
            O => \N__11052\,
            I => \N__11033\
        );

    \I__2339\ : InMux
    port map (
            O => \N__11051\,
            I => \N__11033\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__11042\,
            I => \N__11030\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__11033\,
            I => \DUT.rFifoDataror_0\
        );

    \I__2336\ : Odrv4
    port map (
            O => \N__11030\,
            I => \DUT.rFifoDataror_0\
        );

    \I__2335\ : InMux
    port map (
            O => \N__11025\,
            I => \N__11022\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__11022\,
            I => \N__11019\
        );

    \I__2333\ : Odrv4
    port map (
            O => \N__11019\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_0\
        );

    \I__2332\ : InMux
    port map (
            O => \N__11016\,
            I => \N__11013\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__11013\,
            I => \N__11010\
        );

    \I__2330\ : Odrv4
    port map (
            O => \N__11010\,
            I => \DUT.rFifoDatarxZ0Z_0\
        );

    \I__2329\ : CascadeMux
    port map (
            O => \N__11007\,
            I => \N__11004\
        );

    \I__2328\ : InMux
    port map (
            O => \N__11004\,
            I => \N__11001\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__11001\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_0\
        );

    \I__2326\ : InMux
    port map (
            O => \N__10998\,
            I => \N__10995\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__10995\,
            I => \N__10992\
        );

    \I__2324\ : Odrv4
    port map (
            O => \N__10992\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_5\
        );

    \I__2323\ : InMux
    port map (
            O => \N__10989\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_4\
        );

    \I__2322\ : InMux
    port map (
            O => \N__10986\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5\
        );

    \I__2321\ : InMux
    port map (
            O => \N__10983\,
            I => \N__10980\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__10980\,
            I => \N__10977\
        );

    \I__2319\ : Span4Mux_v
    port map (
            O => \N__10977\,
            I => \N__10974\
        );

    \I__2318\ : Odrv4
    port map (
            O => \N__10974\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_7\
        );

    \I__2317\ : InMux
    port map (
            O => \N__10971\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6\
        );

    \I__2316\ : InMux
    port map (
            O => \N__10968\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_7\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__10965\,
            I => \N__10962\
        );

    \I__2314\ : InMux
    port map (
            O => \N__10962\,
            I => \N__10958\
        );

    \I__2313\ : InMux
    port map (
            O => \N__10961\,
            I => \N__10955\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__10958\,
            I => \N__10952\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__10955\,
            I => \N__10949\
        );

    \I__2310\ : Span4Mux_v
    port map (
            O => \N__10952\,
            I => \N__10943\
        );

    \I__2309\ : Span4Mux_v
    port map (
            O => \N__10949\,
            I => \N__10943\
        );

    \I__2308\ : InMux
    port map (
            O => \N__10948\,
            I => \N__10940\
        );

    \I__2307\ : Odrv4
    port map (
            O => \N__10943\,
            I => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_8\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__10940\,
            I => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_8\
        );

    \I__2305\ : CascadeMux
    port map (
            O => \N__10935\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_\
        );

    \I__2304\ : InMux
    port map (
            O => \N__10932\,
            I => \N__10929\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__10929\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_3\
        );

    \I__2302\ : InMux
    port map (
            O => \N__10926\,
            I => \N__10923\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__10923\,
            I => \DUT.rFifoDatarx_3\
        );

    \I__2300\ : InMux
    port map (
            O => \N__10920\,
            I => \N__10917\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__10917\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_4\
        );

    \I__2298\ : InMux
    port map (
            O => \N__10914\,
            I => \N__10911\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__10911\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_7\
        );

    \I__2296\ : InMux
    port map (
            O => \N__10908\,
            I => \N__10905\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__10905\,
            I => \DUT.rFifoDatarx_7\
        );

    \I__2294\ : InMux
    port map (
            O => \N__10902\,
            I => \N__10899\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__10899\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_5\
        );

    \I__2292\ : InMux
    port map (
            O => \N__10896\,
            I => \N__10893\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__10893\,
            I => \fifo_inst.ft2232h_inst.rFifoState_RNIG8PKZ0Z_4\
        );

    \I__2290\ : CascadeMux
    port map (
            O => \N__10890\,
            I => \N__10886\
        );

    \I__2289\ : InMux
    port map (
            O => \N__10889\,
            I => \N__10883\
        );

    \I__2288\ : InMux
    port map (
            O => \N__10886\,
            I => \N__10879\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__10883\,
            I => \N__10876\
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__10882\,
            I => \N__10873\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__10879\,
            I => \N__10870\
        );

    \I__2284\ : Span4Mux_h
    port map (
            O => \N__10876\,
            I => \N__10867\
        );

    \I__2283\ : InMux
    port map (
            O => \N__10873\,
            I => \N__10864\
        );

    \I__2282\ : Odrv4
    port map (
            O => \N__10870\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_7\
        );

    \I__2281\ : Odrv4
    port map (
            O => \N__10867\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_7\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__10864\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_7\
        );

    \I__2279\ : CascadeMux
    port map (
            O => \N__10857\,
            I => \N__10854\
        );

    \I__2278\ : InMux
    port map (
            O => \N__10854\,
            I => \N__10849\
        );

    \I__2277\ : InMux
    port map (
            O => \N__10853\,
            I => \N__10846\
        );

    \I__2276\ : CascadeMux
    port map (
            O => \N__10852\,
            I => \N__10843\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__10849\,
            I => \N__10840\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__10846\,
            I => \N__10837\
        );

    \I__2273\ : InMux
    port map (
            O => \N__10843\,
            I => \N__10834\
        );

    \I__2272\ : Odrv4
    port map (
            O => \N__10840\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_6\
        );

    \I__2271\ : Odrv4
    port map (
            O => \N__10837\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_6\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__10834\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_6\
        );

    \I__2269\ : InMux
    port map (
            O => \N__10827\,
            I => \N__10824\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__10824\,
            I => \fifo_inst.tx_fifo_inst.un15_rRamRdAddr_5\
        );

    \I__2267\ : CascadeMux
    port map (
            O => \N__10821\,
            I => \fifo_inst.tx_fifo_inst.un15_rRamRdAddr_cascade_\
        );

    \I__2266\ : InMux
    port map (
            O => \N__10818\,
            I => \N__10815\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__10815\,
            I => \N__10812\
        );

    \I__2264\ : Odrv4
    port map (
            O => \N__10812\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddr_0_0\
        );

    \I__2263\ : CascadeMux
    port map (
            O => \N__10809\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddr_rst_cascade_\
        );

    \I__2262\ : InMux
    port map (
            O => \N__10806\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1\
        );

    \I__2261\ : InMux
    port map (
            O => \N__10803\,
            I => \N__10800\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__10800\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_3\
        );

    \I__2259\ : InMux
    port map (
            O => \N__10797\,
            I => \N__10794\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__10794\,
            I => \N__10791\
        );

    \I__2257\ : Span4Mux_v
    port map (
            O => \N__10791\,
            I => \N__10787\
        );

    \I__2256\ : InMux
    port map (
            O => \N__10790\,
            I => \N__10784\
        );

    \I__2255\ : Odrv4
    port map (
            O => \N__10787\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIJ4MZ0Z4\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__10784\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIJ4MZ0Z4\
        );

    \I__2253\ : InMux
    port map (
            O => \N__10779\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2\
        );

    \I__2252\ : InMux
    port map (
            O => \N__10776\,
            I => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3\
        );

    \I__2251\ : CascadeMux
    port map (
            O => \N__10773\,
            I => \N__10770\
        );

    \I__2250\ : InMux
    port map (
            O => \N__10770\,
            I => \N__10767\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__10767\,
            I => \N__10763\
        );

    \I__2248\ : CascadeMux
    port map (
            O => \N__10766\,
            I => \N__10759\
        );

    \I__2247\ : Span4Mux_v
    port map (
            O => \N__10763\,
            I => \N__10756\
        );

    \I__2246\ : InMux
    port map (
            O => \N__10762\,
            I => \N__10753\
        );

    \I__2245\ : InMux
    port map (
            O => \N__10759\,
            I => \N__10750\
        );

    \I__2244\ : Odrv4
    port map (
            O => \N__10756\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_2\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__10753\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_2\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__10750\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_2\
        );

    \I__2241\ : InMux
    port map (
            O => \N__10743\,
            I => \N__10737\
        );

    \I__2240\ : InMux
    port map (
            O => \N__10742\,
            I => \N__10737\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__10737\,
            I => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1_c_RNI5GZ0Z02\
        );

    \I__2238\ : InMux
    port map (
            O => \N__10734\,
            I => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1\
        );

    \I__2237\ : InMux
    port map (
            O => \N__10731\,
            I => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2\
        );

    \I__2236\ : CascadeMux
    port map (
            O => \N__10728\,
            I => \N__10725\
        );

    \I__2235\ : InMux
    port map (
            O => \N__10725\,
            I => \N__10721\
        );

    \I__2234\ : InMux
    port map (
            O => \N__10724\,
            I => \N__10717\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__10721\,
            I => \N__10714\
        );

    \I__2232\ : InMux
    port map (
            O => \N__10720\,
            I => \N__10711\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__10717\,
            I => \N__10708\
        );

    \I__2230\ : Odrv4
    port map (
            O => \N__10714\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_4\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__10711\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_4\
        );

    \I__2228\ : Odrv4
    port map (
            O => \N__10708\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_4\
        );

    \I__2227\ : InMux
    port map (
            O => \N__10701\,
            I => \N__10695\
        );

    \I__2226\ : InMux
    port map (
            O => \N__10700\,
            I => \N__10695\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__10695\,
            I => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_3_c_RNI7KZ0Z22\
        );

    \I__2224\ : InMux
    port map (
            O => \N__10692\,
            I => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_3\
        );

    \I__2223\ : InMux
    port map (
            O => \N__10689\,
            I => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_4\
        );

    \I__2222\ : InMux
    port map (
            O => \N__10686\,
            I => \N__10680\
        );

    \I__2221\ : InMux
    port map (
            O => \N__10685\,
            I => \N__10680\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__10680\,
            I => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_5_c_RNI9OZ0Z42\
        );

    \I__2219\ : InMux
    port map (
            O => \N__10677\,
            I => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_5\
        );

    \I__2218\ : InMux
    port map (
            O => \N__10674\,
            I => \N__10668\
        );

    \I__2217\ : InMux
    port map (
            O => \N__10673\,
            I => \N__10668\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__10668\,
            I => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_6_c_RNIAQZ0Z52\
        );

    \I__2215\ : InMux
    port map (
            O => \N__10665\,
            I => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_6\
        );

    \I__2214\ : InMux
    port map (
            O => \N__10662\,
            I => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_7\
        );

    \I__2213\ : InMux
    port map (
            O => \N__10659\,
            I => \N__10656\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__10656\,
            I => \N__10653\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__10653\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_4\
        );

    \I__2210\ : InMux
    port map (
            O => \N__10650\,
            I => \N__10647\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__10647\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddr_0_7\
        );

    \I__2208\ : InMux
    port map (
            O => \N__10644\,
            I => \N__10641\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__10641\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddr_0_4\
        );

    \I__2206\ : InMux
    port map (
            O => \N__10638\,
            I => \N__10635\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__10635\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddr_0_6\
        );

    \I__2204\ : InMux
    port map (
            O => \N__10632\,
            I => \N__10629\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__10629\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_1_1\
        );

    \I__2202\ : CascadeMux
    port map (
            O => \N__10626\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_\
        );

    \I__2201\ : CascadeMux
    port map (
            O => \N__10623\,
            I => \N__10620\
        );

    \I__2200\ : InMux
    port map (
            O => \N__10620\,
            I => \N__10617\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__10617\,
            I => \N__10614\
        );

    \I__2198\ : Span4Mux_h
    port map (
            O => \N__10614\,
            I => \N__10611\
        );

    \I__2197\ : Odrv4
    port map (
            O => \N__10611\,
            I => \DUT.rFifoDatarx_4\
        );

    \I__2196\ : InMux
    port map (
            O => \N__10608\,
            I => \N__10605\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__10605\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_4\
        );

    \I__2194\ : CascadeMux
    port map (
            O => \N__10602\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_\
        );

    \I__2193\ : InMux
    port map (
            O => \N__10599\,
            I => \N__10596\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__10596\,
            I => \N__10593\
        );

    \I__2191\ : Odrv12
    port map (
            O => \N__10593\,
            I => \DUT.rFifoDatarx_6\
        );

    \I__2190\ : InMux
    port map (
            O => \N__10590\,
            I => \N__10587\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__10587\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_4\
        );

    \I__2188\ : InMux
    port map (
            O => \N__10584\,
            I => \N__10581\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__10581\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_6\
        );

    \I__2186\ : InMux
    port map (
            O => \N__10578\,
            I => \N__10575\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__10575\,
            I => \N__10572\
        );

    \I__2184\ : Odrv4
    port map (
            O => \N__10572\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_6\
        );

    \I__2183\ : InMux
    port map (
            O => \N__10569\,
            I => \N__10566\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__10566\,
            I => \N__10563\
        );

    \I__2181\ : Odrv4
    port map (
            O => \N__10563\,
            I => \DUT.uart_inst0.tx_dataZ0Z_4\
        );

    \I__2180\ : InMux
    port map (
            O => \N__10560\,
            I => \N__10557\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__10557\,
            I => \DUT.uart_inst0.tx_dataZ0Z_7\
        );

    \I__2178\ : InMux
    port map (
            O => \N__10554\,
            I => \N__10551\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__10551\,
            I => \DUT.uart_inst0.tx_dataZ0Z_6\
        );

    \I__2176\ : CascadeMux
    port map (
            O => \N__10548\,
            I => \N__10540\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__10547\,
            I => \N__10530\
        );

    \I__2174\ : CascadeMux
    port map (
            O => \N__10546\,
            I => \N__10527\
        );

    \I__2173\ : InMux
    port map (
            O => \N__10545\,
            I => \N__10523\
        );

    \I__2172\ : InMux
    port map (
            O => \N__10544\,
            I => \N__10516\
        );

    \I__2171\ : InMux
    port map (
            O => \N__10543\,
            I => \N__10516\
        );

    \I__2170\ : InMux
    port map (
            O => \N__10540\,
            I => \N__10516\
        );

    \I__2169\ : InMux
    port map (
            O => \N__10539\,
            I => \N__10513\
        );

    \I__2168\ : InMux
    port map (
            O => \N__10538\,
            I => \N__10510\
        );

    \I__2167\ : InMux
    port map (
            O => \N__10537\,
            I => \N__10504\
        );

    \I__2166\ : InMux
    port map (
            O => \N__10536\,
            I => \N__10504\
        );

    \I__2165\ : CascadeMux
    port map (
            O => \N__10535\,
            I => \N__10495\
        );

    \I__2164\ : CascadeMux
    port map (
            O => \N__10534\,
            I => \N__10492\
        );

    \I__2163\ : InMux
    port map (
            O => \N__10533\,
            I => \N__10481\
        );

    \I__2162\ : InMux
    port map (
            O => \N__10530\,
            I => \N__10481\
        );

    \I__2161\ : InMux
    port map (
            O => \N__10527\,
            I => \N__10481\
        );

    \I__2160\ : InMux
    port map (
            O => \N__10526\,
            I => \N__10481\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__10523\,
            I => \N__10476\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__10516\,
            I => \N__10476\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__10513\,
            I => \N__10472\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__10510\,
            I => \N__10469\
        );

    \I__2155\ : CascadeMux
    port map (
            O => \N__10509\,
            I => \N__10465\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__10504\,
            I => \N__10462\
        );

    \I__2153\ : InMux
    port map (
            O => \N__10503\,
            I => \N__10453\
        );

    \I__2152\ : InMux
    port map (
            O => \N__10502\,
            I => \N__10453\
        );

    \I__2151\ : InMux
    port map (
            O => \N__10501\,
            I => \N__10453\
        );

    \I__2150\ : InMux
    port map (
            O => \N__10500\,
            I => \N__10453\
        );

    \I__2149\ : InMux
    port map (
            O => \N__10499\,
            I => \N__10450\
        );

    \I__2148\ : InMux
    port map (
            O => \N__10498\,
            I => \N__10447\
        );

    \I__2147\ : InMux
    port map (
            O => \N__10495\,
            I => \N__10440\
        );

    \I__2146\ : InMux
    port map (
            O => \N__10492\,
            I => \N__10440\
        );

    \I__2145\ : InMux
    port map (
            O => \N__10491\,
            I => \N__10440\
        );

    \I__2144\ : InMux
    port map (
            O => \N__10490\,
            I => \N__10437\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__10481\,
            I => \N__10434\
        );

    \I__2142\ : Span4Mux_v
    port map (
            O => \N__10476\,
            I => \N__10431\
        );

    \I__2141\ : InMux
    port map (
            O => \N__10475\,
            I => \N__10428\
        );

    \I__2140\ : Span4Mux_h
    port map (
            O => \N__10472\,
            I => \N__10423\
        );

    \I__2139\ : Span4Mux_h
    port map (
            O => \N__10469\,
            I => \N__10423\
        );

    \I__2138\ : InMux
    port map (
            O => \N__10468\,
            I => \N__10420\
        );

    \I__2137\ : InMux
    port map (
            O => \N__10465\,
            I => \N__10417\
        );

    \I__2136\ : Span4Mux_h
    port map (
            O => \N__10462\,
            I => \N__10412\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__10453\,
            I => \N__10412\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__10450\,
            I => \DUT.tx_state_0\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__10447\,
            I => \DUT.tx_state_0\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__10440\,
            I => \DUT.tx_state_0\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__10437\,
            I => \DUT.tx_state_0\
        );

    \I__2130\ : Odrv4
    port map (
            O => \N__10434\,
            I => \DUT.tx_state_0\
        );

    \I__2129\ : Odrv4
    port map (
            O => \N__10431\,
            I => \DUT.tx_state_0\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__10428\,
            I => \DUT.tx_state_0\
        );

    \I__2127\ : Odrv4
    port map (
            O => \N__10423\,
            I => \DUT.tx_state_0\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__10420\,
            I => \DUT.tx_state_0\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__10417\,
            I => \DUT.tx_state_0\
        );

    \I__2124\ : Odrv4
    port map (
            O => \N__10412\,
            I => \DUT.tx_state_0\
        );

    \I__2123\ : InMux
    port map (
            O => \N__10389\,
            I => \N__10386\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__10386\,
            I => \DUT.uart_inst0.tx_dataZ0Z_5\
        );

    \I__2121\ : CEMux
    port map (
            O => \N__10383\,
            I => \N__10380\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__10380\,
            I => \N__10377\
        );

    \I__2119\ : Span4Mux_v
    port map (
            O => \N__10377\,
            I => \N__10373\
        );

    \I__2118\ : CEMux
    port map (
            O => \N__10376\,
            I => \N__10370\
        );

    \I__2117\ : Sp12to4
    port map (
            O => \N__10373\,
            I => \N__10365\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__10370\,
            I => \N__10365\
        );

    \I__2115\ : Odrv12
    port map (
            O => \N__10365\,
            I => \DUT.uart_inst0.N_71_i\
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__10362\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_1_1_cascade_\
        );

    \I__2113\ : InMux
    port map (
            O => \N__10359\,
            I => \N__10355\
        );

    \I__2112\ : InMux
    port map (
            O => \N__10358\,
            I => \N__10352\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__10355\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIZ0Z_1\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__10352\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIZ0Z_1\
        );

    \I__2109\ : InMux
    port map (
            O => \N__10347\,
            I => \N__10341\
        );

    \I__2108\ : InMux
    port map (
            O => \N__10346\,
            I => \N__10341\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__10341\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddr_0_1\
        );

    \I__2106\ : CascadeMux
    port map (
            O => \N__10338\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIZ0Z_1_cascade_\
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__10335\,
            I => \N__10332\
        );

    \I__2104\ : InMux
    port map (
            O => \N__10332\,
            I => \N__10329\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__10329\,
            I => \N__10326\
        );

    \I__2102\ : Span4Mux_h
    port map (
            O => \N__10326\,
            I => \N__10323\
        );

    \I__2101\ : Odrv4
    port map (
            O => \N__10323\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_1\
        );

    \I__2100\ : CascadeMux
    port map (
            O => \N__10320\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_1_cascade_\
        );

    \I__2099\ : CascadeMux
    port map (
            O => \N__10317\,
            I => \N__10313\
        );

    \I__2098\ : InMux
    port map (
            O => \N__10316\,
            I => \N__10308\
        );

    \I__2097\ : InMux
    port map (
            O => \N__10313\,
            I => \N__10308\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__10308\,
            I => \DUT.uart_inst0.tx_dataZ0Z_0\
        );

    \I__2095\ : InMux
    port map (
            O => \N__10305\,
            I => \N__10302\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__10302\,
            I => \DUT.uart_inst0.tx_dataZ0Z_1\
        );

    \I__2093\ : InMux
    port map (
            O => \N__10299\,
            I => \N__10296\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__10296\,
            I => \DUT.uart_inst0.tx_dataZ0Z_3\
        );

    \I__2091\ : InMux
    port map (
            O => \N__10293\,
            I => \N__10290\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__10290\,
            I => \DUT.uart_inst0.tx_dataZ0Z_2\
        );

    \I__2089\ : InMux
    port map (
            O => \N__10287\,
            I => \N__10284\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__10284\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_3\
        );

    \I__2087\ : InMux
    port map (
            O => \N__10281\,
            I => \N__10277\
        );

    \I__2086\ : InMux
    port map (
            O => \N__10280\,
            I => \N__10274\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__10277\,
            I => \N__10268\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__10274\,
            I => \N__10268\
        );

    \I__2083\ : InMux
    port map (
            O => \N__10273\,
            I => \N__10265\
        );

    \I__2082\ : Span4Mux_h
    port map (
            O => \N__10268\,
            I => \N__10260\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__10265\,
            I => \N__10257\
        );

    \I__2080\ : InMux
    port map (
            O => \N__10264\,
            I => \N__10254\
        );

    \I__2079\ : InMux
    port map (
            O => \N__10263\,
            I => \N__10251\
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__10260\,
            I => \DUT.wRxByte_4\
        );

    \I__2077\ : Odrv4
    port map (
            O => \N__10257\,
            I => \DUT.wRxByte_4\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__10254\,
            I => \DUT.wRxByte_4\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__10251\,
            I => \DUT.wRxByte_4\
        );

    \I__2074\ : InMux
    port map (
            O => \N__10242\,
            I => \N__10239\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__10239\,
            I => \N__10236\
        );

    \I__2072\ : Odrv4
    port map (
            O => \N__10236\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_4\
        );

    \I__2071\ : InMux
    port map (
            O => \N__10233\,
            I => \N__10230\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__10230\,
            I => \N__10226\
        );

    \I__2069\ : InMux
    port map (
            O => \N__10229\,
            I => \N__10223\
        );

    \I__2068\ : Span4Mux_h
    port map (
            O => \N__10226\,
            I => \N__10217\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__10223\,
            I => \N__10214\
        );

    \I__2066\ : InMux
    port map (
            O => \N__10222\,
            I => \N__10211\
        );

    \I__2065\ : InMux
    port map (
            O => \N__10221\,
            I => \N__10208\
        );

    \I__2064\ : InMux
    port map (
            O => \N__10220\,
            I => \N__10205\
        );

    \I__2063\ : Odrv4
    port map (
            O => \N__10217\,
            I => \DUT.wRxByte_5\
        );

    \I__2062\ : Odrv4
    port map (
            O => \N__10214\,
            I => \DUT.wRxByte_5\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__10211\,
            I => \DUT.wRxByte_5\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__10208\,
            I => \DUT.wRxByte_5\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__10205\,
            I => \DUT.wRxByte_5\
        );

    \I__2058\ : InMux
    port map (
            O => \N__10194\,
            I => \N__10191\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__10191\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_5\
        );

    \I__2056\ : InMux
    port map (
            O => \N__10188\,
            I => \N__10184\
        );

    \I__2055\ : InMux
    port map (
            O => \N__10187\,
            I => \N__10180\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__10184\,
            I => \N__10177\
        );

    \I__2053\ : InMux
    port map (
            O => \N__10183\,
            I => \N__10174\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__10180\,
            I => \N__10171\
        );

    \I__2051\ : Span4Mux_h
    port map (
            O => \N__10177\,
            I => \N__10166\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__10174\,
            I => \N__10163\
        );

    \I__2049\ : Span4Mux_h
    port map (
            O => \N__10171\,
            I => \N__10160\
        );

    \I__2048\ : InMux
    port map (
            O => \N__10170\,
            I => \N__10157\
        );

    \I__2047\ : InMux
    port map (
            O => \N__10169\,
            I => \N__10154\
        );

    \I__2046\ : Odrv4
    port map (
            O => \N__10166\,
            I => \DUT.wRxByte_6\
        );

    \I__2045\ : Odrv4
    port map (
            O => \N__10163\,
            I => \DUT.wRxByte_6\
        );

    \I__2044\ : Odrv4
    port map (
            O => \N__10160\,
            I => \DUT.wRxByte_6\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__10157\,
            I => \DUT.wRxByte_6\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__10154\,
            I => \DUT.wRxByte_6\
        );

    \I__2041\ : InMux
    port map (
            O => \N__10143\,
            I => \N__10140\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__10140\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_6\
        );

    \I__2039\ : InMux
    port map (
            O => \N__10137\,
            I => \N__10133\
        );

    \I__2038\ : InMux
    port map (
            O => \N__10136\,
            I => \N__10130\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__10133\,
            I => \N__10126\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__10130\,
            I => \N__10123\
        );

    \I__2035\ : InMux
    port map (
            O => \N__10129\,
            I => \N__10120\
        );

    \I__2034\ : Span4Mux_v
    port map (
            O => \N__10126\,
            I => \N__10115\
        );

    \I__2033\ : Span4Mux_h
    port map (
            O => \N__10123\,
            I => \N__10112\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__10120\,
            I => \N__10109\
        );

    \I__2031\ : InMux
    port map (
            O => \N__10119\,
            I => \N__10106\
        );

    \I__2030\ : InMux
    port map (
            O => \N__10118\,
            I => \N__10103\
        );

    \I__2029\ : Odrv4
    port map (
            O => \N__10115\,
            I => \DUT.wRxByte_7\
        );

    \I__2028\ : Odrv4
    port map (
            O => \N__10112\,
            I => \DUT.wRxByte_7\
        );

    \I__2027\ : Odrv4
    port map (
            O => \N__10109\,
            I => \DUT.wRxByte_7\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__10106\,
            I => \DUT.wRxByte_7\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__10103\,
            I => \DUT.wRxByte_7\
        );

    \I__2024\ : InMux
    port map (
            O => \N__10092\,
            I => \N__10089\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__10089\,
            I => \N__10086\
        );

    \I__2022\ : Odrv4
    port map (
            O => \N__10086\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_7\
        );

    \I__2021\ : CEMux
    port map (
            O => \N__10083\,
            I => \N__10079\
        );

    \I__2020\ : InMux
    port map (
            O => \N__10082\,
            I => \N__10076\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__10079\,
            I => \N__10073\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__10076\,
            I => \N__10070\
        );

    \I__2017\ : Span4Mux_h
    port map (
            O => \N__10073\,
            I => \N__10067\
        );

    \I__2016\ : Span4Mux_h
    port map (
            O => \N__10070\,
            I => \N__10064\
        );

    \I__2015\ : Odrv4
    port map (
            O => \N__10067\,
            I => \DUT.fifo_rx_inst.rFifoData_awe2\
        );

    \I__2014\ : Odrv4
    port map (
            O => \N__10064\,
            I => \DUT.fifo_rx_inst.rFifoData_awe2\
        );

    \I__2013\ : InMux
    port map (
            O => \N__10059\,
            I => \N__10055\
        );

    \I__2012\ : InMux
    port map (
            O => \N__10058\,
            I => \N__10051\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__10055\,
            I => \N__10048\
        );

    \I__2010\ : InMux
    port map (
            O => \N__10054\,
            I => \N__10045\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__10051\,
            I => \N__10037\
        );

    \I__2008\ : Span4Mux_v
    port map (
            O => \N__10048\,
            I => \N__10037\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__10045\,
            I => \N__10037\
        );

    \I__2006\ : InMux
    port map (
            O => \N__10044\,
            I => \N__10034\
        );

    \I__2005\ : Span4Mux_h
    port map (
            O => \N__10037\,
            I => \N__10031\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__10034\,
            I => \N__10028\
        );

    \I__2003\ : Odrv4
    port map (
            O => \N__10031\,
            I => \DUT.wRxByte_0\
        );

    \I__2002\ : Odrv12
    port map (
            O => \N__10028\,
            I => \DUT.wRxByte_0\
        );

    \I__2001\ : InMux
    port map (
            O => \N__10023\,
            I => \N__10020\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__10020\,
            I => \N__10017\
        );

    \I__1999\ : Odrv4
    port map (
            O => \N__10017\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_0\
        );

    \I__1998\ : CEMux
    port map (
            O => \N__10014\,
            I => \N__10009\
        );

    \I__1997\ : CEMux
    port map (
            O => \N__10013\,
            I => \N__10006\
        );

    \I__1996\ : CEMux
    port map (
            O => \N__10012\,
            I => \N__10003\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__10009\,
            I => \N__10000\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__10006\,
            I => \N__9997\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__10003\,
            I => \N__9994\
        );

    \I__1992\ : Span4Mux_v
    port map (
            O => \N__10000\,
            I => \N__9989\
        );

    \I__1991\ : Span4Mux_v
    port map (
            O => \N__9997\,
            I => \N__9989\
        );

    \I__1990\ : Span4Mux_h
    port map (
            O => \N__9994\,
            I => \N__9985\
        );

    \I__1989\ : Span4Mux_h
    port map (
            O => \N__9989\,
            I => \N__9982\
        );

    \I__1988\ : InMux
    port map (
            O => \N__9988\,
            I => \N__9979\
        );

    \I__1987\ : Odrv4
    port map (
            O => \N__9985\,
            I => \DUT.fifo_rx_inst.rFifoData_awe0\
        );

    \I__1986\ : Odrv4
    port map (
            O => \N__9982\,
            I => \DUT.fifo_rx_inst.rFifoData_awe0\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__9979\,
            I => \DUT.fifo_rx_inst.rFifoData_awe0\
        );

    \I__1984\ : InMux
    port map (
            O => \N__9972\,
            I => \N__9969\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__9969\,
            I => \fifo_inst.tx_fifo_inst.rRamRdAddr_0_2\
        );

    \I__1982\ : CascadeMux
    port map (
            O => \N__9966\,
            I => \N__9955\
        );

    \I__1981\ : CascadeMux
    port map (
            O => \N__9965\,
            I => \N__9950\
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__9964\,
            I => \N__9947\
        );

    \I__1979\ : InMux
    port map (
            O => \N__9963\,
            I => \N__9934\
        );

    \I__1978\ : InMux
    port map (
            O => \N__9962\,
            I => \N__9934\
        );

    \I__1977\ : InMux
    port map (
            O => \N__9961\,
            I => \N__9934\
        );

    \I__1976\ : InMux
    port map (
            O => \N__9960\,
            I => \N__9934\
        );

    \I__1975\ : InMux
    port map (
            O => \N__9959\,
            I => \N__9934\
        );

    \I__1974\ : InMux
    port map (
            O => \N__9958\,
            I => \N__9927\
        );

    \I__1973\ : InMux
    port map (
            O => \N__9955\,
            I => \N__9927\
        );

    \I__1972\ : InMux
    port map (
            O => \N__9954\,
            I => \N__9927\
        );

    \I__1971\ : InMux
    port map (
            O => \N__9953\,
            I => \N__9918\
        );

    \I__1970\ : InMux
    port map (
            O => \N__9950\,
            I => \N__9918\
        );

    \I__1969\ : InMux
    port map (
            O => \N__9947\,
            I => \N__9918\
        );

    \I__1968\ : InMux
    port map (
            O => \N__9946\,
            I => \N__9918\
        );

    \I__1967\ : CascadeMux
    port map (
            O => \N__9945\,
            I => \N__9914\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__9934\,
            I => \N__9905\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__9927\,
            I => \N__9900\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__9918\,
            I => \N__9900\
        );

    \I__1963\ : InMux
    port map (
            O => \N__9917\,
            I => \N__9895\
        );

    \I__1962\ : InMux
    port map (
            O => \N__9914\,
            I => \N__9895\
        );

    \I__1961\ : CascadeMux
    port map (
            O => \N__9913\,
            I => \N__9892\
        );

    \I__1960\ : InMux
    port map (
            O => \N__9912\,
            I => \N__9887\
        );

    \I__1959\ : InMux
    port map (
            O => \N__9911\,
            I => \N__9887\
        );

    \I__1958\ : InMux
    port map (
            O => \N__9910\,
            I => \N__9884\
        );

    \I__1957\ : InMux
    port map (
            O => \N__9909\,
            I => \N__9879\
        );

    \I__1956\ : InMux
    port map (
            O => \N__9908\,
            I => \N__9879\
        );

    \I__1955\ : Span4Mux_h
    port map (
            O => \N__9905\,
            I => \N__9872\
        );

    \I__1954\ : Span4Mux_v
    port map (
            O => \N__9900\,
            I => \N__9872\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__9895\,
            I => \N__9872\
        );

    \I__1952\ : InMux
    port map (
            O => \N__9892\,
            I => \N__9869\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__9887\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__9884\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__9879\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__1948\ : Odrv4
    port map (
            O => \N__9872\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__9869\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__1946\ : CascadeMux
    port map (
            O => \N__9858\,
            I => \N__9855\
        );

    \I__1945\ : InMux
    port map (
            O => \N__9855\,
            I => \N__9852\
        );

    \I__1944\ : LocalMux
    port map (
            O => \N__9852\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2\
        );

    \I__1943\ : CEMux
    port map (
            O => \N__9849\,
            I => \N__9846\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__9846\,
            I => \N__9842\
        );

    \I__1941\ : CEMux
    port map (
            O => \N__9845\,
            I => \N__9839\
        );

    \I__1940\ : Span4Mux_h
    port map (
            O => \N__9842\,
            I => \N__9836\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__9839\,
            I => \N__9833\
        );

    \I__1938\ : Odrv4
    port map (
            O => \N__9836\,
            I => \N_100_i_0\
        );

    \I__1937\ : Odrv12
    port map (
            O => \N__9833\,
            I => \N_100_i_0\
        );

    \I__1936\ : SRMux
    port map (
            O => \N__9828\,
            I => \N__9824\
        );

    \I__1935\ : SRMux
    port map (
            O => \N__9827\,
            I => \N__9821\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__9824\,
            I => \N__9818\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__9821\,
            I => \N__9815\
        );

    \I__1932\ : Span4Mux_v
    port map (
            O => \N__9818\,
            I => \N__9811\
        );

    \I__1931\ : Span4Mux_h
    port map (
            O => \N__9815\,
            I => \N__9808\
        );

    \I__1930\ : InMux
    port map (
            O => \N__9814\,
            I => \N__9805\
        );

    \I__1929\ : Odrv4
    port map (
            O => \N__9811\,
            I => \rFifoDatarff_0_RNIHJV05\
        );

    \I__1928\ : Odrv4
    port map (
            O => \N__9808\,
            I => \rFifoDatarff_0_RNIHJV05\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__9805\,
            I => \rFifoDatarff_0_RNIHJV05\
        );

    \I__1926\ : InMux
    port map (
            O => \N__9798\,
            I => \N__9795\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__9795\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_1\
        );

    \I__1924\ : InMux
    port map (
            O => \N__9792\,
            I => \N__9789\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__9789\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_0\
        );

    \I__1922\ : InMux
    port map (
            O => \N__9786\,
            I => \N__9783\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__9783\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_2\
        );

    \I__1920\ : InMux
    port map (
            O => \N__9780\,
            I => \N__9777\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__9777\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_4\
        );

    \I__1918\ : InMux
    port map (
            O => \N__9774\,
            I => \N__9769\
        );

    \I__1917\ : CEMux
    port map (
            O => \N__9773\,
            I => \N__9766\
        );

    \I__1916\ : CEMux
    port map (
            O => \N__9772\,
            I => \N__9763\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__9769\,
            I => \N__9760\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__9766\,
            I => \N__9757\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__9763\,
            I => \N__9754\
        );

    \I__1912\ : Span4Mux_v
    port map (
            O => \N__9760\,
            I => \N__9751\
        );

    \I__1911\ : Span4Mux_v
    port map (
            O => \N__9757\,
            I => \N__9748\
        );

    \I__1910\ : Span12Mux_h
    port map (
            O => \N__9754\,
            I => \N__9745\
        );

    \I__1909\ : Span4Mux_h
    port map (
            O => \N__9751\,
            I => \N__9742\
        );

    \I__1908\ : Odrv4
    port map (
            O => \N__9748\,
            I => \DUT.fifo_rx_inst.rFifoData_awe3\
        );

    \I__1907\ : Odrv12
    port map (
            O => \N__9745\,
            I => \DUT.fifo_rx_inst.rFifoData_awe3\
        );

    \I__1906\ : Odrv4
    port map (
            O => \N__9742\,
            I => \DUT.fifo_rx_inst.rFifoData_awe3\
        );

    \I__1905\ : InMux
    port map (
            O => \N__9735\,
            I => \N__9732\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__9732\,
            I => \N__9729\
        );

    \I__1903\ : Odrv12
    port map (
            O => \N__9729\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_0\
        );

    \I__1902\ : InMux
    port map (
            O => \N__9726\,
            I => \N__9722\
        );

    \I__1901\ : InMux
    port map (
            O => \N__9725\,
            I => \N__9719\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__9722\,
            I => \N__9714\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__9719\,
            I => \N__9711\
        );

    \I__1898\ : InMux
    port map (
            O => \N__9718\,
            I => \N__9708\
        );

    \I__1897\ : InMux
    port map (
            O => \N__9717\,
            I => \N__9705\
        );

    \I__1896\ : Span4Mux_h
    port map (
            O => \N__9714\,
            I => \N__9701\
        );

    \I__1895\ : Span4Mux_h
    port map (
            O => \N__9711\,
            I => \N__9698\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__9708\,
            I => \N__9695\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__9705\,
            I => \N__9692\
        );

    \I__1892\ : InMux
    port map (
            O => \N__9704\,
            I => \N__9689\
        );

    \I__1891\ : Odrv4
    port map (
            O => \N__9701\,
            I => \DUT.wRxByte_1\
        );

    \I__1890\ : Odrv4
    port map (
            O => \N__9698\,
            I => \DUT.wRxByte_1\
        );

    \I__1889\ : Odrv4
    port map (
            O => \N__9695\,
            I => \DUT.wRxByte_1\
        );

    \I__1888\ : Odrv4
    port map (
            O => \N__9692\,
            I => \DUT.wRxByte_1\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__9689\,
            I => \DUT.wRxByte_1\
        );

    \I__1886\ : CascadeMux
    port map (
            O => \N__9678\,
            I => \N__9675\
        );

    \I__1885\ : InMux
    port map (
            O => \N__9675\,
            I => \N__9672\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__9672\,
            I => \N__9669\
        );

    \I__1883\ : Odrv4
    port map (
            O => \N__9669\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_1\
        );

    \I__1882\ : InMux
    port map (
            O => \N__9666\,
            I => \N__9662\
        );

    \I__1881\ : InMux
    port map (
            O => \N__9665\,
            I => \N__9659\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__9662\,
            I => \N__9653\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__9659\,
            I => \N__9653\
        );

    \I__1878\ : InMux
    port map (
            O => \N__9658\,
            I => \N__9650\
        );

    \I__1877\ : Span4Mux_v
    port map (
            O => \N__9653\,
            I => \N__9645\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__9650\,
            I => \N__9642\
        );

    \I__1875\ : InMux
    port map (
            O => \N__9649\,
            I => \N__9639\
        );

    \I__1874\ : InMux
    port map (
            O => \N__9648\,
            I => \N__9636\
        );

    \I__1873\ : Odrv4
    port map (
            O => \N__9645\,
            I => \DUT.wRxByte_2\
        );

    \I__1872\ : Odrv4
    port map (
            O => \N__9642\,
            I => \DUT.wRxByte_2\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__9639\,
            I => \DUT.wRxByte_2\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__9636\,
            I => \DUT.wRxByte_2\
        );

    \I__1869\ : InMux
    port map (
            O => \N__9627\,
            I => \N__9624\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__9624\,
            I => \N__9621\
        );

    \I__1867\ : Odrv4
    port map (
            O => \N__9621\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_2\
        );

    \I__1866\ : InMux
    port map (
            O => \N__9618\,
            I => \N__9615\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__9615\,
            I => \N__9611\
        );

    \I__1864\ : InMux
    port map (
            O => \N__9614\,
            I => \N__9608\
        );

    \I__1863\ : Span4Mux_h
    port map (
            O => \N__9611\,
            I => \N__9602\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__9608\,
            I => \N__9599\
        );

    \I__1861\ : InMux
    port map (
            O => \N__9607\,
            I => \N__9596\
        );

    \I__1860\ : InMux
    port map (
            O => \N__9606\,
            I => \N__9593\
        );

    \I__1859\ : InMux
    port map (
            O => \N__9605\,
            I => \N__9590\
        );

    \I__1858\ : Odrv4
    port map (
            O => \N__9602\,
            I => \DUT.wRxByte_3\
        );

    \I__1857\ : Odrv4
    port map (
            O => \N__9599\,
            I => \DUT.wRxByte_3\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__9596\,
            I => \DUT.wRxByte_3\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__9593\,
            I => \DUT.wRxByte_3\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__9590\,
            I => \DUT.wRxByte_3\
        );

    \I__1853\ : InMux
    port map (
            O => \N__9579\,
            I => \N__9575\
        );

    \I__1852\ : InMux
    port map (
            O => \N__9578\,
            I => \N__9572\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__9575\,
            I => \DUT.fifo_rx_inst.rFifoDataro_3\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__9572\,
            I => \DUT.fifo_rx_inst.rFifoDataro_3\
        );

    \I__1849\ : InMux
    port map (
            O => \N__9567\,
            I => \N__9564\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__9564\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_1\
        );

    \I__1847\ : InMux
    port map (
            O => \N__9561\,
            I => \N__9558\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__9558\,
            I => \fifo_inst.ft2232h_inst.N_103\
        );

    \I__1845\ : InMux
    port map (
            O => \N__9555\,
            I => \N__9551\
        );

    \I__1844\ : InMux
    port map (
            O => \N__9554\,
            I => \N__9548\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__9551\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_2\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__9548\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_2\
        );

    \I__1841\ : InMux
    port map (
            O => \N__9543\,
            I => \N__9539\
        );

    \I__1840\ : InMux
    port map (
            O => \N__9542\,
            I => \N__9536\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__9539\,
            I => \DUT.fifo_rx_inst.rFifoDataro_2\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__9536\,
            I => \DUT.fifo_rx_inst.rFifoDataro_2\
        );

    \I__1837\ : CascadeMux
    port map (
            O => \N__9531\,
            I => \N__9528\
        );

    \I__1836\ : InMux
    port map (
            O => \N__9528\,
            I => \N__9521\
        );

    \I__1835\ : InMux
    port map (
            O => \N__9527\,
            I => \N__9516\
        );

    \I__1834\ : InMux
    port map (
            O => \N__9526\,
            I => \N__9516\
        );

    \I__1833\ : InMux
    port map (
            O => \N__9525\,
            I => \N__9511\
        );

    \I__1832\ : InMux
    port map (
            O => \N__9524\,
            I => \N__9511\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__9521\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_0\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__9516\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_0\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__9511\,
            I => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_0\
        );

    \I__1828\ : InMux
    port map (
            O => \N__9504\,
            I => \N__9499\
        );

    \I__1827\ : InMux
    port map (
            O => \N__9503\,
            I => \N__9494\
        );

    \I__1826\ : InMux
    port map (
            O => \N__9502\,
            I => \N__9494\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__9499\,
            I => \N__9491\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__9494\,
            I => \N__9488\
        );

    \I__1823\ : Span4Mux_h
    port map (
            O => \N__9491\,
            I => \N__9485\
        );

    \I__1822\ : Span4Mux_h
    port map (
            O => \N__9488\,
            I => \N__9482\
        );

    \I__1821\ : Span4Mux_v
    port map (
            O => \N__9485\,
            I => \N__9479\
        );

    \I__1820\ : Sp12to4
    port map (
            O => \N__9482\,
            I => \N__9476\
        );

    \I__1819\ : Span4Mux_v
    port map (
            O => \N__9479\,
            I => \N__9473\
        );

    \I__1818\ : Span12Mux_v
    port map (
            O => \N__9476\,
            I => \N__9470\
        );

    \I__1817\ : Span4Mux_v
    port map (
            O => \N__9473\,
            I => \N__9467\
        );

    \I__1816\ : Odrv12
    port map (
            O => \N__9470\,
            I => \iTxE_n_c\
        );

    \I__1815\ : Odrv4
    port map (
            O => \N__9467\,
            I => \iTxE_n_c\
        );

    \I__1814\ : InMux
    port map (
            O => \N__9462\,
            I => \N__9455\
        );

    \I__1813\ : InMux
    port map (
            O => \N__9461\,
            I => \N__9455\
        );

    \I__1812\ : InMux
    port map (
            O => \N__9460\,
            I => \N__9450\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__9455\,
            I => \N__9447\
        );

    \I__1810\ : InMux
    port map (
            O => \N__9454\,
            I => \N__9442\
        );

    \I__1809\ : InMux
    port map (
            O => \N__9453\,
            I => \N__9442\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__9450\,
            I => \N__9435\
        );

    \I__1807\ : Span4Mux_h
    port map (
            O => \N__9447\,
            I => \N__9435\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__9442\,
            I => \N__9435\
        );

    \I__1805\ : Span4Mux_v
    port map (
            O => \N__9435\,
            I => \N__9432\
        );

    \I__1804\ : Sp12to4
    port map (
            O => \N__9432\,
            I => \N__9429\
        );

    \I__1803\ : Span12Mux_h
    port map (
            O => \N__9429\,
            I => \N__9426\
        );

    \I__1802\ : Odrv12
    port map (
            O => \N__9426\,
            I => \iRxF_n_c\
        );

    \I__1801\ : CascadeMux
    port map (
            O => \N__9423\,
            I => \N__9420\
        );

    \I__1800\ : InMux
    port map (
            O => \N__9420\,
            I => \N__9417\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__9417\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_0\
        );

    \I__1798\ : InMux
    port map (
            O => \N__9414\,
            I => \N__9408\
        );

    \I__1797\ : InMux
    port map (
            O => \N__9413\,
            I => \N__9401\
        );

    \I__1796\ : InMux
    port map (
            O => \N__9412\,
            I => \N__9401\
        );

    \I__1795\ : InMux
    port map (
            O => \N__9411\,
            I => \N__9401\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__9408\,
            I => \N__9390\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__9401\,
            I => \N__9387\
        );

    \I__1792\ : InMux
    port map (
            O => \N__9400\,
            I => \N__9382\
        );

    \I__1791\ : InMux
    port map (
            O => \N__9399\,
            I => \N__9382\
        );

    \I__1790\ : InMux
    port map (
            O => \N__9398\,
            I => \N__9374\
        );

    \I__1789\ : InMux
    port map (
            O => \N__9397\,
            I => \N__9374\
        );

    \I__1788\ : InMux
    port map (
            O => \N__9396\,
            I => \N__9374\
        );

    \I__1787\ : InMux
    port map (
            O => \N__9395\,
            I => \N__9367\
        );

    \I__1786\ : InMux
    port map (
            O => \N__9394\,
            I => \N__9367\
        );

    \I__1785\ : InMux
    port map (
            O => \N__9393\,
            I => \N__9367\
        );

    \I__1784\ : Span4Mux_h
    port map (
            O => \N__9390\,
            I => \N__9360\
        );

    \I__1783\ : Span4Mux_v
    port map (
            O => \N__9387\,
            I => \N__9360\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__9382\,
            I => \N__9360\
        );

    \I__1781\ : InMux
    port map (
            O => \N__9381\,
            I => \N__9357\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__9374\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__9367\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__1778\ : Odrv4
    port map (
            O => \N__9360\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__9357\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__1776\ : CascadeMux
    port map (
            O => \N__9348\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_\
        );

    \I__1775\ : CascadeMux
    port map (
            O => \N__9345\,
            I => \N__9342\
        );

    \I__1774\ : InMux
    port map (
            O => \N__9342\,
            I => \N__9339\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__9339\,
            I => \N__9336\
        );

    \I__1772\ : Span4Mux_h
    port map (
            O => \N__9336\,
            I => \N__9333\
        );

    \I__1771\ : Odrv4
    port map (
            O => \N__9333\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7\
        );

    \I__1770\ : InMux
    port map (
            O => \N__9330\,
            I => \N__9327\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__9327\,
            I => \N__9324\
        );

    \I__1768\ : Span4Mux_h
    port map (
            O => \N__9324\,
            I => \N__9321\
        );

    \I__1767\ : Odrv4
    port map (
            O => \N__9321\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_7\
        );

    \I__1766\ : InMux
    port map (
            O => \N__9318\,
            I => \N__9315\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__9315\,
            I => \N__9312\
        );

    \I__1764\ : Span4Mux_h
    port map (
            O => \N__9312\,
            I => \N__9309\
        );

    \I__1763\ : Odrv4
    port map (
            O => \N__9309\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1\
        );

    \I__1762\ : InMux
    port map (
            O => \N__9306\,
            I => \N__9303\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__9303\,
            I => \N__9292\
        );

    \I__1760\ : InMux
    port map (
            O => \N__9302\,
            I => \N__9287\
        );

    \I__1759\ : InMux
    port map (
            O => \N__9301\,
            I => \N__9287\
        );

    \I__1758\ : InMux
    port map (
            O => \N__9300\,
            I => \N__9282\
        );

    \I__1757\ : InMux
    port map (
            O => \N__9299\,
            I => \N__9282\
        );

    \I__1756\ : InMux
    port map (
            O => \N__9298\,
            I => \N__9279\
        );

    \I__1755\ : InMux
    port map (
            O => \N__9297\,
            I => \N__9274\
        );

    \I__1754\ : InMux
    port map (
            O => \N__9296\,
            I => \N__9274\
        );

    \I__1753\ : InMux
    port map (
            O => \N__9295\,
            I => \N__9271\
        );

    \I__1752\ : Span4Mux_h
    port map (
            O => \N__9292\,
            I => \N__9268\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__9287\,
            I => \N__9263\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__9282\,
            I => \N__9263\
        );

    \I__1749\ : LocalMux
    port map (
            O => \N__9279\,
            I => \DUT.uart_inst0.N_77\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__9274\,
            I => \DUT.uart_inst0.N_77\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__9271\,
            I => \DUT.uart_inst0.N_77\
        );

    \I__1746\ : Odrv4
    port map (
            O => \N__9268\,
            I => \DUT.uart_inst0.N_77\
        );

    \I__1745\ : Odrv4
    port map (
            O => \N__9263\,
            I => \DUT.uart_inst0.N_77\
        );

    \I__1744\ : InMux
    port map (
            O => \N__9252\,
            I => \N__9249\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__9249\,
            I => \DUT.uart_inst0.tx_bits_remaining_RNO_0Z0Z_3\
        );

    \I__1742\ : InMux
    port map (
            O => \N__9246\,
            I => \N__9243\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__9243\,
            I => \DUT.uart_inst0.tx_bits_remaining_RNIAIE4LZ0Z_1\
        );

    \I__1740\ : CascadeMux
    port map (
            O => \N__9240\,
            I => \N__9236\
        );

    \I__1739\ : InMux
    port map (
            O => \N__9239\,
            I => \N__9232\
        );

    \I__1738\ : InMux
    port map (
            O => \N__9236\,
            I => \N__9229\
        );

    \I__1737\ : InMux
    port map (
            O => \N__9235\,
            I => \N__9226\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__9232\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_1\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__9229\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_1\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__9226\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_1\
        );

    \I__1733\ : CascadeMux
    port map (
            O => \N__9219\,
            I => \N__9216\
        );

    \I__1732\ : InMux
    port map (
            O => \N__9216\,
            I => \N__9213\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__9213\,
            I => \N__9207\
        );

    \I__1730\ : InMux
    port map (
            O => \N__9212\,
            I => \N__9204\
        );

    \I__1729\ : InMux
    port map (
            O => \N__9211\,
            I => \N__9201\
        );

    \I__1728\ : InMux
    port map (
            O => \N__9210\,
            I => \N__9198\
        );

    \I__1727\ : Span4Mux_h
    port map (
            O => \N__9207\,
            I => \N__9195\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__9204\,
            I => \N__9192\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__9201\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_0\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__9198\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_0\
        );

    \I__1723\ : Odrv4
    port map (
            O => \N__9195\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_0\
        );

    \I__1722\ : Odrv4
    port map (
            O => \N__9192\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_0\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__9183\,
            I => \N__9179\
        );

    \I__1720\ : InMux
    port map (
            O => \N__9182\,
            I => \N__9174\
        );

    \I__1719\ : InMux
    port map (
            O => \N__9179\,
            I => \N__9168\
        );

    \I__1718\ : InMux
    port map (
            O => \N__9178\,
            I => \N__9168\
        );

    \I__1717\ : InMux
    port map (
            O => \N__9177\,
            I => \N__9165\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__9174\,
            I => \N__9162\
        );

    \I__1715\ : InMux
    port map (
            O => \N__9173\,
            I => \N__9159\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__9168\,
            I => \N__9156\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__9165\,
            I => \N__9149\
        );

    \I__1712\ : Span4Mux_h
    port map (
            O => \N__9162\,
            I => \N__9149\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__9159\,
            I => \N__9149\
        );

    \I__1710\ : Odrv12
    port map (
            O => \N__9156\,
            I => \DUT.uart_inst0.N_124\
        );

    \I__1709\ : Odrv4
    port map (
            O => \N__9149\,
            I => \DUT.uart_inst0.N_124\
        );

    \I__1708\ : CascadeMux
    port map (
            O => \N__9144\,
            I => \N__9141\
        );

    \I__1707\ : InMux
    port map (
            O => \N__9141\,
            I => \N__9136\
        );

    \I__1706\ : InMux
    port map (
            O => \N__9140\,
            I => \N__9131\
        );

    \I__1705\ : InMux
    port map (
            O => \N__9139\,
            I => \N__9131\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__9136\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_2\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__9131\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_2\
        );

    \I__1702\ : InMux
    port map (
            O => \N__9126\,
            I => \N__9123\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__9123\,
            I => \DUT.uart_inst0.tx_bits_remaining_RNIBJE4LZ0Z_2\
        );

    \I__1700\ : CascadeMux
    port map (
            O => \N__9120\,
            I => \N__9116\
        );

    \I__1699\ : InMux
    port map (
            O => \N__9119\,
            I => \N__9111\
        );

    \I__1698\ : InMux
    port map (
            O => \N__9116\,
            I => \N__9111\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__9111\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_3\
        );

    \I__1696\ : InMux
    port map (
            O => \N__9108\,
            I => \N__9103\
        );

    \I__1695\ : InMux
    port map (
            O => \N__9107\,
            I => \N__9096\
        );

    \I__1694\ : InMux
    port map (
            O => \N__9106\,
            I => \N__9093\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__9103\,
            I => \N__9090\
        );

    \I__1692\ : InMux
    port map (
            O => \N__9102\,
            I => \N__9083\
        );

    \I__1691\ : InMux
    port map (
            O => \N__9101\,
            I => \N__9083\
        );

    \I__1690\ : InMux
    port map (
            O => \N__9100\,
            I => \N__9083\
        );

    \I__1689\ : InMux
    port map (
            O => \N__9099\,
            I => \N__9080\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__9096\,
            I => \DUT.uart_inst0.N_96\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__9093\,
            I => \DUT.uart_inst0.N_96\
        );

    \I__1686\ : Odrv4
    port map (
            O => \N__9090\,
            I => \DUT.uart_inst0.N_96\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__9083\,
            I => \DUT.uart_inst0.N_96\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__9080\,
            I => \DUT.uart_inst0.N_96\
        );

    \I__1683\ : InMux
    port map (
            O => \N__9069\,
            I => \N__9064\
        );

    \I__1682\ : InMux
    port map (
            O => \N__9068\,
            I => \N__9061\
        );

    \I__1681\ : InMux
    port map (
            O => \N__9067\,
            I => \N__9055\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__9064\,
            I => \N__9050\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__9061\,
            I => \N__9050\
        );

    \I__1678\ : InMux
    port map (
            O => \N__9060\,
            I => \N__9043\
        );

    \I__1677\ : InMux
    port map (
            O => \N__9059\,
            I => \N__9043\
        );

    \I__1676\ : InMux
    port map (
            O => \N__9058\,
            I => \N__9043\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__9055\,
            I => \DUT.uart_inst0.N_99\
        );

    \I__1674\ : Odrv4
    port map (
            O => \N__9050\,
            I => \DUT.uart_inst0.N_99\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__9043\,
            I => \DUT.uart_inst0.N_99\
        );

    \I__1672\ : InMux
    port map (
            O => \N__9036\,
            I => \N__9033\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__9033\,
            I => \DUT.uart_inst0.un1_tx_bits_remaining_axb_3\
        );

    \I__1670\ : IoInMux
    port map (
            O => \N__9030\,
            I => \N__9026\
        );

    \I__1669\ : IoInMux
    port map (
            O => \N__9029\,
            I => \N__9023\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__9026\,
            I => \N__9020\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__9023\,
            I => \N__9017\
        );

    \I__1666\ : Span4Mux_s0_v
    port map (
            O => \N__9020\,
            I => \N__9014\
        );

    \I__1665\ : Span4Mux_s2_v
    port map (
            O => \N__9017\,
            I => \N__9011\
        );

    \I__1664\ : Sp12to4
    port map (
            O => \N__9014\,
            I => \N__9008\
        );

    \I__1663\ : Span4Mux_v
    port map (
            O => \N__9011\,
            I => \N__9005\
        );

    \I__1662\ : Span12Mux_h
    port map (
            O => \N__9008\,
            I => \N__9002\
        );

    \I__1661\ : Span4Mux_v
    port map (
            O => \N__9005\,
            I => \N__8999\
        );

    \I__1660\ : Span12Mux_v
    port map (
            O => \N__9002\,
            I => \N__8995\
        );

    \I__1659\ : Span4Mux_v
    port map (
            O => \N__8999\,
            I => \N__8992\
        );

    \I__1658\ : InMux
    port map (
            O => \N__8998\,
            I => \N__8989\
        );

    \I__1657\ : Odrv12
    port map (
            O => \N__8995\,
            I => \P1A4_c\
        );

    \I__1656\ : Odrv4
    port map (
            O => \N__8992\,
            I => \P1A4_c\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__8989\,
            I => \P1A4_c\
        );

    \I__1654\ : CascadeMux
    port map (
            O => \N__8982\,
            I => \DUT.uart_inst0.tx_countdown_7_i_a3_0_sx_3_cascade_\
        );

    \I__1653\ : InMux
    port map (
            O => \N__8979\,
            I => \N__8976\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__8976\,
            I => \DUT.uart_inst0.N_116\
        );

    \I__1651\ : SRMux
    port map (
            O => \N__8973\,
            I => \N__8969\
        );

    \I__1650\ : SRMux
    port map (
            O => \N__8972\,
            I => \N__8966\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__8969\,
            I => \N__8963\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__8966\,
            I => \N__8960\
        );

    \I__1647\ : Odrv4
    port map (
            O => \N__8963\,
            I => \DUT.uart_inst0.N_76_i\
        );

    \I__1646\ : Odrv4
    port map (
            O => \N__8960\,
            I => \DUT.uart_inst0.N_76_i\
        );

    \I__1645\ : CascadeMux
    port map (
            O => \N__8955\,
            I => \N__8947\
        );

    \I__1644\ : InMux
    port map (
            O => \N__8954\,
            I => \N__8944\
        );

    \I__1643\ : InMux
    port map (
            O => \N__8953\,
            I => \N__8939\
        );

    \I__1642\ : InMux
    port map (
            O => \N__8952\,
            I => \N__8939\
        );

    \I__1641\ : InMux
    port map (
            O => \N__8951\,
            I => \N__8936\
        );

    \I__1640\ : InMux
    port map (
            O => \N__8950\,
            I => \N__8933\
        );

    \I__1639\ : InMux
    port map (
            O => \N__8947\,
            I => \N__8930\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__8944\,
            I => \N__8927\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__8939\,
            I => \N__8924\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__8936\,
            I => \N__8921\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__8933\,
            I => \DUT.uart_inst0.tx_countdown_3_2\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__8930\,
            I => \DUT.uart_inst0.tx_countdown_3_2\
        );

    \I__1633\ : Odrv4
    port map (
            O => \N__8927\,
            I => \DUT.uart_inst0.tx_countdown_3_2\
        );

    \I__1632\ : Odrv4
    port map (
            O => \N__8924\,
            I => \DUT.uart_inst0.tx_countdown_3_2\
        );

    \I__1631\ : Odrv4
    port map (
            O => \N__8921\,
            I => \DUT.uart_inst0.tx_countdown_3_2\
        );

    \I__1630\ : CascadeMux
    port map (
            O => \N__8910\,
            I => \N__8905\
        );

    \I__1629\ : InMux
    port map (
            O => \N__8909\,
            I => \N__8900\
        );

    \I__1628\ : InMux
    port map (
            O => \N__8908\,
            I => \N__8895\
        );

    \I__1627\ : InMux
    port map (
            O => \N__8905\,
            I => \N__8895\
        );

    \I__1626\ : InMux
    port map (
            O => \N__8904\,
            I => \N__8891\
        );

    \I__1625\ : InMux
    port map (
            O => \N__8903\,
            I => \N__8888\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__8900\,
            I => \N__8883\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__8895\,
            I => \N__8883\
        );

    \I__1622\ : InMux
    port map (
            O => \N__8894\,
            I => \N__8880\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__8891\,
            I => \DUT.uart_inst0.tx_countdown_3_4\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__8888\,
            I => \DUT.uart_inst0.tx_countdown_3_4\
        );

    \I__1619\ : Odrv4
    port map (
            O => \N__8883\,
            I => \DUT.uart_inst0.tx_countdown_3_4\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__8880\,
            I => \DUT.uart_inst0.tx_countdown_3_4\
        );

    \I__1617\ : InMux
    port map (
            O => \N__8871\,
            I => \N__8863\
        );

    \I__1616\ : InMux
    port map (
            O => \N__8870\,
            I => \N__8858\
        );

    \I__1615\ : InMux
    port map (
            O => \N__8869\,
            I => \N__8858\
        );

    \I__1614\ : CascadeMux
    port map (
            O => \N__8868\,
            I => \N__8855\
        );

    \I__1613\ : InMux
    port map (
            O => \N__8867\,
            I => \N__8852\
        );

    \I__1612\ : InMux
    port map (
            O => \N__8866\,
            I => \N__8849\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__8863\,
            I => \N__8844\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__8858\,
            I => \N__8844\
        );

    \I__1609\ : InMux
    port map (
            O => \N__8855\,
            I => \N__8841\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__8852\,
            I => \DUT.uart_inst0.tx_countdown_3_1\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__8849\,
            I => \DUT.uart_inst0.tx_countdown_3_1\
        );

    \I__1606\ : Odrv4
    port map (
            O => \N__8844\,
            I => \DUT.uart_inst0.tx_countdown_3_1\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__8841\,
            I => \DUT.uart_inst0.tx_countdown_3_1\
        );

    \I__1604\ : InMux
    port map (
            O => \N__8832\,
            I => \N__8826\
        );

    \I__1603\ : InMux
    port map (
            O => \N__8831\,
            I => \N__8821\
        );

    \I__1602\ : InMux
    port map (
            O => \N__8830\,
            I => \N__8821\
        );

    \I__1601\ : InMux
    port map (
            O => \N__8829\,
            I => \N__8817\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__8826\,
            I => \N__8814\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__8821\,
            I => \N__8811\
        );

    \I__1598\ : InMux
    port map (
            O => \N__8820\,
            I => \N__8808\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__8817\,
            I => \DUT.uart_inst0.tx_countdown_3_3\
        );

    \I__1596\ : Odrv4
    port map (
            O => \N__8814\,
            I => \DUT.uart_inst0.tx_countdown_3_3\
        );

    \I__1595\ : Odrv4
    port map (
            O => \N__8811\,
            I => \DUT.uart_inst0.tx_countdown_3_3\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__8808\,
            I => \DUT.uart_inst0.tx_countdown_3_3\
        );

    \I__1593\ : InMux
    port map (
            O => \N__8799\,
            I => \N__8795\
        );

    \I__1592\ : InMux
    port map (
            O => \N__8798\,
            I => \N__8790\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__8795\,
            I => \N__8786\
        );

    \I__1590\ : InMux
    port map (
            O => \N__8794\,
            I => \N__8781\
        );

    \I__1589\ : InMux
    port map (
            O => \N__8793\,
            I => \N__8781\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__8790\,
            I => \N__8778\
        );

    \I__1587\ : InMux
    port map (
            O => \N__8789\,
            I => \N__8775\
        );

    \I__1586\ : Span4Mux_h
    port map (
            O => \N__8786\,
            I => \N__8772\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__8781\,
            I => \N__8769\
        );

    \I__1584\ : Span4Mux_v
    port map (
            O => \N__8778\,
            I => \N__8764\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__8775\,
            I => \N__8764\
        );

    \I__1582\ : Odrv4
    port map (
            O => \N__8772\,
            I => \DUT.uart_inst0.tx_countdown_3_0\
        );

    \I__1581\ : Odrv4
    port map (
            O => \N__8769\,
            I => \DUT.uart_inst0.tx_countdown_3_0\
        );

    \I__1580\ : Odrv4
    port map (
            O => \N__8764\,
            I => \DUT.uart_inst0.tx_countdown_3_0\
        );

    \I__1579\ : CascadeMux
    port map (
            O => \N__8757\,
            I => \DUT.uart_inst0.N_77_cascade_\
        );

    \I__1578\ : CascadeMux
    port map (
            O => \N__8754\,
            I => \N__8750\
        );

    \I__1577\ : InMux
    port map (
            O => \N__8753\,
            I => \N__8744\
        );

    \I__1576\ : InMux
    port map (
            O => \N__8750\,
            I => \N__8739\
        );

    \I__1575\ : InMux
    port map (
            O => \N__8749\,
            I => \N__8739\
        );

    \I__1574\ : InMux
    port map (
            O => \N__8748\,
            I => \N__8735\
        );

    \I__1573\ : InMux
    port map (
            O => \N__8747\,
            I => \N__8732\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__8744\,
            I => \N__8729\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__8739\,
            I => \N__8726\
        );

    \I__1570\ : InMux
    port map (
            O => \N__8738\,
            I => \N__8723\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__8735\,
            I => \DUT.uart_inst0.tx_countdown_3_5\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__8732\,
            I => \DUT.uart_inst0.tx_countdown_3_5\
        );

    \I__1567\ : Odrv4
    port map (
            O => \N__8729\,
            I => \DUT.uart_inst0.tx_countdown_3_5\
        );

    \I__1566\ : Odrv4
    port map (
            O => \N__8726\,
            I => \DUT.uart_inst0.tx_countdown_3_5\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__8723\,
            I => \DUT.uart_inst0.tx_countdown_3_5\
        );

    \I__1564\ : CascadeMux
    port map (
            O => \N__8712\,
            I => \DUT.uart_inst0.tx_state_RNI9DTT5Z0Z_0_cascade_\
        );

    \I__1563\ : InMux
    port map (
            O => \N__8709\,
            I => \N__8706\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__8706\,
            I => \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIMJ5ECZ0\
        );

    \I__1561\ : CascadeMux
    port map (
            O => \N__8703\,
            I => \DUT.uart_inst0.N_99_cascade_\
        );

    \I__1560\ : InMux
    port map (
            O => \N__8700\,
            I => \N__8697\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__8697\,
            I => \DUT.uart_inst0.un1_tx_bits_remaining_cry_0_c_RNOZ0\
        );

    \I__1558\ : InMux
    port map (
            O => \N__8694\,
            I => \N__8683\
        );

    \I__1557\ : InMux
    port map (
            O => \N__8693\,
            I => \N__8683\
        );

    \I__1556\ : InMux
    port map (
            O => \N__8692\,
            I => \N__8680\
        );

    \I__1555\ : InMux
    port map (
            O => \N__8691\,
            I => \N__8675\
        );

    \I__1554\ : InMux
    port map (
            O => \N__8690\,
            I => \N__8675\
        );

    \I__1553\ : InMux
    port map (
            O => \N__8689\,
            I => \N__8670\
        );

    \I__1552\ : InMux
    port map (
            O => \N__8688\,
            I => \N__8670\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__8683\,
            I => \N__8667\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__8680\,
            I => \DUT.tx_state_1\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__8675\,
            I => \DUT.tx_state_1\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__8670\,
            I => \DUT.tx_state_1\
        );

    \I__1547\ : Odrv4
    port map (
            O => \N__8667\,
            I => \DUT.tx_state_1\
        );

    \I__1546\ : CascadeMux
    port map (
            O => \N__8658\,
            I => \N__8655\
        );

    \I__1545\ : InMux
    port map (
            O => \N__8655\,
            I => \N__8652\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__8652\,
            I => \N__8649\
        );

    \I__1543\ : Span4Mux_v
    port map (
            O => \N__8649\,
            I => \N__8646\
        );

    \I__1542\ : Odrv4
    port map (
            O => \N__8646\,
            I => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_3\
        );

    \I__1541\ : CascadeMux
    port map (
            O => \N__8643\,
            I => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_3_cascade_\
        );

    \I__1540\ : IoInMux
    port map (
            O => \N__8640\,
            I => \N__8637\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__8637\,
            I => \N__8634\
        );

    \I__1538\ : Span4Mux_s2_v
    port map (
            O => \N__8634\,
            I => \N__8631\
        );

    \I__1537\ : Span4Mux_v
    port map (
            O => \N__8631\,
            I => \N__8628\
        );

    \I__1536\ : Span4Mux_v
    port map (
            O => \N__8628\,
            I => \N__8624\
        );

    \I__1535\ : CascadeMux
    port map (
            O => \N__8627\,
            I => \N__8621\
        );

    \I__1534\ : Span4Mux_h
    port map (
            O => \N__8624\,
            I => \N__8617\
        );

    \I__1533\ : InMux
    port map (
            O => \N__8621\,
            I => \N__8614\
        );

    \I__1532\ : InMux
    port map (
            O => \N__8620\,
            I => \N__8611\
        );

    \I__1531\ : Odrv4
    port map (
            O => \N__8617\,
            I => \P1A7_c\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__8614\,
            I => \P1A7_c\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__8611\,
            I => \P1A7_c\
        );

    \I__1528\ : InMux
    port map (
            O => \N__8604\,
            I => \N__8601\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__8601\,
            I => \DUT.uart_inst0.N_112\
        );

    \I__1526\ : CascadeMux
    port map (
            O => \N__8598\,
            I => \DUT.uart_inst0.tx_out_6_iv_0_a3_1_1_cascade_\
        );

    \I__1525\ : CascadeMux
    port map (
            O => \N__8595\,
            I => \DUT.uart_inst0.tx_out_6_iv_0_a3_1_sx_cascade_\
        );

    \I__1524\ : InMux
    port map (
            O => \N__8592\,
            I => \N__8589\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__8589\,
            I => \DUT.uart_inst0.N_113\
        );

    \I__1522\ : CascadeMux
    port map (
            O => \N__8586\,
            I => \N__8583\
        );

    \I__1521\ : InMux
    port map (
            O => \N__8583\,
            I => \N__8580\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__8580\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_3\
        );

    \I__1519\ : InMux
    port map (
            O => \N__8577\,
            I => \N__8574\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__8574\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_3\
        );

    \I__1517\ : CascadeMux
    port map (
            O => \N__8571\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_\
        );

    \I__1516\ : InMux
    port map (
            O => \N__8568\,
            I => \N__8565\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__8565\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6\
        );

    \I__1514\ : InMux
    port map (
            O => \N__8562\,
            I => \N__8559\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__8559\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_6\
        );

    \I__1512\ : InMux
    port map (
            O => \N__8556\,
            I => \N__8553\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__8553\,
            I => \N__8550\
        );

    \I__1510\ : Odrv12
    port map (
            O => \N__8550\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_3\
        );

    \I__1509\ : InMux
    port map (
            O => \N__8547\,
            I => \N__8544\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__8544\,
            I => \N__8541\
        );

    \I__1507\ : Odrv4
    port map (
            O => \N__8541\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_5\
        );

    \I__1506\ : CascadeMux
    port map (
            O => \N__8538\,
            I => \N__8528\
        );

    \I__1505\ : CascadeMux
    port map (
            O => \N__8537\,
            I => \N__8525\
        );

    \I__1504\ : CascadeMux
    port map (
            O => \N__8536\,
            I => \N__8521\
        );

    \I__1503\ : CascadeMux
    port map (
            O => \N__8535\,
            I => \N__8517\
        );

    \I__1502\ : CascadeMux
    port map (
            O => \N__8534\,
            I => \N__8513\
        );

    \I__1501\ : CascadeMux
    port map (
            O => \N__8533\,
            I => \N__8509\
        );

    \I__1500\ : CascadeMux
    port map (
            O => \N__8532\,
            I => \N__8505\
        );

    \I__1499\ : InMux
    port map (
            O => \N__8531\,
            I => \N__8484\
        );

    \I__1498\ : InMux
    port map (
            O => \N__8528\,
            I => \N__8484\
        );

    \I__1497\ : InMux
    port map (
            O => \N__8525\,
            I => \N__8484\
        );

    \I__1496\ : InMux
    port map (
            O => \N__8524\,
            I => \N__8484\
        );

    \I__1495\ : InMux
    port map (
            O => \N__8521\,
            I => \N__8484\
        );

    \I__1494\ : InMux
    port map (
            O => \N__8520\,
            I => \N__8484\
        );

    \I__1493\ : InMux
    port map (
            O => \N__8517\,
            I => \N__8469\
        );

    \I__1492\ : InMux
    port map (
            O => \N__8516\,
            I => \N__8469\
        );

    \I__1491\ : InMux
    port map (
            O => \N__8513\,
            I => \N__8469\
        );

    \I__1490\ : InMux
    port map (
            O => \N__8512\,
            I => \N__8469\
        );

    \I__1489\ : InMux
    port map (
            O => \N__8509\,
            I => \N__8469\
        );

    \I__1488\ : InMux
    port map (
            O => \N__8508\,
            I => \N__8469\
        );

    \I__1487\ : InMux
    port map (
            O => \N__8505\,
            I => \N__8469\
        );

    \I__1486\ : CascadeMux
    port map (
            O => \N__8504\,
            I => \N__8464\
        );

    \I__1485\ : CascadeMux
    port map (
            O => \N__8503\,
            I => \N__8460\
        );

    \I__1484\ : CascadeMux
    port map (
            O => \N__8502\,
            I => \N__8456\
        );

    \I__1483\ : CascadeMux
    port map (
            O => \N__8501\,
            I => \N__8452\
        );

    \I__1482\ : CascadeMux
    port map (
            O => \N__8500\,
            I => \N__8447\
        );

    \I__1481\ : CascadeMux
    port map (
            O => \N__8499\,
            I => \N__8444\
        );

    \I__1480\ : CascadeMux
    port map (
            O => \N__8498\,
            I => \N__8441\
        );

    \I__1479\ : CascadeMux
    port map (
            O => \N__8497\,
            I => \N__8436\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__8484\,
            I => \N__8430\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__8469\,
            I => \N__8430\
        );

    \I__1476\ : InMux
    port map (
            O => \N__8468\,
            I => \N__8427\
        );

    \I__1475\ : InMux
    port map (
            O => \N__8467\,
            I => \N__8410\
        );

    \I__1474\ : InMux
    port map (
            O => \N__8464\,
            I => \N__8410\
        );

    \I__1473\ : InMux
    port map (
            O => \N__8463\,
            I => \N__8410\
        );

    \I__1472\ : InMux
    port map (
            O => \N__8460\,
            I => \N__8410\
        );

    \I__1471\ : InMux
    port map (
            O => \N__8459\,
            I => \N__8410\
        );

    \I__1470\ : InMux
    port map (
            O => \N__8456\,
            I => \N__8410\
        );

    \I__1469\ : InMux
    port map (
            O => \N__8455\,
            I => \N__8410\
        );

    \I__1468\ : InMux
    port map (
            O => \N__8452\,
            I => \N__8410\
        );

    \I__1467\ : InMux
    port map (
            O => \N__8451\,
            I => \N__8407\
        );

    \I__1466\ : InMux
    port map (
            O => \N__8450\,
            I => \N__8392\
        );

    \I__1465\ : InMux
    port map (
            O => \N__8447\,
            I => \N__8392\
        );

    \I__1464\ : InMux
    port map (
            O => \N__8444\,
            I => \N__8392\
        );

    \I__1463\ : InMux
    port map (
            O => \N__8441\,
            I => \N__8392\
        );

    \I__1462\ : InMux
    port map (
            O => \N__8440\,
            I => \N__8392\
        );

    \I__1461\ : InMux
    port map (
            O => \N__8439\,
            I => \N__8392\
        );

    \I__1460\ : InMux
    port map (
            O => \N__8436\,
            I => \N__8392\
        );

    \I__1459\ : InMux
    port map (
            O => \N__8435\,
            I => \N__8389\
        );

    \I__1458\ : Span4Mux_v
    port map (
            O => \N__8430\,
            I => \N__8381\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__8427\,
            I => \N__8381\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__8410\,
            I => \N__8381\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__8407\,
            I => \N__8376\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__8392\,
            I => \N__8376\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__8389\,
            I => \N__8373\
        );

    \I__1452\ : InMux
    port map (
            O => \N__8388\,
            I => \N__8370\
        );

    \I__1451\ : Span4Mux_v
    port map (
            O => \N__8381\,
            I => \N__8365\
        );

    \I__1450\ : Span4Mux_v
    port map (
            O => \N__8376\,
            I => \N__8365\
        );

    \I__1449\ : Span4Mux_v
    port map (
            O => \N__8373\,
            I => \N__8362\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__8370\,
            I => \N__8359\
        );

    \I__1447\ : Odrv4
    port map (
            O => \N__8365\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1446\ : Odrv4
    port map (
            O => \N__8362\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1445\ : Odrv12
    port map (
            O => \N__8359\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1444\ : CascadeMux
    port map (
            O => \N__8352\,
            I => \N__8345\
        );

    \I__1443\ : CascadeMux
    port map (
            O => \N__8351\,
            I => \N__8342\
        );

    \I__1442\ : InMux
    port map (
            O => \N__8350\,
            I => \N__8337\
        );

    \I__1441\ : CascadeMux
    port map (
            O => \N__8349\,
            I => \N__8330\
        );

    \I__1440\ : InMux
    port map (
            O => \N__8348\,
            I => \N__8322\
        );

    \I__1439\ : InMux
    port map (
            O => \N__8345\,
            I => \N__8322\
        );

    \I__1438\ : InMux
    port map (
            O => \N__8342\,
            I => \N__8322\
        );

    \I__1437\ : CascadeMux
    port map (
            O => \N__8341\,
            I => \N__8312\
        );

    \I__1436\ : InMux
    port map (
            O => \N__8340\,
            I => \N__8309\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__8337\,
            I => \N__8306\
        );

    \I__1434\ : InMux
    port map (
            O => \N__8336\,
            I => \N__8303\
        );

    \I__1433\ : InMux
    port map (
            O => \N__8335\,
            I => \N__8298\
        );

    \I__1432\ : InMux
    port map (
            O => \N__8334\,
            I => \N__8293\
        );

    \I__1431\ : InMux
    port map (
            O => \N__8333\,
            I => \N__8293\
        );

    \I__1430\ : InMux
    port map (
            O => \N__8330\,
            I => \N__8288\
        );

    \I__1429\ : InMux
    port map (
            O => \N__8329\,
            I => \N__8288\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__8322\,
            I => \N__8275\
        );

    \I__1427\ : InMux
    port map (
            O => \N__8321\,
            I => \N__8270\
        );

    \I__1426\ : InMux
    port map (
            O => \N__8320\,
            I => \N__8270\
        );

    \I__1425\ : InMux
    port map (
            O => \N__8319\,
            I => \N__8265\
        );

    \I__1424\ : InMux
    port map (
            O => \N__8318\,
            I => \N__8265\
        );

    \I__1423\ : InMux
    port map (
            O => \N__8317\,
            I => \N__8256\
        );

    \I__1422\ : InMux
    port map (
            O => \N__8316\,
            I => \N__8256\
        );

    \I__1421\ : InMux
    port map (
            O => \N__8315\,
            I => \N__8256\
        );

    \I__1420\ : InMux
    port map (
            O => \N__8312\,
            I => \N__8256\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__8309\,
            I => \N__8253\
        );

    \I__1418\ : Span4Mux_v
    port map (
            O => \N__8306\,
            I => \N__8248\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__8303\,
            I => \N__8248\
        );

    \I__1416\ : InMux
    port map (
            O => \N__8302\,
            I => \N__8245\
        );

    \I__1415\ : InMux
    port map (
            O => \N__8301\,
            I => \N__8242\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__8298\,
            I => \N__8235\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__8293\,
            I => \N__8235\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__8288\,
            I => \N__8235\
        );

    \I__1411\ : InMux
    port map (
            O => \N__8287\,
            I => \N__8220\
        );

    \I__1410\ : InMux
    port map (
            O => \N__8286\,
            I => \N__8220\
        );

    \I__1409\ : InMux
    port map (
            O => \N__8285\,
            I => \N__8220\
        );

    \I__1408\ : InMux
    port map (
            O => \N__8284\,
            I => \N__8220\
        );

    \I__1407\ : InMux
    port map (
            O => \N__8283\,
            I => \N__8220\
        );

    \I__1406\ : InMux
    port map (
            O => \N__8282\,
            I => \N__8220\
        );

    \I__1405\ : InMux
    port map (
            O => \N__8281\,
            I => \N__8220\
        );

    \I__1404\ : InMux
    port map (
            O => \N__8280\,
            I => \N__8217\
        );

    \I__1403\ : InMux
    port map (
            O => \N__8279\,
            I => \N__8212\
        );

    \I__1402\ : InMux
    port map (
            O => \N__8278\,
            I => \N__8212\
        );

    \I__1401\ : Span4Mux_v
    port map (
            O => \N__8275\,
            I => \N__8207\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__8270\,
            I => \N__8207\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__8265\,
            I => \N__8202\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__8256\,
            I => \N__8202\
        );

    \I__1397\ : Span4Mux_v
    port map (
            O => \N__8253\,
            I => \N__8199\
        );

    \I__1396\ : Span4Mux_v
    port map (
            O => \N__8248\,
            I => \N__8194\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__8245\,
            I => \N__8194\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__8242\,
            I => \N__8183\
        );

    \I__1393\ : Span4Mux_v
    port map (
            O => \N__8235\,
            I => \N__8183\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__8220\,
            I => \N__8183\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__8217\,
            I => \N__8183\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__8212\,
            I => \N__8183\
        );

    \I__1389\ : Span4Mux_v
    port map (
            O => \N__8207\,
            I => \N__8178\
        );

    \I__1388\ : Span4Mux_v
    port map (
            O => \N__8202\,
            I => \N__8178\
        );

    \I__1387\ : Span4Mux_h
    port map (
            O => \N__8199\,
            I => \N__8171\
        );

    \I__1386\ : Span4Mux_v
    port map (
            O => \N__8194\,
            I => \N__8171\
        );

    \I__1385\ : Span4Mux_v
    port map (
            O => \N__8183\,
            I => \N__8171\
        );

    \I__1384\ : Sp12to4
    port map (
            O => \N__8178\,
            I => \N__8166\
        );

    \I__1383\ : Sp12to4
    port map (
            O => \N__8171\,
            I => \N__8166\
        );

    \I__1382\ : Span12Mux_h
    port map (
            O => \N__8166\,
            I => \N__8163\
        );

    \I__1381\ : Odrv12
    port map (
            O => \N__8163\,
            I => \P1A1_c\
        );

    \I__1380\ : InMux
    port map (
            O => \N__8160\,
            I => \N__8157\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__8157\,
            I => \N__8154\
        );

    \I__1378\ : Span4Mux_h
    port map (
            O => \N__8154\,
            I => \N__8151\
        );

    \I__1377\ : Odrv4
    port map (
            O => \N__8151\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO\
        );

    \I__1376\ : CascadeMux
    port map (
            O => \N__8148\,
            I => \N__8141\
        );

    \I__1375\ : CascadeMux
    port map (
            O => \N__8147\,
            I => \N__8134\
        );

    \I__1374\ : CascadeMux
    port map (
            O => \N__8146\,
            I => \N__8131\
        );

    \I__1373\ : CascadeMux
    port map (
            O => \N__8145\,
            I => \N__8128\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__8144\,
            I => \N__8125\
        );

    \I__1371\ : InMux
    port map (
            O => \N__8141\,
            I => \N__8116\
        );

    \I__1370\ : CascadeMux
    port map (
            O => \N__8140\,
            I => \N__8111\
        );

    \I__1369\ : InMux
    port map (
            O => \N__8139\,
            I => \N__8096\
        );

    \I__1368\ : InMux
    port map (
            O => \N__8138\,
            I => \N__8096\
        );

    \I__1367\ : InMux
    port map (
            O => \N__8137\,
            I => \N__8096\
        );

    \I__1366\ : InMux
    port map (
            O => \N__8134\,
            I => \N__8096\
        );

    \I__1365\ : InMux
    port map (
            O => \N__8131\,
            I => \N__8096\
        );

    \I__1364\ : InMux
    port map (
            O => \N__8128\,
            I => \N__8096\
        );

    \I__1363\ : InMux
    port map (
            O => \N__8125\,
            I => \N__8096\
        );

    \I__1362\ : InMux
    port map (
            O => \N__8124\,
            I => \N__8091\
        );

    \I__1361\ : InMux
    port map (
            O => \N__8123\,
            I => \N__8091\
        );

    \I__1360\ : CascadeMux
    port map (
            O => \N__8122\,
            I => \N__8088\
        );

    \I__1359\ : CascadeMux
    port map (
            O => \N__8121\,
            I => \N__8085\
        );

    \I__1358\ : CascadeMux
    port map (
            O => \N__8120\,
            I => \N__8082\
        );

    \I__1357\ : CascadeMux
    port map (
            O => \N__8119\,
            I => \N__8079\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__8116\,
            I => \N__8074\
        );

    \I__1355\ : InMux
    port map (
            O => \N__8115\,
            I => \N__8071\
        );

    \I__1354\ : InMux
    port map (
            O => \N__8114\,
            I => \N__8065\
        );

    \I__1353\ : InMux
    port map (
            O => \N__8111\,
            I => \N__8065\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__8096\,
            I => \N__8060\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__8091\,
            I => \N__8060\
        );

    \I__1350\ : InMux
    port map (
            O => \N__8088\,
            I => \N__8047\
        );

    \I__1349\ : InMux
    port map (
            O => \N__8085\,
            I => \N__8047\
        );

    \I__1348\ : InMux
    port map (
            O => \N__8082\,
            I => \N__8047\
        );

    \I__1347\ : InMux
    port map (
            O => \N__8079\,
            I => \N__8047\
        );

    \I__1346\ : InMux
    port map (
            O => \N__8078\,
            I => \N__8047\
        );

    \I__1345\ : InMux
    port map (
            O => \N__8077\,
            I => \N__8047\
        );

    \I__1344\ : Span4Mux_v
    port map (
            O => \N__8074\,
            I => \N__8042\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__8071\,
            I => \N__8042\
        );

    \I__1342\ : InMux
    port map (
            O => \N__8070\,
            I => \N__8037\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__8065\,
            I => \N__8034\
        );

    \I__1340\ : Span4Mux_v
    port map (
            O => \N__8060\,
            I => \N__8031\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__8047\,
            I => \N__8026\
        );

    \I__1338\ : Span4Mux_h
    port map (
            O => \N__8042\,
            I => \N__8026\
        );

    \I__1337\ : InMux
    port map (
            O => \N__8041\,
            I => \N__8021\
        );

    \I__1336\ : InMux
    port map (
            O => \N__8040\,
            I => \N__8021\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__8037\,
            I => \DUT.uart_inst0.recv_stateZ0Z_0\
        );

    \I__1334\ : Odrv12
    port map (
            O => \N__8034\,
            I => \DUT.uart_inst0.recv_stateZ0Z_0\
        );

    \I__1333\ : Odrv4
    port map (
            O => \N__8031\,
            I => \DUT.uart_inst0.recv_stateZ0Z_0\
        );

    \I__1332\ : Odrv4
    port map (
            O => \N__8026\,
            I => \DUT.uart_inst0.recv_stateZ0Z_0\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__8021\,
            I => \DUT.uart_inst0.recv_stateZ0Z_0\
        );

    \I__1330\ : CascadeMux
    port map (
            O => \N__8010\,
            I => \N__8006\
        );

    \I__1329\ : CascadeMux
    port map (
            O => \N__8009\,
            I => \N__8003\
        );

    \I__1328\ : InMux
    port map (
            O => \N__8006\,
            I => \N__7999\
        );

    \I__1327\ : InMux
    port map (
            O => \N__8003\,
            I => \N__7996\
        );

    \I__1326\ : InMux
    port map (
            O => \N__8002\,
            I => \N__7993\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__7999\,
            I => \N__7988\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__7996\,
            I => \N__7988\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__7993\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_4\
        );

    \I__1322\ : Odrv12
    port map (
            O => \N__7988\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_4\
        );

    \I__1321\ : CascadeMux
    port map (
            O => \N__7983\,
            I => \N__7980\
        );

    \I__1320\ : InMux
    port map (
            O => \N__7980\,
            I => \N__7977\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__7977\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_6\
        );

    \I__1318\ : CascadeMux
    port map (
            O => \N__7974\,
            I => \N__7971\
        );

    \I__1317\ : InMux
    port map (
            O => \N__7971\,
            I => \N__7968\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__7968\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_7\
        );

    \I__1315\ : CEMux
    port map (
            O => \N__7965\,
            I => \N__7962\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__7962\,
            I => \N__7959\
        );

    \I__1313\ : Span4Mux_h
    port map (
            O => \N__7959\,
            I => \N__7955\
        );

    \I__1312\ : InMux
    port map (
            O => \N__7958\,
            I => \N__7952\
        );

    \I__1311\ : Odrv4
    port map (
            O => \N__7955\,
            I => \DUT.fifo_rx_inst.rFifoData_awe1\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__7952\,
            I => \DUT.fifo_rx_inst.rFifoData_awe1\
        );

    \I__1309\ : InMux
    port map (
            O => \N__7947\,
            I => \N__7944\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__7944\,
            I => \N__7941\
        );

    \I__1307\ : Odrv4
    port map (
            O => \N__7941\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_4\
        );

    \I__1306\ : InMux
    port map (
            O => \N__7938\,
            I => \N__7935\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__7935\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_4\
        );

    \I__1304\ : CascadeMux
    port map (
            O => \N__7932\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4_cascade_\
        );

    \I__1303\ : InMux
    port map (
            O => \N__7929\,
            I => \N__7926\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__7926\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_5\
        );

    \I__1301\ : CascadeMux
    port map (
            O => \N__7923\,
            I => \N__7920\
        );

    \I__1300\ : InMux
    port map (
            O => \N__7920\,
            I => \N__7917\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__7917\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_5\
        );

    \I__1298\ : InMux
    port map (
            O => \N__7914\,
            I => \N__7911\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__7911\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5\
        );

    \I__1296\ : InMux
    port map (
            O => \N__7908\,
            I => \N__7905\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__7905\,
            I => \N_100_i\
        );

    \I__1294\ : InMux
    port map (
            O => \N__7902\,
            I => \N__7899\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__7899\,
            I => \DUT.fifo_rx_inst.rTxByte_52_1\
        );

    \I__1292\ : CascadeMux
    port map (
            O => \N__7896\,
            I => \DUT.fifo_rx_inst.rTxByte_52_0_cascade_\
        );

    \I__1291\ : InMux
    port map (
            O => \N__7893\,
            I => \N__7886\
        );

    \I__1290\ : InMux
    port map (
            O => \N__7892\,
            I => \N__7886\
        );

    \I__1289\ : InMux
    port map (
            O => \N__7891\,
            I => \N__7883\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__7886\,
            I => \N__7880\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__7883\,
            I => \N__7875\
        );

    \I__1286\ : Span4Mux_v
    port map (
            O => \N__7880\,
            I => \N__7875\
        );

    \I__1285\ : Odrv4
    port map (
            O => \N__7875\,
            I => \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1Z0Z_0\
        );

    \I__1284\ : CascadeMux
    port map (
            O => \N__7872\,
            I => \N__7869\
        );

    \I__1283\ : InMux
    port map (
            O => \N__7869\,
            I => \N__7866\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__7866\,
            I => \N__7863\
        );

    \I__1281\ : Odrv4
    port map (
            O => \N__7863\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_2\
        );

    \I__1280\ : CascadeMux
    port map (
            O => \N__7860\,
            I => \N__7857\
        );

    \I__1279\ : InMux
    port map (
            O => \N__7857\,
            I => \N__7854\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__7854\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_1\
        );

    \I__1277\ : InMux
    port map (
            O => \N__7851\,
            I => \N__7848\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__7848\,
            I => \N__7845\
        );

    \I__1275\ : Odrv4
    port map (
            O => \N__7845\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_2\
        );

    \I__1274\ : InMux
    port map (
            O => \N__7842\,
            I => \N__7839\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__7839\,
            I => \DUT.uart_inst0.tx_countdown_3_axb_5\
        );

    \I__1272\ : InMux
    port map (
            O => \N__7836\,
            I => \DUT.uart_inst0.tx_countdown_3_cry_4\
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__7833\,
            I => \N__7829\
        );

    \I__1270\ : CascadeMux
    port map (
            O => \N__7832\,
            I => \N__7826\
        );

    \I__1269\ : InMux
    port map (
            O => \N__7829\,
            I => \N__7823\
        );

    \I__1268\ : InMux
    port map (
            O => \N__7826\,
            I => \N__7820\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__7823\,
            I => \N__7817\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__7820\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__1265\ : Odrv4
    port map (
            O => \N__7817\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__1264\ : InMux
    port map (
            O => \N__7812\,
            I => \N__7809\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__7809\,
            I => \DUT.uart_inst0.tx_countdown_RNI4K692Z0Z_1\
        );

    \I__1262\ : InMux
    port map (
            O => \N__7806\,
            I => \N__7795\
        );

    \I__1261\ : InMux
    port map (
            O => \N__7805\,
            I => \N__7795\
        );

    \I__1260\ : InMux
    port map (
            O => \N__7804\,
            I => \N__7790\
        );

    \I__1259\ : InMux
    port map (
            O => \N__7803\,
            I => \N__7790\
        );

    \I__1258\ : InMux
    port map (
            O => \N__7802\,
            I => \N__7783\
        );

    \I__1257\ : InMux
    port map (
            O => \N__7801\,
            I => \N__7783\
        );

    \I__1256\ : InMux
    port map (
            O => \N__7800\,
            I => \N__7783\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__7795\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_10\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__7790\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_10\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__7783\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_10\
        );

    \I__1252\ : CascadeMux
    port map (
            O => \N__7776\,
            I => \N__7772\
        );

    \I__1251\ : InMux
    port map (
            O => \N__7775\,
            I => \N__7769\
        );

    \I__1250\ : InMux
    port map (
            O => \N__7772\,
            I => \N__7766\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__7769\,
            I => \DUT.uart_inst0.tx_countdownZ1Z_3\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__7766\,
            I => \DUT.uart_inst0.tx_countdownZ1Z_3\
        );

    \I__1247\ : InMux
    port map (
            O => \N__7761\,
            I => \N__7756\
        );

    \I__1246\ : CascadeMux
    port map (
            O => \N__7760\,
            I => \N__7752\
        );

    \I__1245\ : CascadeMux
    port map (
            O => \N__7759\,
            I => \N__7748\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__7756\,
            I => \N__7743\
        );

    \I__1243\ : InMux
    port map (
            O => \N__7755\,
            I => \N__7740\
        );

    \I__1242\ : InMux
    port map (
            O => \N__7752\,
            I => \N__7735\
        );

    \I__1241\ : InMux
    port map (
            O => \N__7751\,
            I => \N__7735\
        );

    \I__1240\ : InMux
    port map (
            O => \N__7748\,
            I => \N__7728\
        );

    \I__1239\ : InMux
    port map (
            O => \N__7747\,
            I => \N__7728\
        );

    \I__1238\ : InMux
    port map (
            O => \N__7746\,
            I => \N__7728\
        );

    \I__1237\ : Odrv12
    port map (
            O => \N__7743\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_8\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__7740\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_8\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__7735\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_8\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__7728\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_8\
        );

    \I__1233\ : InMux
    port map (
            O => \N__7719\,
            I => \N__7710\
        );

    \I__1232\ : InMux
    port map (
            O => \N__7718\,
            I => \N__7705\
        );

    \I__1231\ : InMux
    port map (
            O => \N__7717\,
            I => \N__7705\
        );

    \I__1230\ : InMux
    port map (
            O => \N__7716\,
            I => \N__7696\
        );

    \I__1229\ : InMux
    port map (
            O => \N__7715\,
            I => \N__7696\
        );

    \I__1228\ : InMux
    port map (
            O => \N__7714\,
            I => \N__7696\
        );

    \I__1227\ : InMux
    port map (
            O => \N__7713\,
            I => \N__7696\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__7710\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_9\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__7705\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_9\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__7696\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_9\
        );

    \I__1223\ : InMux
    port map (
            O => \N__7689\,
            I => \N__7686\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__7686\,
            I => \DUT.uart_inst0.tx_countdown_RNI6M692Z0Z_3\
        );

    \I__1221\ : InMux
    port map (
            O => \N__7683\,
            I => \DUT.uart_inst0.un1_tx_bits_remaining_cry_0\
        );

    \I__1220\ : InMux
    port map (
            O => \N__7680\,
            I => \DUT.uart_inst0.un1_tx_bits_remaining_cry_1\
        );

    \I__1219\ : InMux
    port map (
            O => \N__7677\,
            I => \DUT.uart_inst0.un1_tx_bits_remaining_cry_2\
        );

    \I__1218\ : IoInMux
    port map (
            O => \N__7674\,
            I => \N__7671\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__7671\,
            I => \N__7668\
        );

    \I__1216\ : IoSpan4Mux
    port map (
            O => \N__7668\,
            I => \N__7664\
        );

    \I__1215\ : IoInMux
    port map (
            O => \N__7667\,
            I => \N__7661\
        );

    \I__1214\ : Span4Mux_s3_v
    port map (
            O => \N__7664\,
            I => \N__7658\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__7661\,
            I => \N__7655\
        );

    \I__1212\ : Span4Mux_h
    port map (
            O => \N__7658\,
            I => \N__7650\
        );

    \I__1211\ : Span4Mux_s3_v
    port map (
            O => \N__7655\,
            I => \N__7650\
        );

    \I__1210\ : Sp12to4
    port map (
            O => \N__7650\,
            I => \N__7647\
        );

    \I__1209\ : Span12Mux_s11_h
    port map (
            O => \N__7647\,
            I => \N__7643\
        );

    \I__1208\ : InMux
    port map (
            O => \N__7646\,
            I => \N__7640\
        );

    \I__1207\ : Odrv12
    port map (
            O => \N__7643\,
            I => \P1A3_c\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__7640\,
            I => \P1A3_c\
        );

    \I__1205\ : InMux
    port map (
            O => \N__7635\,
            I => \N__7631\
        );

    \I__1204\ : InMux
    port map (
            O => \N__7634\,
            I => \N__7628\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__7631\,
            I => \DUT.uart_inst0.N_82\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__7628\,
            I => \DUT.uart_inst0.N_82\
        );

    \I__1201\ : InMux
    port map (
            O => \N__7623\,
            I => \N__7620\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__7620\,
            I => \DUT.uart_inst0.tx_countdown_3_cry_0_c_RNOZ0\
        );

    \I__1199\ : CascadeMux
    port map (
            O => \N__7617\,
            I => \N__7613\
        );

    \I__1198\ : CascadeMux
    port map (
            O => \N__7616\,
            I => \N__7609\
        );

    \I__1197\ : InMux
    port map (
            O => \N__7613\,
            I => \N__7606\
        );

    \I__1196\ : InMux
    port map (
            O => \N__7612\,
            I => \N__7603\
        );

    \I__1195\ : InMux
    port map (
            O => \N__7609\,
            I => \N__7600\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__7606\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__7603\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__7600\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__1191\ : InMux
    port map (
            O => \N__7593\,
            I => \DUT.uart_inst0.tx_countdown_3_cry_0\
        );

    \I__1190\ : InMux
    port map (
            O => \N__7590\,
            I => \N__7587\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__7587\,
            I => \DUT.uart_inst0.tx_countdown_RNI5L692Z0Z_2\
        );

    \I__1188\ : InMux
    port map (
            O => \N__7584\,
            I => \N__7580\
        );

    \I__1187\ : CascadeMux
    port map (
            O => \N__7583\,
            I => \N__7577\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__7580\,
            I => \N__7574\
        );

    \I__1185\ : InMux
    port map (
            O => \N__7577\,
            I => \N__7571\
        );

    \I__1184\ : Span12Mux_v
    port map (
            O => \N__7574\,
            I => \N__7568\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__7571\,
            I => \N__7565\
        );

    \I__1182\ : Odrv12
    port map (
            O => \N__7568\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_2\
        );

    \I__1181\ : Odrv4
    port map (
            O => \N__7565\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_2\
        );

    \I__1180\ : InMux
    port map (
            O => \N__7560\,
            I => \DUT.uart_inst0.tx_countdown_3_cry_1\
        );

    \I__1179\ : InMux
    port map (
            O => \N__7557\,
            I => \DUT.uart_inst0.tx_countdown_3_cry_2\
        );

    \I__1178\ : InMux
    port map (
            O => \N__7554\,
            I => \N__7551\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__7551\,
            I => \DUT.uart_inst0.tx_countdown_RNI7N692Z0Z_4\
        );

    \I__1176\ : InMux
    port map (
            O => \N__7548\,
            I => \N__7544\
        );

    \I__1175\ : CascadeMux
    port map (
            O => \N__7547\,
            I => \N__7541\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__7544\,
            I => \N__7538\
        );

    \I__1173\ : InMux
    port map (
            O => \N__7541\,
            I => \N__7535\
        );

    \I__1172\ : Odrv4
    port map (
            O => \N__7538\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_4\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__7535\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_4\
        );

    \I__1170\ : InMux
    port map (
            O => \N__7530\,
            I => \DUT.uart_inst0.tx_countdown_3_cry_3\
        );

    \I__1169\ : CascadeMux
    port map (
            O => \N__7527\,
            I => \DUT.uart_inst0.tx_bits_remaining_RNI5UON8Z0Z_3_cascade_\
        );

    \I__1168\ : CascadeMux
    port map (
            O => \N__7524\,
            I => \DUT.uart_inst0.N_109_cascade_\
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__7521\,
            I => \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIKK41CZ0_cascade_\
        );

    \I__1166\ : InMux
    port map (
            O => \N__7518\,
            I => \N__7515\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__7515\,
            I => \DUT.uart_inst0.N_109\
        );

    \I__1164\ : InMux
    port map (
            O => \N__7512\,
            I => \N__7509\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__7509\,
            I => \DUT.uart_inst0.tx_state_ns_i_i_a3_1_0\
        );

    \I__1162\ : InMux
    port map (
            O => \N__7506\,
            I => \N__7503\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__7503\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_6\
        );

    \I__1160\ : CEMux
    port map (
            O => \N__7500\,
            I => \N__7496\
        );

    \I__1159\ : CEMux
    port map (
            O => \N__7499\,
            I => \N__7492\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__7496\,
            I => \N__7489\
        );

    \I__1157\ : CEMux
    port map (
            O => \N__7495\,
            I => \N__7486\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__7492\,
            I => \N__7483\
        );

    \I__1155\ : Span4Mux_h
    port map (
            O => \N__7489\,
            I => \N__7478\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__7486\,
            I => \N__7478\
        );

    \I__1153\ : Span4Mux_h
    port map (
            O => \N__7483\,
            I => \N__7475\
        );

    \I__1152\ : Span4Mux_h
    port map (
            O => \N__7478\,
            I => \N__7472\
        );

    \I__1151\ : Span4Mux_v
    port map (
            O => \N__7475\,
            I => \N__7469\
        );

    \I__1150\ : Span4Mux_v
    port map (
            O => \N__7472\,
            I => \N__7466\
        );

    \I__1149\ : Odrv4
    port map (
            O => \N__7469\,
            I => \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa\
        );

    \I__1148\ : Odrv4
    port map (
            O => \N__7466\,
            I => \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa\
        );

    \I__1147\ : CascadeMux
    port map (
            O => \N__7461\,
            I => \DUT.uart_inst0.g0_0_1_cascade_\
        );

    \I__1146\ : InMux
    port map (
            O => \N__7458\,
            I => \N__7450\
        );

    \I__1145\ : InMux
    port map (
            O => \N__7457\,
            I => \N__7447\
        );

    \I__1144\ : InMux
    port map (
            O => \N__7456\,
            I => \N__7440\
        );

    \I__1143\ : InMux
    port map (
            O => \N__7455\,
            I => \N__7440\
        );

    \I__1142\ : InMux
    port map (
            O => \N__7454\,
            I => \N__7440\
        );

    \I__1141\ : InMux
    port map (
            O => \N__7453\,
            I => \N__7437\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__7450\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_0\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__7447\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_0\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__7440\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_0\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__7437\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_0\
        );

    \I__1136\ : InMux
    port map (
            O => \N__7428\,
            I => \N__7424\
        );

    \I__1135\ : InMux
    port map (
            O => \N__7427\,
            I => \N__7421\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__7424\,
            I => \DUT.uart_inst0.N_62_4\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__7421\,
            I => \DUT.uart_inst0.N_62_4\
        );

    \I__1132\ : InMux
    port map (
            O => \N__7416\,
            I => \N__7407\
        );

    \I__1131\ : InMux
    port map (
            O => \N__7415\,
            I => \N__7407\
        );

    \I__1130\ : InMux
    port map (
            O => \N__7414\,
            I => \N__7403\
        );

    \I__1129\ : InMux
    port map (
            O => \N__7413\,
            I => \N__7398\
        );

    \I__1128\ : InMux
    port map (
            O => \N__7412\,
            I => \N__7398\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__7407\,
            I => \N__7395\
        );

    \I__1126\ : InMux
    port map (
            O => \N__7406\,
            I => \N__7392\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__7403\,
            I => \N__7387\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__7398\,
            I => \N__7380\
        );

    \I__1123\ : Span4Mux_h
    port map (
            O => \N__7395\,
            I => \N__7380\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__7392\,
            I => \N__7380\
        );

    \I__1121\ : InMux
    port map (
            O => \N__7391\,
            I => \N__7375\
        );

    \I__1120\ : InMux
    port map (
            O => \N__7390\,
            I => \N__7375\
        );

    \I__1119\ : Odrv12
    port map (
            O => \N__7387\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__1118\ : Odrv4
    port map (
            O => \N__7380\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__7375\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__1116\ : CascadeMux
    port map (
            O => \N__7368\,
            I => \DUT.uart_inst0.recv_state_srsts_1_2_cascade_\
        );

    \I__1115\ : InMux
    port map (
            O => \N__7365\,
            I => \N__7355\
        );

    \I__1114\ : InMux
    port map (
            O => \N__7364\,
            I => \N__7350\
        );

    \I__1113\ : InMux
    port map (
            O => \N__7363\,
            I => \N__7350\
        );

    \I__1112\ : InMux
    port map (
            O => \N__7362\,
            I => \N__7341\
        );

    \I__1111\ : InMux
    port map (
            O => \N__7361\,
            I => \N__7341\
        );

    \I__1110\ : InMux
    port map (
            O => \N__7360\,
            I => \N__7341\
        );

    \I__1109\ : InMux
    port map (
            O => \N__7359\,
            I => \N__7336\
        );

    \I__1108\ : InMux
    port map (
            O => \N__7358\,
            I => \N__7336\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__7355\,
            I => \N__7333\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__7350\,
            I => \N__7330\
        );

    \I__1105\ : InMux
    port map (
            O => \N__7349\,
            I => \N__7325\
        );

    \I__1104\ : InMux
    port map (
            O => \N__7348\,
            I => \N__7325\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__7341\,
            I => \N__7320\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__7336\,
            I => \N__7320\
        );

    \I__1101\ : Span4Mux_h
    port map (
            O => \N__7333\,
            I => \N__7317\
        );

    \I__1100\ : Odrv4
    port map (
            O => \N__7330\,
            I => \DUT.uart_inst0.N_42\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__7325\,
            I => \DUT.uart_inst0.N_42\
        );

    \I__1098\ : Odrv4
    port map (
            O => \N__7320\,
            I => \DUT.uart_inst0.N_42\
        );

    \I__1097\ : Odrv4
    port map (
            O => \N__7317\,
            I => \DUT.uart_inst0.N_42\
        );

    \I__1096\ : InMux
    port map (
            O => \N__7308\,
            I => \N__7303\
        );

    \I__1095\ : InMux
    port map (
            O => \N__7307\,
            I => \N__7300\
        );

    \I__1094\ : InMux
    port map (
            O => \N__7306\,
            I => \N__7297\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__7303\,
            I => \N__7294\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__7300\,
            I => \N__7289\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__7297\,
            I => \N__7289\
        );

    \I__1090\ : Span4Mux_h
    port map (
            O => \N__7294\,
            I => \N__7277\
        );

    \I__1089\ : Span4Mux_v
    port map (
            O => \N__7289\,
            I => \N__7274\
        );

    \I__1088\ : InMux
    port map (
            O => \N__7288\,
            I => \N__7267\
        );

    \I__1087\ : InMux
    port map (
            O => \N__7287\,
            I => \N__7267\
        );

    \I__1086\ : InMux
    port map (
            O => \N__7286\,
            I => \N__7267\
        );

    \I__1085\ : InMux
    port map (
            O => \N__7285\,
            I => \N__7262\
        );

    \I__1084\ : InMux
    port map (
            O => \N__7284\,
            I => \N__7262\
        );

    \I__1083\ : InMux
    port map (
            O => \N__7283\,
            I => \N__7253\
        );

    \I__1082\ : InMux
    port map (
            O => \N__7282\,
            I => \N__7253\
        );

    \I__1081\ : InMux
    port map (
            O => \N__7281\,
            I => \N__7253\
        );

    \I__1080\ : InMux
    port map (
            O => \N__7280\,
            I => \N__7253\
        );

    \I__1079\ : Odrv4
    port map (
            O => \N__7277\,
            I => \DUT.uart_inst0.recv_stateZ0Z_2\
        );

    \I__1078\ : Odrv4
    port map (
            O => \N__7274\,
            I => \DUT.uart_inst0.recv_stateZ0Z_2\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__7267\,
            I => \DUT.uart_inst0.recv_stateZ0Z_2\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__7262\,
            I => \DUT.uart_inst0.recv_stateZ0Z_2\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__7253\,
            I => \DUT.uart_inst0.recv_stateZ0Z_2\
        );

    \I__1074\ : InMux
    port map (
            O => \N__7242\,
            I => \N__7239\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__7239\,
            I => \DUT.uart_inst0.m5_0_0\
        );

    \I__1072\ : InMux
    port map (
            O => \N__7236\,
            I => \N__7230\
        );

    \I__1071\ : InMux
    port map (
            O => \N__7235\,
            I => \N__7230\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__7230\,
            I => \DUT.fifo_rx_inst.rFifoDataro_0\
        );

    \I__1069\ : InMux
    port map (
            O => \N__7227\,
            I => \N__7221\
        );

    \I__1068\ : InMux
    port map (
            O => \N__7226\,
            I => \N__7221\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__7221\,
            I => \DUT.fifo_rx_inst.rFifoDataro_1\
        );

    \I__1066\ : InMux
    port map (
            O => \N__7218\,
            I => \N__7215\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__7215\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_1\
        );

    \I__1064\ : InMux
    port map (
            O => \N__7212\,
            I => \N__7209\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__7209\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_7\
        );

    \I__1062\ : CascadeMux
    port map (
            O => \N__7206\,
            I => \DUT.uart_inst0.tx_countdown_3_0_cascade_\
        );

    \I__1061\ : CascadeMux
    port map (
            O => \N__7203\,
            I => \N__7200\
        );

    \I__1060\ : InMux
    port map (
            O => \N__7200\,
            I => \N__7196\
        );

    \I__1059\ : InMux
    port map (
            O => \N__7199\,
            I => \N__7193\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__7196\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_11\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__7193\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_11\
        );

    \I__1056\ : InMux
    port map (
            O => \N__7188\,
            I => \N__7184\
        );

    \I__1055\ : InMux
    port map (
            O => \N__7187\,
            I => \N__7181\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__7184\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_10\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__7181\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_10\
        );

    \I__1052\ : CascadeMux
    port map (
            O => \N__7176\,
            I => \N__7173\
        );

    \I__1051\ : InMux
    port map (
            O => \N__7173\,
            I => \N__7169\
        );

    \I__1050\ : InMux
    port map (
            O => \N__7172\,
            I => \N__7166\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__7169\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_9\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__7166\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_9\
        );

    \I__1047\ : InMux
    port map (
            O => \N__7161\,
            I => \N__7157\
        );

    \I__1046\ : InMux
    port map (
            O => \N__7160\,
            I => \N__7154\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__7157\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_8\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__7154\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_8\
        );

    \I__1043\ : InMux
    port map (
            O => \N__7149\,
            I => \N__7145\
        );

    \I__1042\ : InMux
    port map (
            O => \N__7148\,
            I => \N__7142\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__7145\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_1\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__7142\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_1\
        );

    \I__1039\ : CascadeMux
    port map (
            O => \N__7137\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_7_cascade_\
        );

    \I__1038\ : CascadeMux
    port map (
            O => \N__7134\,
            I => \N__7130\
        );

    \I__1037\ : InMux
    port map (
            O => \N__7133\,
            I => \N__7126\
        );

    \I__1036\ : InMux
    port map (
            O => \N__7130\,
            I => \N__7123\
        );

    \I__1035\ : InMux
    port map (
            O => \N__7129\,
            I => \N__7120\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__7126\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_0\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__7123\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_0\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__7120\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_0\
        );

    \I__1031\ : CascadeMux
    port map (
            O => \N__7113\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_10_cascade_\
        );

    \I__1030\ : CascadeMux
    port map (
            O => \N__7110\,
            I => \DUT.uart_inst0.tx_clk_divider_1_sqmuxa_1_0_cascade_\
        );

    \I__1029\ : SRMux
    port map (
            O => \N__7107\,
            I => \N__7103\
        );

    \I__1028\ : SRMux
    port map (
            O => \N__7106\,
            I => \N__7100\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__7103\,
            I => \DUT.uart_inst0.tx_clk_divider_1_sqmuxa_1_i\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__7100\,
            I => \DUT.uart_inst0.tx_clk_divider_1_sqmuxa_1_i\
        );

    \I__1025\ : InMux
    port map (
            O => \N__7095\,
            I => \N__7092\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__7092\,
            I => \N__7089\
        );

    \I__1023\ : Odrv12
    port map (
            O => \N__7089\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_5\
        );

    \I__1022\ : CascadeMux
    port map (
            O => \N__7086\,
            I => \N__7082\
        );

    \I__1021\ : InMux
    port map (
            O => \N__7085\,
            I => \N__7075\
        );

    \I__1020\ : InMux
    port map (
            O => \N__7082\,
            I => \N__7075\
        );

    \I__1019\ : InMux
    port map (
            O => \N__7081\,
            I => \N__7072\
        );

    \I__1018\ : CascadeMux
    port map (
            O => \N__7080\,
            I => \N__7069\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__7075\,
            I => \N__7064\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__7072\,
            I => \N__7064\
        );

    \I__1015\ : InMux
    port map (
            O => \N__7069\,
            I => \N__7061\
        );

    \I__1014\ : Span4Mux_v
    port map (
            O => \N__7064\,
            I => \N__7058\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__7061\,
            I => \N__7054\
        );

    \I__1012\ : Span4Mux_h
    port map (
            O => \N__7058\,
            I => \N__7051\
        );

    \I__1011\ : InMux
    port map (
            O => \N__7057\,
            I => \N__7048\
        );

    \I__1010\ : Odrv12
    port map (
            O => \N__7054\,
            I => \DUT.uart_inst0.N_47\
        );

    \I__1009\ : Odrv4
    port map (
            O => \N__7051\,
            I => \DUT.uart_inst0.N_47\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__7048\,
            I => \DUT.uart_inst0.N_47\
        );

    \I__1007\ : InMux
    port map (
            O => \N__7041\,
            I => \N__7038\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__7038\,
            I => \DUT.uart_inst0.N_68\
        );

    \I__1005\ : CascadeMux
    port map (
            O => \N__7035\,
            I => \N__7031\
        );

    \I__1004\ : CascadeMux
    port map (
            O => \N__7034\,
            I => \N__7028\
        );

    \I__1003\ : InMux
    port map (
            O => \N__7031\,
            I => \N__7024\
        );

    \I__1002\ : InMux
    port map (
            O => \N__7028\,
            I => \N__7019\
        );

    \I__1001\ : InMux
    port map (
            O => \N__7027\,
            I => \N__7019\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__7024\,
            I => \N__7012\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__7019\,
            I => \N__7009\
        );

    \I__998\ : InMux
    port map (
            O => \N__7018\,
            I => \N__7002\
        );

    \I__997\ : InMux
    port map (
            O => \N__7017\,
            I => \N__7002\
        );

    \I__996\ : InMux
    port map (
            O => \N__7016\,
            I => \N__7002\
        );

    \I__995\ : CascadeMux
    port map (
            O => \N__7015\,
            I => \N__6999\
        );

    \I__994\ : Span4Mux_v
    port map (
            O => \N__7012\,
            I => \N__6992\
        );

    \I__993\ : Span4Mux_v
    port map (
            O => \N__7009\,
            I => \N__6992\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__7002\,
            I => \N__6992\
        );

    \I__991\ : InMux
    port map (
            O => \N__6999\,
            I => \N__6989\
        );

    \I__990\ : Span4Mux_h
    port map (
            O => \N__6992\,
            I => \N__6986\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__6989\,
            I => \DUT.uart_inst0.recv_stateZ0Z_5\
        );

    \I__988\ : Odrv4
    port map (
            O => \N__6986\,
            I => \DUT.uart_inst0.recv_stateZ0Z_5\
        );

    \I__987\ : CascadeMux
    port map (
            O => \N__6981\,
            I => \N__6977\
        );

    \I__986\ : InMux
    port map (
            O => \N__6980\,
            I => \N__6974\
        );

    \I__985\ : InMux
    port map (
            O => \N__6977\,
            I => \N__6971\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__6974\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_2\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__6971\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_2\
        );

    \I__982\ : InMux
    port map (
            O => \N__6966\,
            I => \N__6961\
        );

    \I__981\ : InMux
    port map (
            O => \N__6965\,
            I => \N__6956\
        );

    \I__980\ : InMux
    port map (
            O => \N__6964\,
            I => \N__6956\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__6961\,
            I => \DUT.uart_inst0.rx_countdown_3_2\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__6956\,
            I => \DUT.uart_inst0.rx_countdown_3_2\
        );

    \I__977\ : CascadeMux
    port map (
            O => \N__6951\,
            I => \N__6948\
        );

    \I__976\ : InMux
    port map (
            O => \N__6948\,
            I => \N__6945\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__6945\,
            I => \N__6939\
        );

    \I__974\ : InMux
    port map (
            O => \N__6944\,
            I => \N__6934\
        );

    \I__973\ : InMux
    port map (
            O => \N__6943\,
            I => \N__6934\
        );

    \I__972\ : InMux
    port map (
            O => \N__6942\,
            I => \N__6931\
        );

    \I__971\ : Odrv12
    port map (
            O => \N__6939\,
            I => \DUT.uart_inst0.rx_countdown_3_3\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__6934\,
            I => \DUT.uart_inst0.rx_countdown_3_3\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__6931\,
            I => \DUT.uart_inst0.rx_countdown_3_3\
        );

    \I__968\ : InMux
    port map (
            O => \N__6924\,
            I => \N__6918\
        );

    \I__967\ : InMux
    port map (
            O => \N__6923\,
            I => \N__6913\
        );

    \I__966\ : InMux
    port map (
            O => \N__6922\,
            I => \N__6913\
        );

    \I__965\ : InMux
    port map (
            O => \N__6921\,
            I => \N__6910\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__6918\,
            I => \DUT.uart_inst0.rx_countdown_3_4\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__6913\,
            I => \DUT.uart_inst0.rx_countdown_3_4\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__6910\,
            I => \DUT.uart_inst0.rx_countdown_3_4\
        );

    \I__961\ : CascadeMux
    port map (
            O => \N__6903\,
            I => \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa_0_a2_0_a2_1_cascade_\
        );

    \I__960\ : InMux
    port map (
            O => \N__6900\,
            I => \N__6896\
        );

    \I__959\ : InMux
    port map (
            O => \N__6899\,
            I => \N__6893\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__6896\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_2_2\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__6893\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_2_2\
        );

    \I__956\ : InMux
    port map (
            O => \N__6888\,
            I => \N__6884\
        );

    \I__955\ : InMux
    port map (
            O => \N__6887\,
            I => \N__6881\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__6884\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_12\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__6881\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_12\
        );

    \I__952\ : InMux
    port map (
            O => \N__6876\,
            I => \N__6872\
        );

    \I__951\ : InMux
    port map (
            O => \N__6875\,
            I => \N__6869\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__6872\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_7\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__6869\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_7\
        );

    \I__948\ : CascadeMux
    port map (
            O => \N__6864\,
            I => \N__6861\
        );

    \I__947\ : InMux
    port map (
            O => \N__6861\,
            I => \N__6857\
        );

    \I__946\ : InMux
    port map (
            O => \N__6860\,
            I => \N__6854\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__6857\,
            I => \N__6851\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__6854\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_13\
        );

    \I__943\ : Odrv4
    port map (
            O => \N__6851\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_13\
        );

    \I__942\ : CascadeMux
    port map (
            O => \N__6846\,
            I => \N__6843\
        );

    \I__941\ : InMux
    port map (
            O => \N__6843\,
            I => \N__6839\
        );

    \I__940\ : InMux
    port map (
            O => \N__6842\,
            I => \N__6836\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__6839\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_6\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__6836\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_6\
        );

    \I__937\ : CascadeMux
    port map (
            O => \N__6831\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_8_cascade_\
        );

    \I__936\ : CascadeMux
    port map (
            O => \N__6828\,
            I => \N__6825\
        );

    \I__935\ : InMux
    port map (
            O => \N__6825\,
            I => \N__6821\
        );

    \I__934\ : InMux
    port map (
            O => \N__6824\,
            I => \N__6818\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__6821\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_4\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__6818\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_4\
        );

    \I__931\ : InMux
    port map (
            O => \N__6813\,
            I => \N__6809\
        );

    \I__930\ : InMux
    port map (
            O => \N__6812\,
            I => \N__6806\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__6809\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_3\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__6806\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_3\
        );

    \I__927\ : CascadeMux
    port map (
            O => \N__6801\,
            I => \N__6798\
        );

    \I__926\ : InMux
    port map (
            O => \N__6798\,
            I => \N__6794\
        );

    \I__925\ : InMux
    port map (
            O => \N__6797\,
            I => \N__6791\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__6794\,
            I => \N__6788\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__6791\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_5\
        );

    \I__922\ : Odrv4
    port map (
            O => \N__6788\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_5\
        );

    \I__921\ : CascadeMux
    port map (
            O => \N__6783\,
            I => \N__6780\
        );

    \I__920\ : InMux
    port map (
            O => \N__6780\,
            I => \N__6776\
        );

    \I__919\ : InMux
    port map (
            O => \N__6779\,
            I => \N__6773\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__6776\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_2\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__6773\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_2\
        );

    \I__916\ : CascadeMux
    port map (
            O => \N__6768\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_9_cascade_\
        );

    \I__915\ : CascadeMux
    port map (
            O => \N__6765\,
            I => \N__6760\
        );

    \I__914\ : CascadeMux
    port map (
            O => \N__6764\,
            I => \N__6757\
        );

    \I__913\ : InMux
    port map (
            O => \N__6763\,
            I => \N__6753\
        );

    \I__912\ : InMux
    port map (
            O => \N__6760\,
            I => \N__6748\
        );

    \I__911\ : InMux
    port map (
            O => \N__6757\,
            I => \N__6748\
        );

    \I__910\ : InMux
    port map (
            O => \N__6756\,
            I => \N__6745\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__6753\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__6748\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__6745\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__906\ : CascadeMux
    port map (
            O => \N__6738\,
            I => \N__6735\
        );

    \I__905\ : InMux
    port map (
            O => \N__6735\,
            I => \N__6732\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__6732\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_0_c_RNOZ0\
        );

    \I__903\ : InMux
    port map (
            O => \N__6729\,
            I => \N__6725\
        );

    \I__902\ : InMux
    port map (
            O => \N__6728\,
            I => \N__6722\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__6725\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_1\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__6722\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_1\
        );

    \I__899\ : CascadeMux
    port map (
            O => \N__6717\,
            I => \N__6714\
        );

    \I__898\ : InMux
    port map (
            O => \N__6714\,
            I => \N__6711\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__6711\,
            I => \DUT.uart_inst0.rx_countdown_RNICSMA4Z0Z_1\
        );

    \I__896\ : InMux
    port map (
            O => \N__6708\,
            I => \N__6704\
        );

    \I__895\ : InMux
    port map (
            O => \N__6707\,
            I => \N__6701\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__6704\,
            I => \DUT.uart_inst0.rx_countdown_3_1\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__6701\,
            I => \DUT.uart_inst0.rx_countdown_3_1\
        );

    \I__892\ : InMux
    port map (
            O => \N__6696\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_0\
        );

    \I__891\ : InMux
    port map (
            O => \N__6693\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_1\
        );

    \I__890\ : InMux
    port map (
            O => \N__6690\,
            I => \N__6686\
        );

    \I__889\ : InMux
    port map (
            O => \N__6689\,
            I => \N__6683\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__6686\,
            I => \DUT.uart_inst0.rx_countdownZ1Z_3\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__6683\,
            I => \DUT.uart_inst0.rx_countdownZ1Z_3\
        );

    \I__886\ : CascadeMux
    port map (
            O => \N__6678\,
            I => \N__6675\
        );

    \I__885\ : InMux
    port map (
            O => \N__6675\,
            I => \N__6672\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__6672\,
            I => \N__6669\
        );

    \I__883\ : Odrv4
    port map (
            O => \N__6669\,
            I => \DUT.uart_inst0.rx_countdown_RNIEUMA4Z0Z_3\
        );

    \I__882\ : InMux
    port map (
            O => \N__6666\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_2\
        );

    \I__881\ : InMux
    port map (
            O => \N__6663\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_3\
        );

    \I__880\ : InMux
    port map (
            O => \N__6660\,
            I => \N__6657\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__6657\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_5\
        );

    \I__878\ : InMux
    port map (
            O => \N__6654\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_4\
        );

    \I__877\ : CascadeMux
    port map (
            O => \N__6651\,
            I => \N__6648\
        );

    \I__876\ : InMux
    port map (
            O => \N__6648\,
            I => \N__6645\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__6645\,
            I => \N__6641\
        );

    \I__874\ : InMux
    port map (
            O => \N__6644\,
            I => \N__6638\
        );

    \I__873\ : Odrv4
    port map (
            O => \N__6641\,
            I => \DUT.uart_inst0.rx_countdown_3_5\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__6638\,
            I => \DUT.uart_inst0.rx_countdown_3_5\
        );

    \I__871\ : CascadeMux
    port map (
            O => \N__6633\,
            I => \N__6629\
        );

    \I__870\ : InMux
    port map (
            O => \N__6632\,
            I => \N__6624\
        );

    \I__869\ : InMux
    port map (
            O => \N__6629\,
            I => \N__6624\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__6624\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_4\
        );

    \I__867\ : InMux
    port map (
            O => \N__6621\,
            I => \N__6618\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__6618\,
            I => \DUT.uart_inst0.rx_countdown_RNIFVMA4Z0Z_4\
        );

    \I__865\ : InMux
    port map (
            O => \N__6615\,
            I => \N__6604\
        );

    \I__864\ : InMux
    port map (
            O => \N__6614\,
            I => \N__6604\
        );

    \I__863\ : CascadeMux
    port map (
            O => \N__6613\,
            I => \N__6601\
        );

    \I__862\ : CascadeMux
    port map (
            O => \N__6612\,
            I => \N__6597\
        );

    \I__861\ : CascadeMux
    port map (
            O => \N__6611\,
            I => \N__6592\
        );

    \I__860\ : InMux
    port map (
            O => \N__6610\,
            I => \N__6589\
        );

    \I__859\ : InMux
    port map (
            O => \N__6609\,
            I => \N__6586\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__6604\,
            I => \N__6583\
        );

    \I__857\ : InMux
    port map (
            O => \N__6601\,
            I => \N__6578\
        );

    \I__856\ : InMux
    port map (
            O => \N__6600\,
            I => \N__6578\
        );

    \I__855\ : InMux
    port map (
            O => \N__6597\,
            I => \N__6571\
        );

    \I__854\ : InMux
    port map (
            O => \N__6596\,
            I => \N__6571\
        );

    \I__853\ : InMux
    port map (
            O => \N__6595\,
            I => \N__6571\
        );

    \I__852\ : InMux
    port map (
            O => \N__6592\,
            I => \N__6568\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__6589\,
            I => \N__6565\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__6586\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_15\
        );

    \I__849\ : Odrv4
    port map (
            O => \N__6583\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_15\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__6578\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_15\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__6571\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_15\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__6568\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_15\
        );

    \I__845\ : Odrv4
    port map (
            O => \N__6565\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_15\
        );

    \I__844\ : InMux
    port map (
            O => \N__6552\,
            I => \N__6538\
        );

    \I__843\ : InMux
    port map (
            O => \N__6551\,
            I => \N__6538\
        );

    \I__842\ : InMux
    port map (
            O => \N__6550\,
            I => \N__6538\
        );

    \I__841\ : InMux
    port map (
            O => \N__6549\,
            I => \N__6533\
        );

    \I__840\ : InMux
    port map (
            O => \N__6548\,
            I => \N__6533\
        );

    \I__839\ : InMux
    port map (
            O => \N__6547\,
            I => \N__6528\
        );

    \I__838\ : InMux
    port map (
            O => \N__6546\,
            I => \N__6528\
        );

    \I__837\ : InMux
    port map (
            O => \N__6545\,
            I => \N__6525\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__6538\,
            I => \N__6519\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__6533\,
            I => \N__6512\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__6528\,
            I => \N__6512\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__6525\,
            I => \N__6512\
        );

    \I__832\ : InMux
    port map (
            O => \N__6524\,
            I => \N__6507\
        );

    \I__831\ : InMux
    port map (
            O => \N__6523\,
            I => \N__6507\
        );

    \I__830\ : InMux
    port map (
            O => \N__6522\,
            I => \N__6504\
        );

    \I__829\ : Span4Mux_h
    port map (
            O => \N__6519\,
            I => \N__6497\
        );

    \I__828\ : Span4Mux_v
    port map (
            O => \N__6512\,
            I => \N__6497\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__6507\,
            I => \N__6497\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__6504\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_14\
        );

    \I__825\ : Odrv4
    port map (
            O => \N__6497\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_14\
        );

    \I__824\ : InMux
    port map (
            O => \N__6492\,
            I => \N__6489\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__6489\,
            I => \DUT.uart_inst0.rx_countdown_RNIDTMA4Z0Z_2\
        );

    \I__822\ : IoInMux
    port map (
            O => \N__6486\,
            I => \N__6483\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__6483\,
            I => \wPllLocked_i\
        );

    \I__820\ : InMux
    port map (
            O => \N__6480\,
            I => \N__6477\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__6477\,
            I => \N__6474\
        );

    \I__818\ : Odrv4
    port map (
            O => \N__6474\,
            I => \DUT.uart_inst0.rx_clk_divider_1_5\
        );

    \I__817\ : InMux
    port map (
            O => \N__6471\,
            I => \N__6467\
        );

    \I__816\ : InMux
    port map (
            O => \N__6470\,
            I => \N__6464\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__6467\,
            I => \N__6459\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__6464\,
            I => \N__6459\
        );

    \I__813\ : Odrv12
    port map (
            O => \N__6459\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_5\
        );

    \I__812\ : InMux
    port map (
            O => \N__6456\,
            I => \N__6453\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__6453\,
            I => \N__6450\
        );

    \I__810\ : Odrv4
    port map (
            O => \N__6450\,
            I => \DUT.uart_inst0.rx_clk_divider_1_6\
        );

    \I__809\ : CascadeMux
    port map (
            O => \N__6447\,
            I => \N__6444\
        );

    \I__808\ : InMux
    port map (
            O => \N__6444\,
            I => \N__6440\
        );

    \I__807\ : InMux
    port map (
            O => \N__6443\,
            I => \N__6437\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__6440\,
            I => \N__6432\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__6437\,
            I => \N__6432\
        );

    \I__804\ : Span4Mux_h
    port map (
            O => \N__6432\,
            I => \N__6429\
        );

    \I__803\ : Odrv4
    port map (
            O => \N__6429\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_6\
        );

    \I__802\ : InMux
    port map (
            O => \N__6426\,
            I => \N__6423\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__6423\,
            I => \DUT.fifo_rx_inst.un1_i11_2_i\
        );

    \I__800\ : CascadeMux
    port map (
            O => \N__6420\,
            I => \DUT.fifo_rx_inst.un1_i11_2_i_cascade_\
        );

    \I__799\ : CascadeMux
    port map (
            O => \N__6417\,
            I => \N__6413\
        );

    \I__798\ : InMux
    port map (
            O => \N__6416\,
            I => \N__6408\
        );

    \I__797\ : InMux
    port map (
            O => \N__6413\,
            I => \N__6401\
        );

    \I__796\ : InMux
    port map (
            O => \N__6412\,
            I => \N__6401\
        );

    \I__795\ : InMux
    port map (
            O => \N__6411\,
            I => \N__6401\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__6408\,
            I => \DUT.fifo_rx_inst.N_88\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__6401\,
            I => \DUT.fifo_rx_inst.N_88\
        );

    \I__792\ : InMux
    port map (
            O => \N__6396\,
            I => \N__6386\
        );

    \I__791\ : InMux
    port map (
            O => \N__6395\,
            I => \N__6386\
        );

    \I__790\ : InMux
    port map (
            O => \N__6394\,
            I => \N__6386\
        );

    \I__789\ : CascadeMux
    port map (
            O => \N__6393\,
            I => \N__6381\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__6386\,
            I => \N__6378\
        );

    \I__787\ : InMux
    port map (
            O => \N__6385\,
            I => \N__6371\
        );

    \I__786\ : InMux
    port map (
            O => \N__6384\,
            I => \N__6371\
        );

    \I__785\ : InMux
    port map (
            O => \N__6381\,
            I => \N__6371\
        );

    \I__784\ : Odrv4
    port map (
            O => \N__6378\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_0\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__6371\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_0\
        );

    \I__782\ : InMux
    port map (
            O => \N__6366\,
            I => \N__6360\
        );

    \I__781\ : InMux
    port map (
            O => \N__6365\,
            I => \N__6355\
        );

    \I__780\ : InMux
    port map (
            O => \N__6364\,
            I => \N__6355\
        );

    \I__779\ : CascadeMux
    port map (
            O => \N__6363\,
            I => \N__6352\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__6360\,
            I => \N__6346\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__6355\,
            I => \N__6346\
        );

    \I__776\ : InMux
    port map (
            O => \N__6352\,
            I => \N__6341\
        );

    \I__775\ : InMux
    port map (
            O => \N__6351\,
            I => \N__6341\
        );

    \I__774\ : Odrv4
    port map (
            O => \N__6346\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_1\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__6341\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_1\
        );

    \I__772\ : InMux
    port map (
            O => \N__6336\,
            I => \N__6327\
        );

    \I__771\ : InMux
    port map (
            O => \N__6335\,
            I => \N__6327\
        );

    \I__770\ : InMux
    port map (
            O => \N__6334\,
            I => \N__6320\
        );

    \I__769\ : InMux
    port map (
            O => \N__6333\,
            I => \N__6320\
        );

    \I__768\ : InMux
    port map (
            O => \N__6332\,
            I => \N__6320\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__6327\,
            I => \DUT.fifo_rx_inst.N_85\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__6320\,
            I => \DUT.fifo_rx_inst.N_85\
        );

    \I__765\ : CascadeMux
    port map (
            O => \N__6315\,
            I => \N__6309\
        );

    \I__764\ : CascadeMux
    port map (
            O => \N__6314\,
            I => \N__6306\
        );

    \I__763\ : InMux
    port map (
            O => \N__6313\,
            I => \N__6302\
        );

    \I__762\ : InMux
    port map (
            O => \N__6312\,
            I => \N__6293\
        );

    \I__761\ : InMux
    port map (
            O => \N__6309\,
            I => \N__6293\
        );

    \I__760\ : InMux
    port map (
            O => \N__6306\,
            I => \N__6293\
        );

    \I__759\ : InMux
    port map (
            O => \N__6305\,
            I => \N__6293\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__6302\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_1\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__6293\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_1\
        );

    \I__756\ : CascadeMux
    port map (
            O => \N__6288\,
            I => \DUT.uart_inst0.m5_1_cascade_\
        );

    \I__755\ : CascadeMux
    port map (
            O => \N__6285\,
            I => \N__6282\
        );

    \I__754\ : InMux
    port map (
            O => \N__6282\,
            I => \N__6279\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__6279\,
            I => \N__6276\
        );

    \I__752\ : Odrv4
    port map (
            O => \N__6276\,
            I => \DUT.uart_inst0.N_6_0\
        );

    \I__751\ : CascadeMux
    port map (
            O => \N__6273\,
            I => \DUT.uart_inst0.N_12_cascade_\
        );

    \I__750\ : CascadeMux
    port map (
            O => \N__6270\,
            I => \DUT.uart_inst0.N_7_0_cascade_\
        );

    \I__749\ : CascadeMux
    port map (
            O => \N__6267\,
            I => \N__6262\
        );

    \I__748\ : InMux
    port map (
            O => \N__6266\,
            I => \N__6255\
        );

    \I__747\ : InMux
    port map (
            O => \N__6265\,
            I => \N__6255\
        );

    \I__746\ : InMux
    port map (
            O => \N__6262\,
            I => \N__6255\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__6255\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_3\
        );

    \I__744\ : CascadeMux
    port map (
            O => \N__6252\,
            I => \DUT.uart_inst0.m5_0_1_cascade_\
        );

    \I__743\ : CascadeMux
    port map (
            O => \N__6249\,
            I => \DUT.uart_inst0.N_6_cascade_\
        );

    \I__742\ : InMux
    port map (
            O => \N__6246\,
            I => \N__6234\
        );

    \I__741\ : InMux
    port map (
            O => \N__6245\,
            I => \N__6234\
        );

    \I__740\ : InMux
    port map (
            O => \N__6244\,
            I => \N__6234\
        );

    \I__739\ : InMux
    port map (
            O => \N__6243\,
            I => \N__6234\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__6234\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_2\
        );

    \I__737\ : InMux
    port map (
            O => \N__6231\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_4\
        );

    \I__736\ : InMux
    port map (
            O => \N__6228\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_5\
        );

    \I__735\ : InMux
    port map (
            O => \N__6225\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_6\
        );

    \I__734\ : InMux
    port map (
            O => \N__6222\,
            I => \bfn_12_15_0_\
        );

    \I__733\ : InMux
    port map (
            O => \N__6219\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_8\
        );

    \I__732\ : InMux
    port map (
            O => \N__6216\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_9\
        );

    \I__731\ : InMux
    port map (
            O => \N__6213\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_10\
        );

    \I__730\ : InMux
    port map (
            O => \N__6210\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_11\
        );

    \I__729\ : InMux
    port map (
            O => \N__6207\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_12\
        );

    \I__728\ : CascadeMux
    port map (
            O => \N__6204\,
            I => \DUT.uart_inst0.rx_countdown_RNI8KQG9Z0Z_0_cascade_\
        );

    \I__727\ : CascadeMux
    port map (
            O => \N__6201\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_2_2_cascade_\
        );

    \I__726\ : CascadeMux
    port map (
            O => \N__6198\,
            I => \DUT.uart_inst0.N_42_cascade_\
        );

    \I__725\ : InMux
    port map (
            O => \N__6195\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_0\
        );

    \I__724\ : InMux
    port map (
            O => \N__6192\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_1\
        );

    \I__723\ : InMux
    port map (
            O => \N__6189\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_2\
        );

    \I__722\ : InMux
    port map (
            O => \N__6186\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_3\
        );

    \I__721\ : InMux
    port map (
            O => \N__6183\,
            I => \N__6180\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__6180\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO\
        );

    \I__719\ : CascadeMux
    port map (
            O => \N__6177\,
            I => \N__6172\
        );

    \I__718\ : InMux
    port map (
            O => \N__6176\,
            I => \N__6169\
        );

    \I__717\ : InMux
    port map (
            O => \N__6175\,
            I => \N__6166\
        );

    \I__716\ : InMux
    port map (
            O => \N__6172\,
            I => \N__6163\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__6169\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_13\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__6166\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_13\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__6163\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_13\
        );

    \I__712\ : CascadeMux
    port map (
            O => \N__6156\,
            I => \N__6153\
        );

    \I__711\ : InMux
    port map (
            O => \N__6153\,
            I => \N__6150\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__6150\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO\
        );

    \I__709\ : CascadeMux
    port map (
            O => \N__6147\,
            I => \N__6143\
        );

    \I__708\ : InMux
    port map (
            O => \N__6146\,
            I => \N__6139\
        );

    \I__707\ : InMux
    port map (
            O => \N__6143\,
            I => \N__6136\
        );

    \I__706\ : InMux
    port map (
            O => \N__6142\,
            I => \N__6133\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__6139\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_14\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__6136\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_14\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__6133\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_14\
        );

    \I__702\ : InMux
    port map (
            O => \N__6126\,
            I => \N__6123\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__6123\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO\
        );

    \I__700\ : InMux
    port map (
            O => \N__6120\,
            I => \N__6115\
        );

    \I__699\ : InMux
    port map (
            O => \N__6119\,
            I => \N__6112\
        );

    \I__698\ : InMux
    port map (
            O => \N__6118\,
            I => \N__6109\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__6115\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_15\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__6112\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_15\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__6109\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_15\
        );

    \I__694\ : CascadeMux
    port map (
            O => \N__6102\,
            I => \N__6099\
        );

    \I__693\ : InMux
    port map (
            O => \N__6099\,
            I => \N__6096\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__6096\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO\
        );

    \I__691\ : CascadeMux
    port map (
            O => \N__6093\,
            I => \N__6089\
        );

    \I__690\ : InMux
    port map (
            O => \N__6092\,
            I => \N__6085\
        );

    \I__689\ : InMux
    port map (
            O => \N__6089\,
            I => \N__6082\
        );

    \I__688\ : InMux
    port map (
            O => \N__6088\,
            I => \N__6079\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__6085\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_16\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__6082\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_16\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__6079\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_16\
        );

    \I__684\ : CascadeMux
    port map (
            O => \N__6072\,
            I => \DUT.uart_inst0.N_46_cascade_\
        );

    \I__683\ : InMux
    port map (
            O => \N__6069\,
            I => \N__6066\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__6066\,
            I => \DUT.uart_inst0.rx_countdown_3_0\
        );

    \I__681\ : InMux
    port map (
            O => \N__6063\,
            I => \N__6060\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__6060\,
            I => \DUT.fifo_rx_inst.N_97\
        );

    \I__679\ : CascadeMux
    port map (
            O => \N__6057\,
            I => \N__6054\
        );

    \I__678\ : InMux
    port map (
            O => \N__6054\,
            I => \N__6047\
        );

    \I__677\ : InMux
    port map (
            O => \N__6053\,
            I => \N__6044\
        );

    \I__676\ : InMux
    port map (
            O => \N__6052\,
            I => \N__6037\
        );

    \I__675\ : InMux
    port map (
            O => \N__6051\,
            I => \N__6037\
        );

    \I__674\ : InMux
    port map (
            O => \N__6050\,
            I => \N__6037\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__6047\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_0\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__6044\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_0\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__6037\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_0\
        );

    \I__670\ : InMux
    port map (
            O => \N__6030\,
            I => \N__6020\
        );

    \I__669\ : InMux
    port map (
            O => \N__6029\,
            I => \N__6015\
        );

    \I__668\ : InMux
    port map (
            O => \N__6028\,
            I => \N__6015\
        );

    \I__667\ : InMux
    port map (
            O => \N__6027\,
            I => \N__6012\
        );

    \I__666\ : InMux
    port map (
            O => \N__6026\,
            I => \N__6009\
        );

    \I__665\ : InMux
    port map (
            O => \N__6025\,
            I => \N__6004\
        );

    \I__664\ : InMux
    port map (
            O => \N__6024\,
            I => \N__6004\
        );

    \I__663\ : InMux
    port map (
            O => \N__6023\,
            I => \N__6001\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__6020\,
            I => \N__5996\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__6015\,
            I => \N__5996\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__6012\,
            I => \DUT.wRcvd\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__6009\,
            I => \DUT.wRcvd\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__6004\,
            I => \DUT.wRcvd\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__6001\,
            I => \DUT.wRcvd\
        );

    \I__656\ : Odrv4
    port map (
            O => \N__5996\,
            I => \DUT.wRcvd\
        );

    \I__655\ : CascadeMux
    port map (
            O => \N__5985\,
            I => \N__5982\
        );

    \I__654\ : InMux
    port map (
            O => \N__5982\,
            I => \N__5973\
        );

    \I__653\ : InMux
    port map (
            O => \N__5981\,
            I => \N__5970\
        );

    \I__652\ : InMux
    port map (
            O => \N__5980\,
            I => \N__5965\
        );

    \I__651\ : InMux
    port map (
            O => \N__5979\,
            I => \N__5965\
        );

    \I__650\ : InMux
    port map (
            O => \N__5978\,
            I => \N__5958\
        );

    \I__649\ : InMux
    port map (
            O => \N__5977\,
            I => \N__5958\
        );

    \I__648\ : InMux
    port map (
            O => \N__5976\,
            I => \N__5958\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__5973\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__5970\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__5965\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__5958\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\
        );

    \I__643\ : InMux
    port map (
            O => \N__5949\,
            I => \N__5944\
        );

    \I__642\ : InMux
    port map (
            O => \N__5948\,
            I => \N__5941\
        );

    \I__641\ : InMux
    port map (
            O => \N__5947\,
            I => \N__5938\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__5944\,
            I => \DUT.uart_inst0.rx_clk_dividerZ1Z_1\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__5941\,
            I => \DUT.uart_inst0.rx_clk_dividerZ1Z_1\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__5938\,
            I => \DUT.uart_inst0.rx_clk_dividerZ1Z_1\
        );

    \I__637\ : InMux
    port map (
            O => \N__5931\,
            I => \N__5927\
        );

    \I__636\ : InMux
    port map (
            O => \N__5930\,
            I => \N__5924\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__5927\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_3\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__5924\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_3\
        );

    \I__633\ : CascadeMux
    port map (
            O => \N__5919\,
            I => \N__5916\
        );

    \I__632\ : InMux
    port map (
            O => \N__5916\,
            I => \N__5912\
        );

    \I__631\ : InMux
    port map (
            O => \N__5915\,
            I => \N__5908\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__5912\,
            I => \N__5905\
        );

    \I__629\ : InMux
    port map (
            O => \N__5911\,
            I => \N__5902\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__5908\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_2\
        );

    \I__627\ : Odrv4
    port map (
            O => \N__5905\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_2\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__5902\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_2\
        );

    \I__625\ : CascadeMux
    port map (
            O => \N__5895\,
            I => \N__5891\
        );

    \I__624\ : InMux
    port map (
            O => \N__5894\,
            I => \N__5887\
        );

    \I__623\ : InMux
    port map (
            O => \N__5891\,
            I => \N__5884\
        );

    \I__622\ : InMux
    port map (
            O => \N__5890\,
            I => \N__5881\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__5887\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_1\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__5884\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_1\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__5881\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_1\
        );

    \I__618\ : CascadeMux
    port map (
            O => \N__5874\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_9_cascade_\
        );

    \I__617\ : CascadeMux
    port map (
            O => \N__5871\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_15_cascade_\
        );

    \I__616\ : CascadeMux
    port map (
            O => \N__5868\,
            I => \N__5864\
        );

    \I__615\ : InMux
    port map (
            O => \N__5867\,
            I => \N__5861\
        );

    \I__614\ : InMux
    port map (
            O => \N__5864\,
            I => \N__5858\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__5861\,
            I => \N__5855\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__5858\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_17\
        );

    \I__611\ : Odrv4
    port map (
            O => \N__5855\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_17\
        );

    \I__610\ : InMux
    port map (
            O => \N__5850\,
            I => \N__5847\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__5847\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_12\
        );

    \I__608\ : InMux
    port map (
            O => \N__5844\,
            I => \N__5841\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__5841\,
            I => \DUT.uart_inst0.N_50\
        );

    \I__606\ : CascadeMux
    port map (
            O => \N__5838\,
            I => \DUT.uart_inst0.recv_state_srsts_1_3_cascade_\
        );

    \I__605\ : InMux
    port map (
            O => \N__5835\,
            I => \N__5826\
        );

    \I__604\ : InMux
    port map (
            O => \N__5834\,
            I => \N__5826\
        );

    \I__603\ : InMux
    port map (
            O => \N__5833\,
            I => \N__5826\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__5826\,
            I => \DUT.uart_inst0.recv_stateZ0Z_3\
        );

    \I__601\ : CascadeMux
    port map (
            O => \N__5823\,
            I => \DUT.fifo_rx_inst.N_88_cascade_\
        );

    \I__600\ : CascadeMux
    port map (
            O => \N__5820\,
            I => \N__5817\
        );

    \I__599\ : InMux
    port map (
            O => \N__5817\,
            I => \N__5814\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__5814\,
            I => \DUT.fifo_rx_inst.rFifoCount_RNIK3G92Z0Z_1\
        );

    \I__597\ : CascadeMux
    port map (
            O => \N__5811\,
            I => \N__5806\
        );

    \I__596\ : InMux
    port map (
            O => \N__5810\,
            I => \N__5802\
        );

    \I__595\ : InMux
    port map (
            O => \N__5809\,
            I => \N__5795\
        );

    \I__594\ : InMux
    port map (
            O => \N__5806\,
            I => \N__5795\
        );

    \I__593\ : InMux
    port map (
            O => \N__5805\,
            I => \N__5795\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__5802\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_1\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__5795\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_1\
        );

    \I__590\ : CascadeMux
    port map (
            O => \N__5790\,
            I => \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1Z0Z_0_cascade_\
        );

    \I__589\ : CascadeMux
    port map (
            O => \N__5787\,
            I => \DUT.fifo_rx_inst.N_97_cascade_\
        );

    \I__588\ : CascadeMux
    port map (
            O => \N__5784\,
            I => \N__5781\
        );

    \I__587\ : InMux
    port map (
            O => \N__5781\,
            I => \N__5778\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__5778\,
            I => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0\
        );

    \I__585\ : InMux
    port map (
            O => \N__5775\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_12\
        );

    \I__584\ : InMux
    port map (
            O => \N__5772\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_13\
        );

    \I__583\ : InMux
    port map (
            O => \N__5769\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_14\
        );

    \I__582\ : InMux
    port map (
            O => \N__5766\,
            I => \bfn_11_13_0_\
        );

    \I__581\ : InMux
    port map (
            O => \N__5763\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_16\
        );

    \I__580\ : InMux
    port map (
            O => \N__5760\,
            I => \N__5754\
        );

    \I__579\ : InMux
    port map (
            O => \N__5759\,
            I => \N__5754\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__5754\,
            I => \DUT.uart_inst0.recv_stateZ0Z_4\
        );

    \I__577\ : CascadeMux
    port map (
            O => \N__5751\,
            I => \DUT.uart_inst0.recv_state_ns_0_0_0_cascade_\
        );

    \I__576\ : InMux
    port map (
            O => \N__5748\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_4\
        );

    \I__575\ : InMux
    port map (
            O => \N__5745\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_5\
        );

    \I__574\ : InMux
    port map (
            O => \N__5742\,
            I => \N__5737\
        );

    \I__573\ : InMux
    port map (
            O => \N__5741\,
            I => \N__5734\
        );

    \I__572\ : InMux
    port map (
            O => \N__5740\,
            I => \N__5731\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__5737\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_7\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__5734\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_7\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__5731\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_7\
        );

    \I__568\ : InMux
    port map (
            O => \N__5724\,
            I => \N__5721\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__5721\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO\
        );

    \I__566\ : InMux
    port map (
            O => \N__5718\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_6\
        );

    \I__565\ : CascadeMux
    port map (
            O => \N__5715\,
            I => \N__5711\
        );

    \I__564\ : InMux
    port map (
            O => \N__5714\,
            I => \N__5707\
        );

    \I__563\ : InMux
    port map (
            O => \N__5711\,
            I => \N__5704\
        );

    \I__562\ : InMux
    port map (
            O => \N__5710\,
            I => \N__5701\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__5707\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_8\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__5704\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_8\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__5701\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_8\
        );

    \I__558\ : InMux
    port map (
            O => \N__5694\,
            I => \N__5691\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__5691\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO\
        );

    \I__556\ : InMux
    port map (
            O => \N__5688\,
            I => \bfn_11_12_0_\
        );

    \I__555\ : InMux
    port map (
            O => \N__5685\,
            I => \N__5680\
        );

    \I__554\ : InMux
    port map (
            O => \N__5684\,
            I => \N__5677\
        );

    \I__553\ : InMux
    port map (
            O => \N__5683\,
            I => \N__5674\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__5680\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_9\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__5677\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_9\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__5674\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_9\
        );

    \I__549\ : InMux
    port map (
            O => \N__5667\,
            I => \N__5664\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__5664\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO\
        );

    \I__547\ : InMux
    port map (
            O => \N__5661\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_8\
        );

    \I__546\ : CascadeMux
    port map (
            O => \N__5658\,
            I => \N__5654\
        );

    \I__545\ : InMux
    port map (
            O => \N__5657\,
            I => \N__5650\
        );

    \I__544\ : InMux
    port map (
            O => \N__5654\,
            I => \N__5647\
        );

    \I__543\ : InMux
    port map (
            O => \N__5653\,
            I => \N__5644\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__5650\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_10\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__5647\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_10\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__5644\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_10\
        );

    \I__539\ : InMux
    port map (
            O => \N__5637\,
            I => \N__5634\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__5634\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO\
        );

    \I__537\ : InMux
    port map (
            O => \N__5631\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_9\
        );

    \I__536\ : InMux
    port map (
            O => \N__5628\,
            I => \N__5623\
        );

    \I__535\ : InMux
    port map (
            O => \N__5627\,
            I => \N__5620\
        );

    \I__534\ : InMux
    port map (
            O => \N__5626\,
            I => \N__5617\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__5623\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_11\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__5620\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_11\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__5617\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_11\
        );

    \I__530\ : InMux
    port map (
            O => \N__5610\,
            I => \N__5607\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__5607\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO\
        );

    \I__528\ : InMux
    port map (
            O => \N__5604\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_10\
        );

    \I__527\ : CascadeMux
    port map (
            O => \N__5601\,
            I => \N__5596\
        );

    \I__526\ : CascadeMux
    port map (
            O => \N__5600\,
            I => \N__5593\
        );

    \I__525\ : InMux
    port map (
            O => \N__5599\,
            I => \N__5590\
        );

    \I__524\ : InMux
    port map (
            O => \N__5596\,
            I => \N__5587\
        );

    \I__523\ : InMux
    port map (
            O => \N__5593\,
            I => \N__5584\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__5590\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_12\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__5587\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_12\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__5584\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_12\
        );

    \I__519\ : CascadeMux
    port map (
            O => \N__5577\,
            I => \N__5574\
        );

    \I__518\ : InMux
    port map (
            O => \N__5574\,
            I => \N__5571\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__5571\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO\
        );

    \I__516\ : InMux
    port map (
            O => \N__5568\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_11\
        );

    \I__515\ : CascadeMux
    port map (
            O => \N__5565\,
            I => \DUT.fifo_rx_inst.un1_i11_i_cascade_\
        );

    \I__514\ : InMux
    port map (
            O => \N__5562\,
            I => \N__5559\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__5559\,
            I => \DUT.fifo_rx_inst.un1_i11_i\
        );

    \I__512\ : InMux
    port map (
            O => \N__5556\,
            I => \N__5553\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__5553\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO\
        );

    \I__510\ : InMux
    port map (
            O => \N__5550\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_0\
        );

    \I__509\ : CascadeMux
    port map (
            O => \N__5547\,
            I => \N__5544\
        );

    \I__508\ : InMux
    port map (
            O => \N__5544\,
            I => \N__5541\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__5541\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO\
        );

    \I__506\ : InMux
    port map (
            O => \N__5538\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_1\
        );

    \I__505\ : InMux
    port map (
            O => \N__5535\,
            I => \N__5532\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__5532\,
            I => \DUT.uart_inst0.rx_clk_divider_1_3\
        );

    \I__503\ : InMux
    port map (
            O => \N__5529\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_2\
        );

    \I__502\ : InMux
    port map (
            O => \N__5526\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_3\
        );

    \I__501\ : InMux
    port map (
            O => \N__5523\,
            I => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0\
        );

    \I__500\ : InMux
    port map (
            O => \N__5520\,
            I => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1\
        );

    \I__499\ : CascadeMux
    port map (
            O => \N__5517\,
            I => \DUT.fifo_rx_inst.rFifoData_awe3_cascade_\
        );

    \I__498\ : IoInMux
    port map (
            O => \N__5514\,
            I => \N__5511\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__5511\,
            I => \N__5508\
        );

    \I__496\ : Span12Mux_s3_v
    port map (
            O => \N__5508\,
            I => \N__5505\
        );

    \I__495\ : Odrv12
    port map (
            O => \N__5505\,
            I => \wTxRdData_4\
        );

    \I__494\ : IoInMux
    port map (
            O => \N__5502\,
            I => \N__5499\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__5499\,
            I => \N__5496\
        );

    \I__492\ : Span4Mux_s3_v
    port map (
            O => \N__5496\,
            I => \N__5493\
        );

    \I__491\ : Span4Mux_v
    port map (
            O => \N__5493\,
            I => \N__5490\
        );

    \I__490\ : Span4Mux_h
    port map (
            O => \N__5490\,
            I => \N__5487\
        );

    \I__489\ : Odrv4
    port map (
            O => \N__5487\,
            I => \wTxRdData_1\
        );

    \I__488\ : InMux
    port map (
            O => \N__5484\,
            I => \N__5481\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__5481\,
            I => \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO\
        );

    \I__486\ : CascadeMux
    port map (
            O => \N__5478\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_3_cascade_\
        );

    \I__485\ : InMux
    port map (
            O => \N__5475\,
            I => \N__5472\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__5472\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_11\
        );

    \I__483\ : IoInMux
    port map (
            O => \N__5469\,
            I => \N__5466\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__5466\,
            I => \N__5463\
        );

    \I__481\ : Sp12to4
    port map (
            O => \N__5463\,
            I => \N__5460\
        );

    \I__480\ : Span12Mux_v
    port map (
            O => \N__5460\,
            I => \N__5457\
        );

    \I__479\ : Odrv12
    port map (
            O => \N__5457\,
            I => \wTxRdData_7\
        );

    \I__478\ : IoInMux
    port map (
            O => \N__5454\,
            I => \N__5451\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__5451\,
            I => \N__5448\
        );

    \I__476\ : Span4Mux_s1_v
    port map (
            O => \N__5448\,
            I => \N__5445\
        );

    \I__475\ : Span4Mux_v
    port map (
            O => \N__5445\,
            I => \N__5442\
        );

    \I__474\ : Span4Mux_v
    port map (
            O => \N__5442\,
            I => \N__5439\
        );

    \I__473\ : Span4Mux_h
    port map (
            O => \N__5439\,
            I => \N__5436\
        );

    \I__472\ : Odrv4
    port map (
            O => \N__5436\,
            I => \wTxRdData_0\
        );

    \I__471\ : IoInMux
    port map (
            O => \N__5433\,
            I => \N__5430\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__5430\,
            I => \N__5427\
        );

    \I__469\ : Span12Mux_s9_v
    port map (
            O => \N__5427\,
            I => \N__5424\
        );

    \I__468\ : Span12Mux_v
    port map (
            O => \N__5424\,
            I => \N__5421\
        );

    \I__467\ : Odrv12
    port map (
            O => \N__5421\,
            I => \BTN_N_c\
        );

    \I__466\ : IoInMux
    port map (
            O => \N__5418\,
            I => \N__5415\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__5415\,
            I => \N__5412\
        );

    \I__464\ : Span4Mux_s1_v
    port map (
            O => \N__5412\,
            I => \N__5409\
        );

    \I__463\ : Span4Mux_v
    port map (
            O => \N__5409\,
            I => \N__5406\
        );

    \I__462\ : Span4Mux_v
    port map (
            O => \N__5406\,
            I => \N__5403\
        );

    \I__461\ : Odrv4
    port map (
            O => \N__5403\,
            I => \wTxRdData_3\
        );

    \I__460\ : IoInMux
    port map (
            O => \N__5400\,
            I => \N__5397\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__5397\,
            I => \N__5394\
        );

    \I__458\ : Span12Mux_s8_v
    port map (
            O => \N__5394\,
            I => \N__5391\
        );

    \I__457\ : Odrv12
    port map (
            O => \N__5391\,
            I => \wTxRdData_5\
        );

    \I__456\ : IoInMux
    port map (
            O => \N__5388\,
            I => \N__5385\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__5385\,
            I => \N__5382\
        );

    \I__454\ : Span4Mux_s1_v
    port map (
            O => \N__5382\,
            I => \N__5379\
        );

    \I__453\ : Span4Mux_v
    port map (
            O => \N__5379\,
            I => \N__5376\
        );

    \I__452\ : Span4Mux_v
    port map (
            O => \N__5376\,
            I => \N__5373\
        );

    \I__451\ : Odrv4
    port map (
            O => \N__5373\,
            I => \wTxRdData_2\
        );

    \I__450\ : IoInMux
    port map (
            O => \N__5370\,
            I => \N__5367\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__5367\,
            I => \N__5364\
        );

    \I__448\ : Span12Mux_s10_v
    port map (
            O => \N__5364\,
            I => \N__5361\
        );

    \I__447\ : Odrv12
    port map (
            O => \N__5361\,
            I => \wTxRdData_6\
        );

    \IN_MUX_bfv_17_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_12_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_14_0_\
        );

    \IN_MUX_bfv_12_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_14_0_\
        );

    \IN_MUX_bfv_12_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DUT.uart_inst0.tx_clk_divider_cry_7\,
            carryinitout => \bfn_12_15_0_\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_12_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_11_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DUT.uart_inst0.rx_clk_divider_1_cry_7\,
            carryinitout => \bfn_11_12_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DUT.uart_inst0.rx_clk_divider_1_cry_15\,
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_20_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_17_0_\
        );

    \IN_MUX_bfv_10_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_16_0_\
        );

    \wPllLocked_i_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__6486\,
            GLOBALBUFFEROUTPUT => \wPllLocked_i_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \top_pll_inst.top_pll_inst_RNISDA2\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__12454\,
            GLOBALBUFFEROUTPUT => \wPllLocked_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5484\,
            lcout => \wPllLocked\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIL7JJ_7_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5710\,
            in2 => \_gnd_net_\,
            in3 => \N__5740\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.un2_rx_clk_divider_a_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIHKFQ1_5_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__6443\,
            in1 => \N__6470\,
            in2 => \N__5478\,
            in3 => \N__5475\,
            lcout => \DUT.uart_inst0.un2_rx_clk_divider_a_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIB99J_10_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5683\,
            in1 => \N__5626\,
            in2 => \N__5600\,
            in3 => \N__5653\,
            lcout => \DUT.uart_inst0.un2_rx_clk_divider_a_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_8_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110000100011"
        )
    port map (
            in0 => \N__8319\,
            in1 => \N__5694\,
            in2 => \N__8120\,
            in3 => \N__5714\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13474\,
            ce => \N__12011\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_12_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000000001011"
        )
    port map (
            in0 => \N__8315\,
            in1 => \N__8078\,
            in2 => \N__5577\,
            in3 => \N__5599\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13474\,
            ce => \N__12011\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_7_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101001000101"
        )
    port map (
            in0 => \N__5724\,
            in1 => \N__8316\,
            in2 => \N__8121\,
            in3 => \N__5742\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13474\,
            ce => \N__12011\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_9_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101001000101"
        )
    port map (
            in0 => \N__5667\,
            in1 => \N__8317\,
            in2 => \N__8122\,
            in3 => \N__5685\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13474\,
            ce => \N__12011\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_10_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001001010001"
        )
    port map (
            in0 => \N__5637\,
            in1 => \N__8077\,
            in2 => \N__8341\,
            in3 => \N__5657\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13474\,
            ce => \N__12011\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_11_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110000100011"
        )
    port map (
            in0 => \N__8318\,
            in1 => \N__5610\,
            in2 => \N__8119\,
            in3 => \N__5628\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13474\,
            ce => \N__12011\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_5_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__12296\,
            in1 => \N__5844\,
            in2 => \_gnd_net_\,
            in3 => \N__7365\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13463\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6053\,
            in2 => \N__5784\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_16_0_\,
            carryout => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_1_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5810\,
            in2 => \N__5820\,
            in3 => \N__5523\,
            lcout => \DUT.fifo_rx_inst.rFifoCountZ0Z_1\,
            ltout => OPEN,
            carryin => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0\,
            carryout => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1\,
            clk => \N__13452\,
            ce => 'H',
            sr => \N__13280\
        );

    \DUT.fifo_rx_inst.rFifoCount_2_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001111011100001"
        )
    port map (
            in0 => \N__6027\,
            in1 => \N__6416\,
            in2 => \N__5985\,
            in3 => \N__5520\,
            lcout => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13452\,
            ce => 'H',
            sr => \N__13280\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI96D91_2_1_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6030\,
            in1 => \N__6351\,
            in2 => \N__6393\,
            in3 => \N__5981\,
            lcout => \DUT.fifo_rx_inst.rFifoData_awe3\,
            ltout => \DUT.fifo_rx_inst.rFifoData_awe3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1_1_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__12188\,
            in1 => \_gnd_net_\,
            in2 => \N__5517\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.un1_i11_i\,
            ltout => \DUT.fifo_rx_inst.un1_i11_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_0_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000101"
        )
    port map (
            in0 => \N__6384\,
            in1 => \_gnd_net_\,
            in2 => \N__5565\,
            in3 => \N__6335\,
            lcout => \DUT.fifo_rx_inst.rWritePtrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13448\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_1_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010110100"
        )
    port map (
            in0 => \N__6336\,
            in1 => \N__6385\,
            in2 => \N__6363\,
            in3 => \N__5562\,
            lcout => \DUT.fifo_rx_inst.rWritePtrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13448\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_3_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111111001111"
        )
    port map (
            in0 => \N__6609\,
            in1 => \N__5535\,
            in2 => \N__7080\,
            in3 => \N__6522\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13481\,
            ce => \N__12008\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110000100011"
        )
    port map (
            in0 => \N__8278\,
            in1 => \N__5556\,
            in2 => \N__8140\,
            in3 => \N__5949\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13481\,
            ce => \N__12008\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_2_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000010010100101"
        )
    port map (
            in0 => \N__5915\,
            in1 => \N__8279\,
            in2 => \N__5547\,
            in3 => \N__8114\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13481\,
            ce => \N__12008\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5895\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5948\,
            in2 => \N__8497\,
            in3 => \N__5550\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_0\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8439\,
            in2 => \N__5919\,
            in3 => \N__5538\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_1\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNO_0_3_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5931\,
            in2 => \N__8499\,
            in3 => \N__5529\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_3\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_2\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8440\,
            in2 => \N__8010\,
            in3 => \N__5526\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_3\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNO_0_5_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6471\,
            in2 => \N__8500\,
            in3 => \N__5748\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_5\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_4\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNO_0_6_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8450\,
            in2 => \N__6447\,
            in3 => \N__5745\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_6\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_5\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5741\,
            in2 => \N__8498\,
            in3 => \N__5718\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_6\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8463\,
            in2 => \N__5715\,
            in3 => \N__5688\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_11_12_0_\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5684\,
            in2 => \N__8504\,
            in3 => \N__5661\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_8\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_LUT4_0_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8467\,
            in2 => \N__5658\,
            in3 => \N__5631\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_9\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_LUT4_0_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5627\,
            in2 => \N__8501\,
            in3 => \N__5604\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_10\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_LUT4_0_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8455\,
            in2 => \N__5601\,
            in3 => \N__5568\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_11\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_LUT4_0_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6175\,
            in2 => \N__8502\,
            in3 => \N__5775\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_12\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_LUT4_0_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8459\,
            in2 => \N__6147\,
            in3 => \N__5772\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_13\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_LUT4_0_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6119\,
            in2 => \N__8503\,
            in3 => \N__5769\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_14\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_LUT4_0_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8468\,
            in2 => \N__6093\,
            in3 => \N__5766\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_17_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000000001011"
        )
    port map (
            in0 => \N__8302\,
            in1 => \N__8070\,
            in2 => \N__5868\,
            in3 => \N__5763\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13464\,
            ce => \N__12012\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNI237O_0_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__8329\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8040\,
            lcout => \DUT.uart_inst0.N_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_4_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__12298\,
            in1 => \N__5760\,
            in2 => \N__7015\,
            in3 => \N__7349\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_0_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100010101"
        )
    port map (
            in0 => \N__6026\,
            in1 => \N__8041\,
            in2 => \N__8349\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.recv_state_ns_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_0_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111111011111"
        )
    port map (
            in0 => \N__12297\,
            in1 => \N__5759\,
            in2 => \N__5751\,
            in3 => \N__7348\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13457\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_5_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8334\,
            in1 => \N__5833\,
            in2 => \_gnd_net_\,
            in3 => \N__7406\,
            lcout => \DUT.uart_inst0.N_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_6_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__8333\,
            in1 => \N__5835\,
            in2 => \N__12368\,
            in3 => \N__7358\,
            lcout => \DUT.wRcvd\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13453\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_3_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7308\,
            in2 => \_gnd_net_\,
            in3 => \N__7427\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.recv_state_srsts_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_3_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000001010"
        )
    port map (
            in0 => \N__12320\,
            in1 => \N__5834\,
            in2 => \N__5838\,
            in3 => \N__7359\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13453\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNI9EGD1_0_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110111"
        )
    port map (
            in0 => \N__6051\,
            in1 => \N__13015\,
            in2 => \N__5811\,
            in3 => \N__5977\,
            lcout => \DUT.fifo_rx_inst.N_88\,
            ltout => \DUT.fifo_rx_inst.N_88_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNIK3G92_1_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6025\,
            in2 => \N__5823\,
            in3 => \N__5809\,
            lcout => \DUT.fifo_rx_inst.rFifoCount_RNIK3G92Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5976\,
            in1 => \N__5805\,
            in2 => \_gnd_net_\,
            in3 => \N__6050\,
            lcout => \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1Z0Z_0\,
            ltout => \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNIPTFQ1_0_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6023\,
            in2 => \N__5790\,
            in3 => \N__13016\,
            lcout => \DUT.fifo_rx_inst.N_97\,
            ltout => \DUT.fifo_rx_inst.N_97_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000111"
        )
    port map (
            in0 => \N__5978\,
            in1 => \N__6024\,
            in2 => \N__5787\,
            in3 => \N__6052\,
            lcout => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_0_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110000110100101"
        )
    port map (
            in0 => \N__6063\,
            in1 => \N__6029\,
            in2 => \N__6057\,
            in3 => \N__5980\,
            lcout => \DUT.fifo_rx_inst.rFifoCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13443\,
            ce => 'H',
            sr => \N__13278\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6028\,
            in2 => \_gnd_net_\,
            in3 => \N__5979\,
            lcout => \DUT.fifo_rx_inst.N_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_0_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010111011"
        )
    port map (
            in0 => \N__8280\,
            in1 => \N__8115\,
            in2 => \_gnd_net_\,
            in3 => \N__5894\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13473\,
            ce => \N__12007\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIMQ571_1_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5947\,
            in1 => \N__5930\,
            in2 => \N__8009\,
            in3 => \N__5911\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.un2_rx_clk_divider_a_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIMSP02_16_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6088\,
            in1 => \N__5890\,
            in2 => \N__5874\,
            in3 => \N__5850\,
            lcout => \DUT.uart_inst0.un2_rx_clk_divider_a_15\,
            ltout => \DUT.uart_inst0.un2_rx_clk_divider_a_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_0_c_RNO_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \N__6763\,
            in1 => \_gnd_net_\,
            in2 => \N__5871\,
            in3 => \N__6523\,
            lcout => \DUT.uart_inst0.rx_countdown_3_cry_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNI3ALC_17_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6142\,
            in1 => \N__6118\,
            in2 => \N__6177\,
            in3 => \N__5867\,
            lcout => \DUT.uart_inst0.un2_rx_clk_divider_a_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNICSMA4_1_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__6524\,
            in1 => \N__6729\,
            in2 => \N__6611\,
            in3 => \_gnd_net_\,
            lcout => \DUT.uart_inst0.rx_countdown_RNICSMA4Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_1_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101010000"
        )
    port map (
            in0 => \N__8286\,
            in1 => \N__7018\,
            in2 => \N__8147\,
            in3 => \N__6708\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13462\,
            ce => \N__12009\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_5_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000001010000"
        )
    port map (
            in0 => \N__7016\,
            in1 => \N__8287\,
            in2 => \N__6651\,
            in3 => \N__8137\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13462\,
            ce => \N__12009\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_0_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100000000"
        )
    port map (
            in0 => \N__8285\,
            in1 => \N__7017\,
            in2 => \N__8146\,
            in3 => \N__6069\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13462\,
            ce => \N__12009\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_13_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110000100011"
        )
    port map (
            in0 => \N__8281\,
            in1 => \N__6183\,
            in2 => \N__8144\,
            in3 => \N__6176\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13462\,
            ce => \N__12009\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_14_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000010010100101"
        )
    port map (
            in0 => \N__6146\,
            in1 => \N__8282\,
            in2 => \N__6156\,
            in3 => \N__8138\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13462\,
            ce => \N__12009\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_15_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110000100011"
        )
    port map (
            in0 => \N__8283\,
            in1 => \N__6126\,
            in2 => \N__8145\,
            in3 => \N__6120\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13462\,
            ce => \N__12009\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_16_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000010010100101"
        )
    port map (
            in0 => \N__6092\,
            in1 => \N__8284\,
            in2 => \N__6102\,
            in3 => \N__8139\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13462\,
            ce => \N__12009\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__8301\,
            in1 => \N__7390\,
            in2 => \_gnd_net_\,
            in3 => \N__7306\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_46_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6944\,
            in1 => \N__6923\,
            in2 => \N__6072\,
            in3 => \N__6899\,
            lcout => \DUT.uart_inst0.N_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_0_0_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__6615\,
            in1 => \_gnd_net_\,
            in2 => \N__6765\,
            in3 => \N__6549\,
            lcout => \DUT.uart_inst0.rx_countdown_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNI8KQG9_0_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111011111100"
        )
    port map (
            in0 => \N__6614\,
            in1 => \N__6707\,
            in2 => \N__6764\,
            in3 => \N__6548\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.rx_countdown_RNI8KQG9Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNI8EL7E_0_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__6644\,
            in1 => \_gnd_net_\,
            in2 => \N__6204\,
            in3 => \N__8451\,
            lcout => \DUT.uart_inst0.rx_countdown_8_i_o2_2_2\,
            ltout => \DUT.uart_inst0.rx_countdown_8_i_o2_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_1_c_RNIHH7QT_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6922\,
            in1 => \N__6966\,
            in2 => \N__6201\,
            in3 => \N__6943\,
            lcout => \DUT.uart_inst0.N_42\,
            ltout => \DUT.uart_inst0.N_42_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_1_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000011001100"
        )
    port map (
            in0 => \N__7391\,
            in1 => \N__12366\,
            in2 => \N__6198\,
            in3 => \N__7057\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13456\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7134\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_14_0_\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_1_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7149\,
            in2 => \N__8532\,
            in3 => \N__6195\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_1\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_0\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_1\,
            clk => \N__13451\,
            ce => 'H',
            sr => \N__7107\
        );

    \DUT.uart_inst0.tx_clk_divider_2_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8508\,
            in2 => \N__6783\,
            in3 => \N__6192\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_2\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_1\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_2\,
            clk => \N__13451\,
            ce => 'H',
            sr => \N__7107\
        );

    \DUT.uart_inst0.tx_clk_divider_3_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6813\,
            in2 => \N__8533\,
            in3 => \N__6189\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_3\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_2\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_3\,
            clk => \N__13451\,
            ce => 'H',
            sr => \N__7107\
        );

    \DUT.uart_inst0.tx_clk_divider_4_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8512\,
            in2 => \N__6828\,
            in3 => \N__6186\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_4\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_3\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_4\,
            clk => \N__13451\,
            ce => 'H',
            sr => \N__7107\
        );

    \DUT.uart_inst0.tx_clk_divider_5_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6797\,
            in2 => \N__8534\,
            in3 => \N__6231\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_5\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_4\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_5\,
            clk => \N__13451\,
            ce => 'H',
            sr => \N__7107\
        );

    \DUT.uart_inst0.tx_clk_divider_6_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8516\,
            in2 => \N__6846\,
            in3 => \N__6228\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_6\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_5\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_6\,
            clk => \N__13451\,
            ce => 'H',
            sr => \N__7107\
        );

    \DUT.uart_inst0.tx_clk_divider_7_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6876\,
            in2 => \N__8535\,
            in3 => \N__6225\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_7\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_6\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_7\,
            clk => \N__13451\,
            ce => 'H',
            sr => \N__7107\
        );

    \DUT.uart_inst0.tx_clk_divider_8_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7161\,
            in2 => \N__8538\,
            in3 => \N__6222\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_12_15_0_\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_8\,
            clk => \N__13447\,
            ce => 'H',
            sr => \N__7106\
        );

    \DUT.uart_inst0.tx_clk_divider_9_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8531\,
            in2 => \N__7176\,
            in3 => \N__6219\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_9\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_8\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_9\,
            clk => \N__13447\,
            ce => 'H',
            sr => \N__7106\
        );

    \DUT.uart_inst0.tx_clk_divider_10_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7188\,
            in2 => \N__8536\,
            in3 => \N__6216\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_10\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_9\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_10\,
            clk => \N__13447\,
            ce => 'H',
            sr => \N__7106\
        );

    \DUT.uart_inst0.tx_clk_divider_11_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8524\,
            in2 => \N__7203\,
            in3 => \N__6213\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_11\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_10\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_11\,
            clk => \N__13447\,
            ce => 'H',
            sr => \N__7106\
        );

    \DUT.uart_inst0.tx_clk_divider_12_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6888\,
            in2 => \N__8537\,
            in3 => \N__6210\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_12\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_11\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_12\,
            clk => \N__13447\,
            ce => 'H',
            sr => \N__7106\
        );

    \DUT.uart_inst0.tx_clk_divider_13_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6860\,
            in2 => \_gnd_net_\,
            in3 => \N__6207\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13447\,
            ce => 'H',
            sr => \N__7106\
        );

    \DUT.uart_inst0.tx_clk_divider_0_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__8520\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7133\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13447\,
            ce => 'H',
            sr => \N__7106\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNIUJI11_3_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__6243\,
            in1 => \N__6305\,
            in2 => \N__6267\,
            in3 => \N__7454\,
            lcout => \DUT.uart_inst0.N_62_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_1_3_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__7455\,
            in1 => \N__7286\,
            in2 => \N__6314\,
            in3 => \N__6244\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_0_3_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010100100001"
        )
    port map (
            in0 => \N__6265\,
            in1 => \N__7413\,
            in2 => \N__6273\,
            in3 => \N__7242\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_3_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111100000100"
        )
    port map (
            in0 => \N__7362\,
            in1 => \N__12326\,
            in2 => \N__6270\,
            in3 => \N__6266\,
            lcout => \DUT.uart_inst0.rx_bits_remainingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13442\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_1_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__12324\,
            in1 => \N__7360\,
            in2 => \N__6285\,
            in3 => \N__6312\,
            lcout => \DUT.uart_inst0.rx_bits_remainingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13442\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_1_2_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011111011"
        )
    port map (
            in0 => \N__7456\,
            in1 => \N__7287\,
            in2 => \N__6315\,
            in3 => \N__6245\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.m5_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_0_2_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001111"
        )
    port map (
            in0 => \N__7288\,
            in1 => \N__8336\,
            in2 => \N__6252\,
            in3 => \N__7412\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_2_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101101000000"
        )
    port map (
            in0 => \N__7361\,
            in1 => \N__12325\,
            in2 => \N__6249\,
            in3 => \N__6246\,
            lcout => \DUT.uart_inst0.rx_bits_remainingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13442\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rReadPtr_1_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000101000100"
        )
    port map (
            in0 => \N__6426\,
            in1 => \N__9912\,
            in2 => \N__6417\,
            in3 => \N__9398\,
            lcout => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13439\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__6394\,
            in1 => \N__6364\,
            in2 => \_gnd_net_\,
            in3 => \N__6332\,
            lcout => \DUT.fifo_rx_inst.rFifoData_awe1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rReadPtr_RNI4NC92_0_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100001111"
        )
    port map (
            in0 => \N__6411\,
            in1 => \N__9911\,
            in2 => \N__12192\,
            in3 => \N__9396\,
            lcout => \DUT.fifo_rx_inst.un1_i11_2_i\,
            ltout => \DUT.fifo_rx_inst.un1_i11_2_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rReadPtr_0_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000101"
        )
    port map (
            in0 => \N__9397\,
            in1 => \_gnd_net_\,
            in2 => \N__6420\,
            in3 => \N__6412\,
            lcout => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13439\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6333\,
            in1 => \N__6395\,
            in2 => \_gnd_net_\,
            in3 => \N__6366\,
            lcout => \DUT.fifo_rx_inst.rFifoData_awe0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6396\,
            in1 => \N__6365\,
            in2 => \_gnd_net_\,
            in3 => \N__6334\,
            lcout => \DUT.fifo_rx_inst.rFifoData_awe2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_1_1_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110011001"
        )
    port map (
            in0 => \N__7284\,
            in1 => \N__6313\,
            in2 => \_gnd_net_\,
            in3 => \N__7453\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.m5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_0_1_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100001011"
        )
    port map (
            in0 => \N__8335\,
            in1 => \N__7414\,
            in2 => \N__6288\,
            in3 => \N__7285\,
            lcout => \DUT.uart_inst0.N_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10187\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13436\,
            ce => \N__10013\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9717\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13436\,
            ce => \N__10013\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10118\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13436\,
            ce => \N__10013\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_4_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10222\,
            lcout => \DUT.wRxByte_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13434\,
            ce => \N__7499\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_7_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8350\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.wRxByte_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13434\,
            ce => \N__7499\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_0_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9704\,
            lcout => \DUT.wRxByte_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13433\,
            ce => \N__7500\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.wPllLocked_i_LC_12_30_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12191\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \wPllLocked_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_5_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111110101111"
        )
    port map (
            in0 => \N__6480\,
            in1 => \N__6596\,
            in2 => \N__7086\,
            in3 => \N__6551\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13475\,
            ce => \N__12010\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_6_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011111111"
        )
    port map (
            in0 => \N__6552\,
            in1 => \N__6456\,
            in2 => \N__6612\,
            in3 => \N__7085\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13475\,
            ce => \N__12010\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNIEUMA4_3_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__6690\,
            in1 => \N__6595\,
            in2 => \_gnd_net_\,
            in3 => \N__6550\,
            lcout => \DUT.uart_inst0.rx_countdown_RNIEUMA4Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100011111100"
        )
    port map (
            in0 => \N__8320\,
            in1 => \N__7027\,
            in2 => \N__6951\,
            in3 => \N__8124\,
            lcout => \DUT.uart_inst0.rx_countdownZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13475\,
            ce => \N__12010\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_4_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100000000"
        )
    port map (
            in0 => \N__8123\,
            in1 => \N__8321\,
            in2 => \N__7034\,
            in3 => \N__6924\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13475\,
            ce => \N__12010\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_0_c_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6756\,
            in2 => \N__6738\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_12_0_\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_0_c_RNITO365_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6728\,
            in2 => \N__6717\,
            in3 => \N__6696\,
            lcout => \DUT.uart_inst0.rx_countdown_3_1\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_countdown_3_cry_0\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_1_c_RNI0T465_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6492\,
            in2 => \N__6981\,
            in3 => \N__6693\,
            lcout => \DUT.uart_inst0.rx_countdown_3_2\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_countdown_3_cry_1\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_2_c_RNI31665_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6689\,
            in2 => \N__6678\,
            in3 => \N__6666\,
            lcout => \DUT.uart_inst0.rx_countdown_3_3\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_countdown_3_cry_2\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_3_c_RNI65765_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6621\,
            in2 => \N__6633\,
            in3 => \N__6663\,
            lcout => \DUT.uart_inst0.rx_countdown_3_4\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_countdown_3_cry_3\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_4_c_RNI0QQM4_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001101101100"
        )
    port map (
            in0 => \N__6547\,
            in1 => \N__6660\,
            in2 => \N__6613\,
            in3 => \N__6654\,
            lcout => \DUT.uart_inst0.rx_countdown_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNIFVMA4_4_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__6632\,
            in1 => \N__6600\,
            in2 => \_gnd_net_\,
            in3 => \N__6546\,
            lcout => \DUT.uart_inst0.rx_countdown_RNIFVMA4Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNIDTMA4_2_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \N__6980\,
            in1 => \N__6610\,
            in2 => \_gnd_net_\,
            in3 => \N__6545\,
            lcout => \DUT.uart_inst0.rx_countdown_RNIDTMA4Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_2_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011001100"
        )
    port map (
            in0 => \N__7081\,
            in1 => \N__7041\,
            in2 => \N__7035\,
            in3 => \N__6965\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13465\,
            ce => \N__12013\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_1_c_RNI93IIF_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6964\,
            in1 => \N__6942\,
            in2 => \_gnd_net_\,
            in3 => \N__6921\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa_0_a2_0_a2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNIPAH9U_2_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__7307\,
            in1 => \N__12367\,
            in2 => \N__6903\,
            in3 => \N__6900\,
            lcout => \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_5_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__10536\,
            in1 => \N__8748\,
            in2 => \_gnd_net_\,
            in3 => \N__9302\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13458\,
            ce => \N__12021\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_13_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6887\,
            in1 => \N__6875\,
            in2 => \N__6864\,
            in3 => \N__6842\,
            lcout => \DUT.uart_inst0.un1_tx_clk_divider_8\,
            ltout => \DUT.uart_inst0.un1_tx_clk_divider_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNI7N692_4_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \N__7548\,
            in1 => \N__7719\,
            in2 => \N__6831\,
            in3 => \N__7805\,
            lcout => \DUT.uart_inst0.tx_countdown_RNI7N692Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_RNI2V95_2_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6824\,
            in1 => \N__6812\,
            in2 => \N__6801\,
            in3 => \N__6779\,
            lcout => \DUT.uart_inst0.un1_tx_clk_divider_9\,
            ltout => \DUT.uart_inst0.un1_tx_clk_divider_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNI3J692_0_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__7612\,
            in1 => \N__7755\,
            in2 => \N__6768\,
            in3 => \N__7806\,
            lcout => \DUT.uart_inst0.tx_countdown_3_0\,
            ltout => \DUT.uart_inst0.tx_countdown_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_0_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__9301\,
            in1 => \_gnd_net_\,
            in2 => \N__7206\,
            in3 => \N__10537\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13458\,
            ce => \N__12021\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_RNIR5NO_9_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__7199\,
            in1 => \N__7187\,
            in2 => \_gnd_net_\,
            in3 => \N__7172\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.un1_tx_clk_divider_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_RNIJJMS_0_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__7160\,
            in1 => \N__7148\,
            in2 => \N__7137\,
            in3 => \N__7129\,
            lcout => \DUT.uart_inst0.un1_tx_clk_divider_10\,
            ltout => \DUT.uart_inst0.un1_tx_clk_divider_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNI5L692_2_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__7747\,
            in1 => \N__7584\,
            in2 => \N__7113\,
            in3 => \N__7714\,
            lcout => \DUT.uart_inst0.tx_countdown_RNI5L692Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNI8CH01_0_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__12166\,
            in1 => \N__10538\,
            in2 => \_gnd_net_\,
            in3 => \N__9306\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_clk_divider_1_sqmuxa_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNI5PJS2_0_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__7802\,
            in1 => \N__7761\,
            in2 => \N__7110\,
            in3 => \N__7716\,
            lcout => \DUT.uart_inst0.tx_clk_divider_1_sqmuxa_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_3_cry_0_c_RNO_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7713\,
            in1 => \N__7746\,
            in2 => \N__7617\,
            in3 => \N__7800\,
            lcout => \DUT.uart_inst0.tx_countdown_3_cry_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNI8O692_5_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__7801\,
            in1 => \N__7095\,
            in2 => \N__7759\,
            in3 => \N__7715\,
            lcout => \DUT.uart_inst0.tx_countdown_3_axb_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_0_0_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000100100010"
        )
    port map (
            in0 => \N__7281\,
            in1 => \N__7415\,
            in2 => \N__8352\,
            in3 => \N__7457\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_0_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__12313\,
            in1 => \N__7458\,
            in2 => \N__7461\,
            in3 => \N__7364\,
            lcout => \DUT.uart_inst0.rx_bits_remainingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13449\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_2_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100100010"
        )
    port map (
            in0 => \N__7282\,
            in1 => \N__7428\,
            in2 => \N__8351\,
            in3 => \N__7416\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.recv_state_srsts_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_2_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__12312\,
            in1 => \N__7283\,
            in2 => \N__7368\,
            in3 => \N__7363\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13449\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_2_3_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8348\,
            in2 => \_gnd_net_\,
            in3 => \N__7280\,
            lcout => \DUT.uart_inst0.m5_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_0_RNI0AQO1_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011110111"
        )
    port map (
            in0 => \N__9381\,
            in1 => \N__7226\,
            in2 => \N__9913\,
            in3 => \N__7235\,
            lcout => \DUT.fifo_rx_inst.rTxByte_52_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_0_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__7236\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9988\,
            lcout => \DUT.fifo_rx_inst.rFifoDataro_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13444\,
            ce => 'H',
            sr => \N__13279\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_1_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7958\,
            in2 => \_gnd_net_\,
            in3 => \N__7227\,
            lcout => \DUT.fifo_rx_inst.rFifoDataro_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13444\,
            ce => 'H',
            sr => \N__13279\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__7218\,
            in1 => \N__9908\,
            in2 => \N__7860\,
            in3 => \N__9394\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__9393\,
            in1 => \N__7212\,
            in2 => \N__7974\,
            in3 => \N__9910\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__7506\,
            in1 => \N__9909\,
            in2 => \N__7983\,
            in3 => \N__9395\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10220\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13437\,
            ce => \N__10012\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9606\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13437\,
            ce => \N__10012\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10263\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13437\,
            ce => \N__10012\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9649\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13437\,
            ce => \N__10012\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_2_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9605\,
            lcout => \DUT.wRxByte_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13435\,
            ce => \N__7495\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_3_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10264\,
            lcout => \DUT.wRxByte_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13435\,
            ce => \N__7495\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_1_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9648\,
            lcout => \DUT.wRxByte_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13435\,
            ce => \N__7495\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_5_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10169\,
            lcout => \DUT.wRxByte_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13435\,
            ce => \N__7495\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_6_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10119\,
            lcout => \DUT.wRxByte_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13435\,
            ce => \N__7495\,
            sr => \_gnd_net_\
        );

    \DUT.rTransmit_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__13119\,
            in1 => \N__10499\,
            in2 => \_gnd_net_\,
            in3 => \N__8692\,
            lcout => \DUT.rTransmitZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13482\,
            ce => 'H',
            sr => \N__13286\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNI5UON8_3_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__9182\,
            in1 => \N__8908\,
            in2 => \N__8754\,
            in3 => \N__8793\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_bits_remaining_RNI5UON8Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNIVQ9CI_0_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7527\,
            in3 => \N__7512\,
            lcout => \DUT.uart_inst0.N_109\,
            ltout => \DUT.uart_inst0.N_109_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_1_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__8690\,
            in1 => \N__7634\,
            in2 => \N__7524\,
            in3 => \N__8953\,
            lcout => \DUT.tx_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13476\,
            ce => 'H',
            sr => \N__13285\
        );

    \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIKK41C_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__8831\,
            in1 => \N__8749\,
            in2 => \N__8910\,
            in3 => \N__8870\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIKK41CZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNIN7BAE_0_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8435\,
            in2 => \N__7521\,
            in3 => \N__8794\,
            lcout => \DUT.uart_inst0.N_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_0_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110010"
        )
    port map (
            in0 => \N__10490\,
            in1 => \N__8691\,
            in2 => \N__13078\,
            in3 => \N__7518\,
            lcout => \DUT.tx_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13476\,
            ce => 'H',
            sr => \N__13285\
        );

    \DUT.uart_inst0.tx_state_RNIQSGK9_0_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__8869\,
            in1 => \N__8952\,
            in2 => \N__10509\,
            in3 => \N__8830\,
            lcout => \DUT.uart_inst0.tx_state_ns_i_i_a3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_1_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__10491\,
            in1 => \N__9298\,
            in2 => \_gnd_net_\,
            in3 => \N__8867\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13470\,
            ce => \N__12022\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_4_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__10498\,
            in1 => \N__9297\,
            in2 => \_gnd_net_\,
            in3 => \N__8904\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13470\,
            ce => \N__12022\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_3_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__9296\,
            in1 => \N__8979\,
            in2 => \N__10535\,
            in3 => \N__8829\,
            lcout => \DUT.uart_inst0.tx_countdownZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13470\,
            ce => \N__12022\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_2_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100010101"
        )
    port map (
            in0 => \N__9107\,
            in1 => \N__7635\,
            in2 => \N__10534\,
            in3 => \N__8950\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13470\,
            ce => \N__12022\,
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNISDA2_0_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11889\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12165\,
            lcout => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_3_cry_0_c_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7623\,
            in2 => \N__7616\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_14_0_\,
            carryout => \DUT.uart_inst0.tx_countdown_3_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_3_cry_0_c_RNIPMF33_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7812\,
            in2 => \N__7833\,
            in3 => \N__7593\,
            lcout => \DUT.uart_inst0.tx_countdown_3_1\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_countdown_3_cry_0\,
            carryout => \DUT.uart_inst0.tx_countdown_3_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_3_cry_1_c_RNISQG33_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7590\,
            in2 => \N__7583\,
            in3 => \N__7560\,
            lcout => \DUT.uart_inst0.tx_countdown_3_2\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_countdown_3_cry_1\,
            carryout => \DUT.uart_inst0.tx_countdown_3_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIVUH33_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7689\,
            in2 => \N__7776\,
            in3 => \N__7557\,
            lcout => \DUT.uart_inst0.tx_countdown_3_3\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_countdown_3_cry_2\,
            carryout => \DUT.uart_inst0.tx_countdown_3_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_3_cry_3_c_RNI23J33_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7554\,
            in2 => \N__7547\,
            in3 => \N__7530\,
            lcout => \DUT.uart_inst0.tx_countdown_3_4\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_countdown_3_cry_3\,
            carryout => \DUT.uart_inst0.tx_countdown_3_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_3_cry_4_c_RNIQRFM2_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__7842\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7836\,
            lcout => \DUT.uart_inst0.tx_countdown_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNI4K692_1_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7717\,
            in1 => \N__7751\,
            in2 => \N__7832\,
            in3 => \N__7803\,
            lcout => \DUT.uart_inst0.tx_countdown_RNI4K692Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNI6M692_3_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__7804\,
            in1 => \N__7775\,
            in2 => \N__7760\,
            in3 => \N__7718\,
            lcout => \DUT.uart_inst0.tx_countdown_RNI6M692Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.un1_tx_bits_remaining_cry_0_c_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8700\,
            in2 => \N__9219\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \DUT.uart_inst0.un1_tx_bits_remaining_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_1_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9246\,
            in2 => \N__9240\,
            in3 => \N__7683\,
            lcout => \DUT.uart_inst0.tx_bits_remainingZ0Z_1\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.un1_tx_bits_remaining_cry_0\,
            carryout => \DUT.uart_inst0.un1_tx_bits_remaining_cry_1\,
            clk => \N__13459\,
            ce => 'H',
            sr => \N__8973\
        );

    \DUT.uart_inst0.tx_bits_remaining_2_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9126\,
            in2 => \N__9144\,
            in3 => \N__7680\,
            lcout => \DUT.uart_inst0.tx_bits_remainingZ0Z_2\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.un1_tx_bits_remaining_cry_1\,
            carryout => \DUT.uart_inst0.un1_tx_bits_remaining_cry_2\,
            clk => \N__13459\,
            ce => 'H',
            sr => \N__8973\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9036\,
            in2 => \_gnd_net_\,
            in3 => \N__7677\,
            lcout => \DUT.uart_inst0.tx_bits_remaining_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ft2232h_inst.rRx_n_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100111010101110"
        )
    port map (
            in0 => \N__9555\,
            in1 => \N__7646\,
            in2 => \N__9531\,
            in3 => \N__9460\,
            lcout => \P1A3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13454\,
            ce => 'H',
            sr => \N__13281\
        );

    \rRxRead_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7891\,
            lcout => \rRxReadZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13454\,
            ce => 'H',
            sr => \N__13281\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_0_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11078\,
            in2 => \_gnd_net_\,
            in3 => \N__13173\,
            lcout => \DUT.fifo_tx_inst.rFifoDataro_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13454\,
            ce => 'H',
            sr => \N__13281\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNI250E6_0_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9814\,
            in2 => \_gnd_net_\,
            in3 => \N__7908\,
            lcout => \N_100_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_0_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7892\,
            lcout => \N_100_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100111111"
        )
    port map (
            in0 => \N__9578\,
            in1 => \N__9542\,
            in2 => \N__9945\,
            in3 => \N__9399\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rTxByte_52_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_0_RNIHJV05_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111010101"
        )
    port map (
            in0 => \N__12187\,
            in1 => \N__7902\,
            in2 => \N__7896\,
            in3 => \N__7893\,
            lcout => \rFifoDatarff_0_RNIHJV05\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__9400\,
            in1 => \N__7851\,
            in2 => \N__7872\,
            in3 => \N__9917\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10054\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13445\,
            ce => \N__7965\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9718\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13445\,
            ce => \N__7965\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9658\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13445\,
            ce => \N__7965\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9614\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13445\,
            ce => \N__7965\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10280\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13445\,
            ce => \N__7965\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10229\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13445\,
            ce => \N__7965\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10183\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13445\,
            ce => \N__7965\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10136\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13445\,
            ce => \N__7965\,
            sr => \_gnd_net_\
        );

    \rTxByte_esr_5_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001111"
        )
    port map (
            in0 => \N__10194\,
            in1 => \N__8547\,
            in2 => \N__9964\,
            in3 => \N__7914\,
            lcout => \rTxByteZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13440\,
            ce => \N__9849\,
            sr => \N__9828\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010000110111"
        )
    port map (
            in0 => \N__7947\,
            in1 => \N__9413\,
            in2 => \N__9966\,
            in3 => \N__7938\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rTxByte_esr_4_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__9780\,
            in1 => \N__9958\,
            in2 => \N__7932\,
            in3 => \N__10242\,
            lcout => \rTxByteZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13440\,
            ce => \N__9849\,
            sr => \N__9828\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__7929\,
            in1 => \N__9946\,
            in2 => \N__7923\,
            in3 => \N__9411\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001010111"
        )
    port map (
            in0 => \N__9412\,
            in1 => \N__9954\,
            in2 => \N__8586\,
            in3 => \N__8577\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rTxByte_esr_3_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__8556\,
            in1 => \N__10287\,
            in2 => \N__8571\,
            in3 => \N__9953\,
            lcout => \rTxByteZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13440\,
            ce => \N__9849\,
            sr => \N__9828\
        );

    \rTxByte_esr_6_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001111"
        )
    port map (
            in0 => \N__10143\,
            in1 => \N__8562\,
            in2 => \N__9965\,
            in3 => \N__8568\,
            lcout => \rTxByteZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13440\,
            ce => \N__9849\,
            sr => \N__9828\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10137\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13438\,
            ce => \N__9773\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10170\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13438\,
            ce => \N__9773\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9607\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13438\,
            ce => \N__9773\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10221\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13438\,
            ce => \N__9773\,
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_4_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110000100011"
        )
    port map (
            in0 => \N__8340\,
            in1 => \N__8160\,
            in2 => \N__8148\,
            in3 => \N__8002\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13486\,
            ce => \N__12014\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__8604\,
            in1 => \N__8592\,
            in2 => \N__8627\,
            in3 => \N__9069\,
            lcout => \P1A7_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13486\,
            ce => \N__12014\,
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIFI07_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__11628\,
            in1 => \N__12161\,
            in2 => \_gnd_net_\,
            in3 => \N__10797\,
            lcout => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_3\,
            ltout => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIFI07_2_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__11753\,
            in1 => \_gnd_net_\,
            in2 => \N__8643\,
            in3 => \N__10961\,
            lcout => \fifo_inst.tx_fifo_inst.un18_rRamWrAddr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNIPNAVK_0_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__12424\,
            in1 => \N__9108\,
            in2 => \_gnd_net_\,
            in3 => \N__9068\,
            lcout => \DUT.uart_inst0.N_71_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_RNO_0_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__8689\,
            in1 => \N__8620\,
            in2 => \N__9183\,
            in3 => \N__10316\,
            lcout => \DUT.uart_inst0.N_112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_RNO_3_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__10468\,
            in1 => \N__9178\,
            in2 => \N__10317\,
            in3 => \N__8688\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_out_6_iv_0_a3_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_RNO_2_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__8832\,
            in1 => \N__8954\,
            in2 => \N__8598\,
            in3 => \N__8871\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_out_6_iv_0_a3_1_sx_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_RNO_1_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8798\,
            in1 => \N__8753\,
            in2 => \N__8595\,
            in3 => \N__8909\,
            lcout => \DUT.uart_inst0.N_113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_0_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010011100"
        )
    port map (
            in0 => \N__9106\,
            in1 => \N__9210\,
            in2 => \N__12455\,
            in3 => \N__9067\,
            lcout => \DUT.uart_inst0.tx_bits_remainingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13477\,
            ce => 'H',
            sr => \N__8972\
        );

    \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111111"
        )
    port map (
            in0 => \N__9177\,
            in1 => \N__8866\,
            in2 => \N__8955\,
            in3 => \N__10475\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_countdown_7_i_a3_0_sx_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8799\,
            in1 => \N__8747\,
            in2 => \N__8982\,
            in3 => \N__8903\,
            lcout => \DUT.uart_inst0.N_116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNI8CH01_0_0_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__10503\,
            in1 => \N__12175\,
            in2 => \_gnd_net_\,
            in3 => \N__9300\,
            lcout => \DUT.uart_inst0.N_76_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIMJ5EC_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8951\,
            in1 => \N__8894\,
            in2 => \N__8868\,
            in3 => \N__8820\,
            lcout => \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIMJ5ECZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNI6I8K_1_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8693\,
            in2 => \_gnd_net_\,
            in3 => \N__13052\,
            lcout => \DUT.uart_inst0.N_77\,
            ltout => \DUT.uart_inst0.N_77_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNI9DTT5_0_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__10500\,
            in1 => \N__8789\,
            in2 => \N__8757\,
            in3 => \N__8738\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_state_RNI9DTT5Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNIBV9AJ_0_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011101110"
        )
    port map (
            in0 => \N__9299\,
            in1 => \N__10501\,
            in2 => \N__8712\,
            in3 => \N__8709\,
            lcout => \DUT.uart_inst0.N_99\,
            ltout => \DUT.uart_inst0.N_99_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.un1_tx_bits_remaining_cry_0_c_RNO_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \N__9211\,
            in1 => \N__12381\,
            in2 => \N__8703\,
            in3 => \N__9099\,
            lcout => \DUT.uart_inst0.un1_tx_bits_remaining_cry_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNIIAMI1_1_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001111"
        )
    port map (
            in0 => \N__9173\,
            in1 => \N__8694\,
            in2 => \N__13065\,
            in3 => \N__10502\,
            lcout => \DUT.uart_inst0.N_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_3_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__9295\,
            in1 => \N__10539\,
            in2 => \N__12417\,
            in3 => \N__9252\,
            lcout => \DUT.uart_inst0.tx_bits_remainingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13466\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNIAIE4L_1_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \N__9239\,
            in1 => \N__9100\,
            in2 => \N__12418\,
            in3 => \N__9058\,
            lcout => \DUT.uart_inst0.tx_bits_remaining_RNIAIE4LZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_3_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9139\,
            in1 => \N__9235\,
            in2 => \N__9120\,
            in3 => \N__9212\,
            lcout => \DUT.uart_inst0.N_124\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ft2232h_inst.rFifoState_RNIRPB71_0_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__9461\,
            in1 => \N__9502\,
            in2 => \_gnd_net_\,
            in3 => \N__9524\,
            lcout => \fifo_inst.ft2232h_inst.rFifoStatec_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNIBJE4L_2_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \N__9140\,
            in1 => \N__9101\,
            in2 => \N__12419\,
            in3 => \N__9059\,
            lcout => \DUT.uart_inst0.tx_bits_remaining_RNIBJE4LZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ft2232h_inst.rFifoState_RNO_0_0_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9462\,
            in1 => \N__9503\,
            in2 => \_gnd_net_\,
            in3 => \N__9525\,
            lcout => \fifo_inst.ft2232h_inst.N_103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNO_1_3_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010011010"
        )
    port map (
            in0 => \N__9119\,
            in1 => \N__9102\,
            in2 => \N__12420\,
            in3 => \N__9060\,
            lcout => \DUT.uart_inst0.un1_tx_bits_remaining_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ft2232h_inst.rFifoState_1_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__9453\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9527\,
            lcout => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13460\,
            ce => 'H',
            sr => \N__13282\
        );

    \fifo_inst.ft2232h_inst.rTx_n_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100000011101010"
        )
    port map (
            in0 => \N__8998\,
            in1 => \N__13920\,
            in2 => \N__13872\,
            in3 => \N__12959\,
            lcout => \P1A4_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13460\,
            ce => 'H',
            sr => \N__13282\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_3_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9774\,
            in2 => \_gnd_net_\,
            in3 => \N__9579\,
            lcout => \DUT.fifo_rx_inst.rFifoDataro_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13460\,
            ce => 'H',
            sr => \N__13282\
        );

    \fifo_inst.ft2232h_inst.rFifoState_2_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9567\,
            lcout => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13460\,
            ce => 'H',
            sr => \N__13282\
        );

    \fifo_inst.ft2232h_inst.rFifoState_0_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__9561\,
            in1 => \N__13919\,
            in2 => \N__13871\,
            in3 => \N__9554\,
            lcout => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13460\,
            ce => 'H',
            sr => \N__13282\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_2_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10082\,
            in2 => \_gnd_net_\,
            in3 => \N__9543\,
            lcout => \DUT.fifo_rx_inst.rFifoDataro_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13460\,
            ce => 'H',
            sr => \N__13282\
        );

    \fifo_inst.ft2232h_inst.rFifoState_3_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__9526\,
            in1 => \N__9504\,
            in2 => \_gnd_net_\,
            in3 => \N__9454\,
            lcout => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13460\,
            ce => 'H',
            sr => \N__13282\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__10023\,
            in1 => \N__9959\,
            in2 => \N__9423\,
            in3 => \N__9414\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rTxByte_esr_0_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__9960\,
            in1 => \N__9792\,
            in2 => \N__9348\,
            in3 => \N__9735\,
            lcout => \rTxByteZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13455\,
            ce => \N__9845\,
            sr => \N__9827\
        );

    \rTxByte_esr_7_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__10092\,
            in1 => \N__9963\,
            in2 => \N__9345\,
            in3 => \N__9330\,
            lcout => \rTxByteZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13455\,
            ce => \N__9845\,
            sr => \N__9827\
        );

    \rTxByte_esr_1_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010111011"
        )
    port map (
            in0 => \N__9798\,
            in1 => \N__9961\,
            in2 => \N__9678\,
            in3 => \N__9318\,
            lcout => \rTxByteZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13455\,
            ce => \N__9845\,
            sr => \N__9827\
        );

    \rTxByte_esr_2_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000011"
        )
    port map (
            in0 => \N__9627\,
            in1 => \N__9962\,
            in2 => \N__9858\,
            in3 => \N__9786\,
            lcout => \rTxByteZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13455\,
            ce => \N__9845\,
            sr => \N__9827\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9726\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13450\,
            ce => \N__9772\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10058\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13450\,
            ce => \N__9772\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9666\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13450\,
            ce => \N__9772\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10281\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13450\,
            ce => \N__9772\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10059\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13446\,
            ce => \N__10083\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9725\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13446\,
            ce => \N__10083\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9665\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13446\,
            ce => \N__10083\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9618\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13446\,
            ce => \N__10083\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10273\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13446\,
            ce => \N__10083\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10233\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13446\,
            ce => \N__10083\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10188\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13446\,
            ce => \N__10083\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10129\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13446\,
            ce => \N__10083\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10044\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13441\,
            ce => \N__10014\,
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIGLV01_2_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__9972\,
            in1 => \N__11577\,
            in2 => \N__12476\,
            in3 => \N__10742\,
            lcout => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_2_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10743\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12160\,
            lcout => \fifo_inst.tx_fifo_inst.rRamRdAddr_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13491\,
            ce => \N__11288\,
            sr => \N__13289\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_1_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12159\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10359\,
            lcout => \fifo_inst.tx_fifo_inst.rRamRdAddr_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13491\,
            ce => \N__11288\,
            sr => \N__13289\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIFI07_0_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__10790\,
            in1 => \N__12164\,
            in2 => \_gnd_net_\,
            in3 => \N__11627\,
            lcout => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_0_1_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__10346\,
            in1 => \N__11575\,
            in2 => \N__12456\,
            in3 => \N__10358\,
            lcout => \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_1_1\,
            ltout => \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_RNI_1_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__11476\,
            in1 => \_gnd_net_\,
            in2 => \N__10362\,
            in3 => \_gnd_net_\,
            lcout => \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIZ0Z_1\,
            ltout => \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_1_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__10347\,
            in1 => \N__12428\,
            in2 => \N__10338\,
            in3 => \N__11576\,
            lcout => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_1\,
            ltout => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_2_1_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11660\,
            in1 => \N__10762\,
            in2 => \N__10320\,
            in3 => \N__10724\,
            lcout => \fifo_inst.tx_fifo_inst.un15_rRamRdAddr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_0_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000001010"
        )
    port map (
            in0 => \N__11016\,
            in1 => \N__10305\,
            in2 => \N__11061\,
            in3 => \N__10533\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13487\,
            ce => \N__10376\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_3_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010101100"
        )
    port map (
            in0 => \N__10569\,
            in1 => \N__10926\,
            in2 => \N__10547\,
            in3 => \N__11060\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13487\,
            ce => \N__10376\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_1_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__11055\,
            in1 => \N__10526\,
            in2 => \N__11094\,
            in3 => \N__10293\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13487\,
            ce => \N__10376\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_2_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010101100"
        )
    port map (
            in0 => \N__10299\,
            in1 => \N__12648\,
            in2 => \N__10546\,
            in3 => \N__11059\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13487\,
            ce => \N__10376\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_7_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__11052\,
            in1 => \N__10908\,
            in2 => \_gnd_net_\,
            in3 => \N__10545\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13483\,
            ce => \N__10383\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_4_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__10389\,
            in1 => \N__11053\,
            in2 => \N__10623\,
            in3 => \N__10543\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13483\,
            ce => \N__10383\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_6_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010000000100"
        )
    port map (
            in0 => \N__11051\,
            in1 => \N__10599\,
            in2 => \N__10548\,
            in3 => \N__10560\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13483\,
            ce => \N__10383\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_5_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000110000"
        )
    port map (
            in0 => \N__10554\,
            in1 => \N__11054\,
            in2 => \N__11112\,
            in3 => \N__10544\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13483\,
            ce => \N__10383\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12876\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13478\,
            ce => \N__11157\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13231\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13478\,
            ce => \N__11157\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12918\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13478\,
            ce => \N__11157\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14012\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13478\,
            ce => \N__11157\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12522\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13478\,
            ce => \N__11157\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111110011"
        )
    port map (
            in0 => \N__10659\,
            in1 => \N__10608\,
            in2 => \N__12759\,
            in3 => \N__12849\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__11202\,
            in1 => \N__10590\,
            in2 => \N__10626\,
            in3 => \N__12757\,
            lcout => \DUT.rFifoDatarx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11242\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13471\,
            ce => \N__13181\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14004\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13471\,
            ce => \N__13181\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111110011"
        )
    port map (
            in0 => \N__10578\,
            in1 => \N__12543\,
            in2 => \N__12758\,
            in3 => \N__12848\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__11190\,
            in1 => \N__10584\,
            in2 => \N__10602\,
            in3 => \N__12756\,
            lcout => \DUT.rFifoDatarx_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12613\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13467\,
            ce => \N__11156\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11243\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13467\,
            ce => \N__11156\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12583\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13467\,
            ce => \N__11156\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12582\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13461\,
            ce => \N__13954\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11247\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13461\,
            ce => \N__13954\,
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIDL6N_7_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__10650\,
            in1 => \N__13854\,
            in2 => \N__12480\,
            in3 => \N__10673\,
            lcout => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_7_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__10674\,
            in1 => \_gnd_net_\,
            in2 => \N__12477\,
            in3 => \_gnd_net_\,
            lcout => \fifo_inst.tx_fifo_inst.rRamRdAddr_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13497\,
            ce => \N__11287\,
            sr => \N__13292\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_4_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10701\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12462\,
            lcout => \fifo_inst.tx_fifo_inst.rRamRdAddr_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13497\,
            ce => \N__11287\,
            sr => \N__13292\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIKR111_4_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__11580\,
            in1 => \N__10644\,
            in2 => \N__12478\,
            in3 => \N__10700\,
            lcout => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_6_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10686\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12463\,
            lcout => \fifo_inst.tx_fifo_inst.rRamRdAddr_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13497\,
            ce => \N__11287\,
            sr => \N__13292\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIO1411_6_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__11579\,
            in1 => \N__10638\,
            in2 => \N__12479\,
            in3 => \N__10685\,
            lcout => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_0_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__12461\,
            in1 => \N__11494\,
            in2 => \_gnd_net_\,
            in3 => \N__11543\,
            lcout => \fifo_inst.tx_fifo_inst.rRamRdAddr_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13497\,
            ce => \N__11287\,
            sr => \N__13292\
        );

    \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1_c_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10632\,
            in2 => \N__11495\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1_c_RNI5G02_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10766\,
            in3 => \N__10734\,
            lcout => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1_c_RNI5GZ0Z02\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1\,
            carryout => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI6I12_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11516\,
            in3 => \N__10731\,
            lcout => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI6IZ0Z12\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2\,
            carryout => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_3_c_RNI7K22_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10720\,
            in2 => \_gnd_net_\,
            in3 => \N__10692\,
            lcout => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_3_c_RNI7KZ0Z22\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_3\,
            carryout => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_4_c_RNI44E4_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__12162\,
            in1 => \_gnd_net_\,
            in2 => \N__11659\,
            in3 => \N__10689\,
            lcout => \fifo_inst.tx_fifo_inst.rRamRdAddr_rst_4\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_4\,
            carryout => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_5_c_RNI9O42_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10852\,
            in3 => \N__10677\,
            lcout => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_5_c_RNI9OZ0Z42\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_5\,
            carryout => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_6_c_RNIAQ52_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10882\,
            in3 => \N__10665\,
            lcout => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_6_c_RNIAQZ0Z52\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_6\,
            carryout => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_7_c_RNI7AH4_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__11443\,
            in1 => \N__12163\,
            in2 => \_gnd_net_\,
            in3 => \N__10662\,
            lcout => \fifo_inst.tx_fifo_inst.rRamRdAddr_rst_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ft2232h_inst.rTxRdEn_RNIS0VN_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10896\,
            in2 => \_gnd_net_\,
            in3 => \N__13828\,
            lcout => \fifo_inst.rTxRdEn_RNIS0VN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNISDA2_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__12171\,
            in1 => \N__11620\,
            in2 => \_gnd_net_\,
            in3 => \N__11744\,
            lcout => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ft2232h_inst.rFifoState_RNIG8PK_4_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__13827\,
            in1 => \N__12169\,
            in2 => \_gnd_net_\,
            in3 => \N__13911\,
            lcout => \fifo_inst.ft2232h_inst.rFifoState_RNIG8PKZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_3_1_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__10889\,
            in1 => \N__10853\,
            in2 => \N__11421\,
            in3 => \N__10827\,
            lcout => \fifo_inst.tx_fifo_inst.un15_rRamRdAddr\,
            ltout => \fifo_inst.tx_fifo_inst.un15_rRamRdAddr_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_RNISDA2_0_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12453\,
            in2 => \N__10821\,
            in3 => \N__11486\,
            lcout => OPEN,
            ltout => \fifo_inst.tx_fifo_inst.rRamRdAddr_rst_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_RNISJ0L_0_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10818\,
            in2 => \N__10809\,
            in3 => \N__13826\,
            lcout => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ft2232h_inst.rTxRdEn_fast_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__13829\,
            in1 => \N__12170\,
            in2 => \_gnd_net_\,
            in3 => \N__13912\,
            lcout => \fifo_inst.rTxRdEn_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13492\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11745\,
            in2 => \N__11775\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_12_0_\,
            carryout => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNII2L4_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11604\,
            in2 => \_gnd_net_\,
            in3 => \N__10806\,
            lcout => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNII2LZ0Z4\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1\,
            carryout => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIJ4M4_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10803\,
            in2 => \_gnd_net_\,
            in3 => \N__10779\,
            lcout => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIJ4MZ0Z4\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2\,
            carryout => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIK6N4_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10920\,
            in2 => \_gnd_net_\,
            in3 => \N__10776\,
            lcout => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIK6NZ0Z4\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3\,
            carryout => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_4_c_RNIHM27_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__12179\,
            in1 => \_gnd_net_\,
            in2 => \N__11822\,
            in3 => \N__10989\,
            lcout => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_5\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_4\,
            carryout => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNIIO37_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11928\,
            in2 => \_gnd_net_\,
            in3 => \N__10986\,
            lcout => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNIIOZ0Z37\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5\,
            carryout => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNIJQ47_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10983\,
            in2 => \_gnd_net_\,
            in3 => \N__10971\,
            lcout => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNIJQZ0Z47\,
            ltout => OPEN,
            carryin => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6\,
            carryout => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_7_c_RNIKS57_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__10948\,
            in1 => \N__12180\,
            in2 => \_gnd_net_\,
            in3 => \N__10968\,
            lcout => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__13194\,
            in1 => \N__12724\,
            in2 => \N__11904\,
            in3 => \N__12845\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__12725\,
            in1 => \N__11256\,
            in2 => \N__10935\,
            in3 => \N__10932\,
            lcout => \DUT.rFifoDatarx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIGK17_0_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12186\,
            in2 => \_gnd_net_\,
            in3 => \N__11852\,
            lcout => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__10914\,
            in1 => \N__12726\,
            in2 => \N__11184\,
            in3 => \N__11691\,
            lcout => \DUT.rFifoDatarx_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__12837\,
            in1 => \N__13971\,
            in2 => \N__12748\,
            in3 => \N__10902\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__12723\,
            in1 => \N__10998\,
            in2 => \N__11121\,
            in3 => \N__11118\,
            lcout => \DUT.rFifoDatarx_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111110011"
        )
    port map (
            in0 => \N__11910\,
            in1 => \N__12855\,
            in2 => \N__12747\,
            in3 => \N__12836\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__11103\,
            in1 => \N__11196\,
            in2 => \N__11097\,
            in3 => \N__12722\,
            lcout => \DUT.rFifoDatarx_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000111111"
        )
    port map (
            in0 => \N__13518\,
            in1 => \N__11136\,
            in2 => \N__12746\,
            in3 => \N__12835\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoDataror_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_0_RNIJBAM_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110101"
        )
    port map (
            in0 => \N__11172\,
            in1 => \N__11082\,
            in2 => \N__11064\,
            in3 => \N__12721\,
            lcout => \DUT.rFifoDataror_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__12720\,
            in1 => \N__11025\,
            in2 => \N__11007\,
            in3 => \N__12939\,
            lcout => \DUT.rFifoDatarxZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12928\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13479\,
            ce => \N__13538\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14005\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13479\,
            ce => \N__13538\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12635\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13479\,
            ce => \N__13538\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13238\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13479\,
            ce => \N__13538\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11241\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13479\,
            ce => \N__13538\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12886\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13479\,
            ce => \N__13538\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12588\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13479\,
            ce => \N__13538\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12530\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13479\,
            ce => \N__13538\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_1_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11171\,
            in2 => \_gnd_net_\,
            in3 => \N__13945\,
            lcout => \DUT.fifo_tx_inst.rFifoDataro_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13472\,
            ce => 'H',
            sr => \N__13284\
        );

    \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_1_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__11337\,
            in1 => \N__11363\,
            in2 => \_gnd_net_\,
            in3 => \N__13139\,
            lcout => \DUT.fifo_tx_inst.N_105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__13140\,
            in1 => \N__11364\,
            in2 => \_gnd_net_\,
            in3 => \N__11338\,
            lcout => \DUT.fifo_tx_inst.rFifoData_awe2\,
            ltout => \DUT.fifo_tx_inst.rFifoData_awe2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_2_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11139\,
            in3 => \N__11135\,
            lcout => \DUT.fifo_tx_inst.rFifoDataro_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13472\,
            ce => 'H',
            sr => \N__13284\
        );

    \DUT.fifo_tx_inst.rWritePtr_1_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100000100"
        )
    port map (
            in0 => \N__13138\,
            in1 => \N__11336\,
            in2 => \N__11376\,
            in3 => \N__11362\,
            lcout => \DUT.fifo_tx_inst.rWritePtrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13468\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_RNIN79A_2_1_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__11360\,
            in1 => \N__13022\,
            in2 => \N__11339\,
            in3 => \N__13573\,
            lcout => \DUT.fifo_tx_inst.rFifoData_awe3\,
            ltout => \DUT.fifo_tx_inst.rFifoData_awe3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_RNIJLJC_1_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__12190\,
            in1 => \_gnd_net_\,
            in2 => \N__11379\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_tx_inst.un1_i11_i\,
            ltout => \DUT.fifo_tx_inst.un1_i11_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_0_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000101"
        )
    port map (
            in0 => \N__11335\,
            in1 => \_gnd_net_\,
            in2 => \N__11367\,
            in3 => \N__13137\,
            lcout => \DUT.fifo_tx_inst.rWritePtrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13468\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_RNIN79A_0_1_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__11361\,
            in1 => \_gnd_net_\,
            in2 => \N__11340\,
            in3 => \N__13136\,
            lcout => \DUT.fifo_tx_inst.rFifoData_awe1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIFO7N_8_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11298\,
            in1 => \N__13843\,
            in2 => \_gnd_net_\,
            in3 => \N__11309\,
            lcout => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_5_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11684\,
            lcout => \fifo_inst.tx_fifo_inst.rRamRdAddr_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13498\,
            ce => \N__11292\,
            sr => \N__13293\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_8_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11310\,
            lcout => \fifo_inst.tx_fifo_inst.rRamRdAddr_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13498\,
            ce => \N__11292\,
            sr => \N__13293\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_3_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__12460\,
            in1 => \_gnd_net_\,
            in2 => \N__11544\,
            in3 => \N__11597\,
            lcout => \fifo_inst.tx_fifo_inst.rRamRdAddr_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13498\,
            ce => \N__11292\,
            sr => \N__13293\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_RNI9F4N_5_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__11685\,
            in1 => \_gnd_net_\,
            in2 => \N__13838\,
            in3 => \N__11673\,
            lcout => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNI111S_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__11864\,
            in1 => \N__11781\,
            in2 => \N__11402\,
            in3 => \N__11637\,
            lcout => \fifo_inst.tx_fifo_inst.un18_rRamWrAddr\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIEGV6_0_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12177\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11411\,
            lcout => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI20C4_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12436\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11598\,
            lcout => OPEN,
            ltout => \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI20CZ0Z4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIIO011_3_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__11586\,
            in1 => \N__11578\,
            in2 => \N__11547\,
            in3 => \N__11536\,
            lcout => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_3\,
            ltout => \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.rRamRdAddr_RNI_8_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__11487\,
            in1 => \_gnd_net_\,
            in2 => \N__11448\,
            in3 => \N__11444\,
            lcout => \fifo_inst.tx_fifo_inst.un15_rRamRdAddr_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ft2232h_inst.rTxRdEn_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010100000101000"
        )
    port map (
            in0 => \N__12176\,
            in1 => \N__13913\,
            in2 => \N__13839\,
            in3 => \_gnd_net_\,
            lcout => \fifo_inst.wTxRdEn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13495\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIEGV6_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11412\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12178\,
            lcout => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNISDA2_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12184\,
            in2 => \_gnd_net_\,
            in3 => \N__11939\,
            lcout => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNISDA2_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12185\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11882\,
            lcout => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIGK17_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11853\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12183\,
            lcout => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_4\,
            ltout => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIQIBG_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11818\,
            in1 => \N__11795\,
            in2 => \N__11784\,
            in3 => \N__11702\,
            lcout => \fifo_inst.tx_fifo_inst.un18_rRamWrAddr_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNISDA2_2_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11718\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12182\,
            lcout => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_1\,
            ltout => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNI_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11763\,
            in3 => \N__11749\,
            lcout => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIZ0\,
            ltout => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNISDA2_1_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11712\,
            in3 => \N__12181\,
            lcout => \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__12834\,
            in1 => \N__11895\,
            in2 => \N__12745\,
            in3 => \N__12492\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rReadPtr_RNINFEP_0_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__12846\,
            in1 => \N__13114\,
            in2 => \_gnd_net_\,
            in3 => \N__13082\,
            lcout => \DUT.fifo_tx_inst.N_101\,
            ltout => \DUT.fifo_tx_inst.N_101_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rReadPtr_RNILV421_1_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011111111"
        )
    port map (
            in0 => \N__12713\,
            in1 => \_gnd_net_\,
            in2 => \N__12483\,
            in3 => \N__12435\,
            lcout => \DUT.fifo_tx_inst.un1_i11_2_i\,
            ltout => \DUT.fifo_tx_inst.un1_i11_2_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rReadPtr_0_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000001010"
        )
    port map (
            in0 => \N__12847\,
            in1 => \N__13115\,
            in2 => \N__12195\,
            in3 => \N__13083\,
            lcout => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13489\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNISDA2_0_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12189\,
            in2 => \_gnd_net_\,
            in3 => \N__11940\,
            lcout => \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rReadPtr_1_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__12730\,
            in1 => \N__11922\,
            in2 => \_gnd_net_\,
            in3 => \N__11916\,
            lcout => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13489\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12933\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13488\,
            ce => \N__13961\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12891\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13488\,
            ce => \N__13961\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13239\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13488\,
            ce => \N__13961\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12531\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13488\,
            ce => \N__13961\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12636\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13488\,
            ce => \N__13961\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__12838\,
            in1 => \N__12945\,
            in2 => \N__12749\,
            in3 => \N__12897\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12929\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13484\,
            ce => \N__13185\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12887\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13484\,
            ce => \N__13185\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001101100111"
        )
    port map (
            in0 => \N__12734\,
            in1 => \N__12839\,
            in2 => \N__12597\,
            in3 => \N__12786\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__12780\,
            in1 => \N__12774\,
            in2 => \N__12762\,
            in3 => \N__12735\,
            lcout => \DUT.rFifoDatarx_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12631\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13480\,
            ce => \N__13174\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12584\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13480\,
            ce => \N__13174\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12529\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13480\,
            ce => \N__13174\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13221\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13480\,
            ce => \N__13174\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNIN9O8_0_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__13567\,
            in1 => \N__13610\,
            in2 => \_gnd_net_\,
            in3 => \N__13656\,
            lcout => \DUT.N_93\,
            ltout => \DUT.N_93_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNIEBIJ_0_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13017\,
            in2 => \N__13146\,
            in3 => \N__13079\,
            lcout => \DUT.fifo_tx_inst.N_98\,
            ltout => \DUT.fifo_tx_inst.N_98_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000111"
        )
    port map (
            in0 => \N__13569\,
            in1 => \N__13019\,
            in2 => \N__13143\,
            in3 => \N__13657\,
            lcout => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNIMBD3_2_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__13568\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13018\,
            lcout => \DUT.fifo_tx_inst.N_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNO_0_2_LC_18_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001011110000"
        )
    port map (
            in0 => \N__13081\,
            in1 => \N__13021\,
            in2 => \N__13577\,
            in3 => \N__13110\,
            lcout => \DUT.fifo_tx_inst.un1_rFifoCount_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNIBPFM_1_LC_18_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__13020\,
            in1 => \N__13109\,
            in2 => \N__13614\,
            in3 => \N__13080\,
            lcout => \DUT.fifo_tx_inst.rFifoCount_RNIBPFMZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_0_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010000111"
        )
    port map (
            in0 => \N__13026\,
            in1 => \N__13578\,
            in2 => \N__13667\,
            in3 => \N__12972\,
            lcout => \DUT.fifo_tx_inst.rFifoCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13469\,
            ce => 'H',
            sr => \N__13283\
        );

    \fifo_inst.ft2232h_inst.rFifoState_4_LC_20_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__12966\,
            in1 => \N__13898\,
            in2 => \_gnd_net_\,
            in3 => \N__13863\,
            lcout => \fifo_inst.ft2232h_inst.rFifoStateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13496\,
            ce => 'H',
            sr => \N__13291\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_20_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14016\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13493\,
            ce => \N__13962\,
            sr => \_gnd_net_\
        );

    \fifo_inst.ft2232h_inst.rTxBusReady_LC_20_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110101010"
        )
    port map (
            in0 => \N__13929\,
            in1 => \N__13907\,
            in2 => \N__13870\,
            in3 => \N__13686\,
            lcout => \rTxBusReady\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13490\,
            ce => 'H',
            sr => \N__13288\
        );

    \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13668\,
            in2 => \N__13638\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_20_17_0_\,
            carryout => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_1_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13609\,
            in2 => \N__13626\,
            in3 => \N__13593\,
            lcout => \DUT.fifo_tx_inst.rFifoCountZ0Z_1\,
            ltout => OPEN,
            carryin => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0\,
            carryout => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1\,
            clk => \N__13485\,
            ce => 'H',
            sr => \N__13287\
        );

    \DUT.fifo_tx_inst.rFifoCount_2_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13590\,
            in2 => \_gnd_net_\,
            in3 => \N__13581\,
            lcout => \DUT.fifo_tx_inst.rFifoCountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13485\,
            ce => 'H',
            sr => \N__13287\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_3_LC_21_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13539\,
            in2 => \_gnd_net_\,
            in3 => \N__13514\,
            lcout => \DUT.fifo_tx_inst.rFifoDataro_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__13494\,
            ce => 'H',
            sr => \N__13290\
        );
end \INTERFACE\;
