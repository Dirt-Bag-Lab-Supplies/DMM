// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Mar 30 2020 12:32:26

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    ioFifoData,
    P1A9,
    P1A1,
    P1A8,
    oRx_n,
    P1A7,
    P1A3,
    iTxE_n,
    iRxF_n,
    iClk,
    P1A2,
    BTN_N,
    BTN1,
    oTx_n,
    P1A4);

    output [7:0] ioFifoData;
    output P1A9;
    input P1A1;
    output P1A8;
    output oRx_n;
    output P1A7;
    output P1A3;
    input iTxE_n;
    input iRxF_n;
    input iClk;
    output P1A2;
    input BTN_N;
    input BTN1;
    output oTx_n;
    output P1A4;

    wire N__14220;
    wire N__14206;
    wire N__14205;
    wire N__14204;
    wire N__14197;
    wire N__14196;
    wire N__14195;
    wire N__14188;
    wire N__14187;
    wire N__14186;
    wire N__14179;
    wire N__14178;
    wire N__14177;
    wire N__14170;
    wire N__14169;
    wire N__14168;
    wire N__14161;
    wire N__14160;
    wire N__14159;
    wire N__14152;
    wire N__14151;
    wire N__14150;
    wire N__14143;
    wire N__14142;
    wire N__14141;
    wire N__14134;
    wire N__14133;
    wire N__14132;
    wire N__14125;
    wire N__14124;
    wire N__14123;
    wire N__14116;
    wire N__14115;
    wire N__14114;
    wire N__14107;
    wire N__14106;
    wire N__14105;
    wire N__14098;
    wire N__14097;
    wire N__14096;
    wire N__14089;
    wire N__14088;
    wire N__14087;
    wire N__14080;
    wire N__14079;
    wire N__14078;
    wire N__14071;
    wire N__14070;
    wire N__14069;
    wire N__14062;
    wire N__14061;
    wire N__14060;
    wire N__14053;
    wire N__14052;
    wire N__14051;
    wire N__14044;
    wire N__14043;
    wire N__14042;
    wire N__14035;
    wire N__14034;
    wire N__14033;
    wire N__14016;
    wire N__14013;
    wire N__14012;
    wire N__14009;
    wire N__14006;
    wire N__14005;
    wire N__14004;
    wire N__14001;
    wire N__13998;
    wire N__13995;
    wire N__13992;
    wire N__13987;
    wire N__13982;
    wire N__13979;
    wire N__13976;
    wire N__13971;
    wire N__13968;
    wire N__13965;
    wire N__13962;
    wire N__13961;
    wire N__13958;
    wire N__13955;
    wire N__13954;
    wire N__13949;
    wire N__13946;
    wire N__13945;
    wire N__13942;
    wire N__13939;
    wire N__13936;
    wire N__13929;
    wire N__13926;
    wire N__13923;
    wire N__13920;
    wire N__13919;
    wire N__13914;
    wire N__13913;
    wire N__13912;
    wire N__13911;
    wire N__13908;
    wire N__13907;
    wire N__13904;
    wire N__13899;
    wire N__13898;
    wire N__13895;
    wire N__13892;
    wire N__13887;
    wire N__13884;
    wire N__13877;
    wire N__13872;
    wire N__13871;
    wire N__13870;
    wire N__13867;
    wire N__13864;
    wire N__13863;
    wire N__13860;
    wire N__13855;
    wire N__13854;
    wire N__13853;
    wire N__13850;
    wire N__13847;
    wire N__13844;
    wire N__13843;
    wire N__13840;
    wire N__13839;
    wire N__13838;
    wire N__13835;
    wire N__13830;
    wire N__13829;
    wire N__13828;
    wire N__13827;
    wire N__13826;
    wire N__13823;
    wire N__13820;
    wire N__13817;
    wire N__13814;
    wire N__13811;
    wire N__13808;
    wire N__13805;
    wire N__13796;
    wire N__13791;
    wire N__13788;
    wire N__13783;
    wire N__13770;
    wire N__13769;
    wire N__13766;
    wire N__13765;
    wire N__13764;
    wire N__13763;
    wire N__13762;
    wire N__13759;
    wire N__13756;
    wire N__13753;
    wire N__13750;
    wire N__13749;
    wire N__13746;
    wire N__13743;
    wire N__13740;
    wire N__13733;
    wire N__13730;
    wire N__13729;
    wire N__13724;
    wire N__13719;
    wire N__13716;
    wire N__13713;
    wire N__13710;
    wire N__13705;
    wire N__13702;
    wire N__13699;
    wire N__13696;
    wire N__13693;
    wire N__13690;
    wire N__13687;
    wire N__13686;
    wire N__13683;
    wire N__13678;
    wire N__13675;
    wire N__13668;
    wire N__13667;
    wire N__13664;
    wire N__13661;
    wire N__13658;
    wire N__13657;
    wire N__13656;
    wire N__13653;
    wire N__13650;
    wire N__13645;
    wire N__13638;
    wire N__13635;
    wire N__13632;
    wire N__13629;
    wire N__13626;
    wire N__13623;
    wire N__13620;
    wire N__13617;
    wire N__13614;
    wire N__13611;
    wire N__13610;
    wire N__13609;
    wire N__13604;
    wire N__13601;
    wire N__13598;
    wire N__13593;
    wire N__13590;
    wire N__13587;
    wire N__13584;
    wire N__13581;
    wire N__13578;
    wire N__13577;
    wire N__13574;
    wire N__13573;
    wire N__13570;
    wire N__13569;
    wire N__13568;
    wire N__13567;
    wire N__13564;
    wire N__13561;
    wire N__13552;
    wire N__13549;
    wire N__13544;
    wire N__13539;
    wire N__13538;
    wire N__13535;
    wire N__13532;
    wire N__13529;
    wire N__13526;
    wire N__13523;
    wire N__13518;
    wire N__13515;
    wire N__13514;
    wire N__13511;
    wire N__13508;
    wire N__13505;
    wire N__13500;
    wire N__13499;
    wire N__13498;
    wire N__13497;
    wire N__13496;
    wire N__13495;
    wire N__13494;
    wire N__13493;
    wire N__13492;
    wire N__13491;
    wire N__13490;
    wire N__13489;
    wire N__13488;
    wire N__13487;
    wire N__13486;
    wire N__13485;
    wire N__13484;
    wire N__13483;
    wire N__13482;
    wire N__13481;
    wire N__13480;
    wire N__13479;
    wire N__13478;
    wire N__13477;
    wire N__13476;
    wire N__13475;
    wire N__13474;
    wire N__13473;
    wire N__13472;
    wire N__13471;
    wire N__13470;
    wire N__13469;
    wire N__13468;
    wire N__13467;
    wire N__13466;
    wire N__13465;
    wire N__13464;
    wire N__13463;
    wire N__13462;
    wire N__13461;
    wire N__13460;
    wire N__13459;
    wire N__13458;
    wire N__13457;
    wire N__13456;
    wire N__13455;
    wire N__13454;
    wire N__13453;
    wire N__13452;
    wire N__13451;
    wire N__13450;
    wire N__13449;
    wire N__13448;
    wire N__13447;
    wire N__13446;
    wire N__13445;
    wire N__13444;
    wire N__13443;
    wire N__13442;
    wire N__13441;
    wire N__13440;
    wire N__13439;
    wire N__13438;
    wire N__13437;
    wire N__13436;
    wire N__13435;
    wire N__13434;
    wire N__13433;
    wire N__13296;
    wire N__13293;
    wire N__13292;
    wire N__13291;
    wire N__13290;
    wire N__13289;
    wire N__13288;
    wire N__13287;
    wire N__13286;
    wire N__13285;
    wire N__13284;
    wire N__13283;
    wire N__13282;
    wire N__13281;
    wire N__13280;
    wire N__13279;
    wire N__13278;
    wire N__13245;
    wire N__13242;
    wire N__13239;
    wire N__13238;
    wire N__13235;
    wire N__13232;
    wire N__13231;
    wire N__13228;
    wire N__13225;
    wire N__13222;
    wire N__13221;
    wire N__13214;
    wire N__13211;
    wire N__13208;
    wire N__13205;
    wire N__13202;
    wire N__13199;
    wire N__13194;
    wire N__13191;
    wire N__13188;
    wire N__13185;
    wire N__13182;
    wire N__13181;
    wire N__13178;
    wire N__13175;
    wire N__13174;
    wire N__13173;
    wire N__13168;
    wire N__13165;
    wire N__13162;
    wire N__13159;
    wire N__13156;
    wire N__13153;
    wire N__13146;
    wire N__13143;
    wire N__13140;
    wire N__13139;
    wire N__13138;
    wire N__13137;
    wire N__13136;
    wire N__13131;
    wire N__13124;
    wire N__13119;
    wire N__13116;
    wire N__13115;
    wire N__13114;
    wire N__13111;
    wire N__13110;
    wire N__13109;
    wire N__13104;
    wire N__13101;
    wire N__13098;
    wire N__13095;
    wire N__13092;
    wire N__13083;
    wire N__13082;
    wire N__13081;
    wire N__13080;
    wire N__13079;
    wire N__13078;
    wire N__13073;
    wire N__13066;
    wire N__13065;
    wire N__13062;
    wire N__13059;
    wire N__13056;
    wire N__13053;
    wire N__13052;
    wire N__13049;
    wire N__13044;
    wire N__13041;
    wire N__13038;
    wire N__13029;
    wire N__13026;
    wire N__13023;
    wire N__13022;
    wire N__13021;
    wire N__13020;
    wire N__13019;
    wire N__13018;
    wire N__13017;
    wire N__13016;
    wire N__13015;
    wire N__13012;
    wire N__13009;
    wire N__13000;
    wire N__12997;
    wire N__12992;
    wire N__12983;
    wire N__12980;
    wire N__12977;
    wire N__12972;
    wire N__12969;
    wire N__12966;
    wire N__12963;
    wire N__12960;
    wire N__12959;
    wire N__12956;
    wire N__12953;
    wire N__12950;
    wire N__12945;
    wire N__12942;
    wire N__12939;
    wire N__12936;
    wire N__12933;
    wire N__12930;
    wire N__12929;
    wire N__12928;
    wire N__12925;
    wire N__12922;
    wire N__12919;
    wire N__12918;
    wire N__12911;
    wire N__12908;
    wire N__12905;
    wire N__12902;
    wire N__12897;
    wire N__12894;
    wire N__12891;
    wire N__12888;
    wire N__12887;
    wire N__12886;
    wire N__12883;
    wire N__12880;
    wire N__12877;
    wire N__12876;
    wire N__12869;
    wire N__12866;
    wire N__12863;
    wire N__12860;
    wire N__12855;
    wire N__12852;
    wire N__12849;
    wire N__12848;
    wire N__12847;
    wire N__12846;
    wire N__12845;
    wire N__12840;
    wire N__12839;
    wire N__12838;
    wire N__12837;
    wire N__12836;
    wire N__12835;
    wire N__12834;
    wire N__12829;
    wire N__12826;
    wire N__12823;
    wire N__12820;
    wire N__12817;
    wire N__12810;
    wire N__12807;
    wire N__12800;
    wire N__12795;
    wire N__12786;
    wire N__12783;
    wire N__12780;
    wire N__12777;
    wire N__12774;
    wire N__12771;
    wire N__12768;
    wire N__12765;
    wire N__12762;
    wire N__12759;
    wire N__12758;
    wire N__12757;
    wire N__12756;
    wire N__12753;
    wire N__12750;
    wire N__12749;
    wire N__12748;
    wire N__12747;
    wire N__12746;
    wire N__12745;
    wire N__12736;
    wire N__12735;
    wire N__12734;
    wire N__12731;
    wire N__12730;
    wire N__12727;
    wire N__12726;
    wire N__12725;
    wire N__12724;
    wire N__12723;
    wire N__12722;
    wire N__12721;
    wire N__12720;
    wire N__12717;
    wire N__12714;
    wire N__12713;
    wire N__12710;
    wire N__12707;
    wire N__12700;
    wire N__12697;
    wire N__12694;
    wire N__12687;
    wire N__12674;
    wire N__12669;
    wire N__12666;
    wire N__12663;
    wire N__12648;
    wire N__12645;
    wire N__12642;
    wire N__12639;
    wire N__12636;
    wire N__12635;
    wire N__12632;
    wire N__12631;
    wire N__12628;
    wire N__12625;
    wire N__12622;
    wire N__12619;
    wire N__12614;
    wire N__12613;
    wire N__12610;
    wire N__12607;
    wire N__12604;
    wire N__12597;
    wire N__12594;
    wire N__12591;
    wire N__12588;
    wire N__12585;
    wire N__12584;
    wire N__12583;
    wire N__12582;
    wire N__12579;
    wire N__12576;
    wire N__12573;
    wire N__12570;
    wire N__12567;
    wire N__12562;
    wire N__12559;
    wire N__12556;
    wire N__12553;
    wire N__12550;
    wire N__12543;
    wire N__12540;
    wire N__12537;
    wire N__12534;
    wire N__12531;
    wire N__12530;
    wire N__12529;
    wire N__12526;
    wire N__12523;
    wire N__12522;
    wire N__12519;
    wire N__12514;
    wire N__12511;
    wire N__12508;
    wire N__12505;
    wire N__12502;
    wire N__12499;
    wire N__12492;
    wire N__12489;
    wire N__12486;
    wire N__12483;
    wire N__12480;
    wire N__12479;
    wire N__12478;
    wire N__12477;
    wire N__12476;
    wire N__12473;
    wire N__12470;
    wire N__12467;
    wire N__12464;
    wire N__12463;
    wire N__12462;
    wire N__12461;
    wire N__12460;
    wire N__12457;
    wire N__12456;
    wire N__12455;
    wire N__12454;
    wire N__12453;
    wire N__12450;
    wire N__12437;
    wire N__12436;
    wire N__12435;
    wire N__12432;
    wire N__12429;
    wire N__12428;
    wire N__12425;
    wire N__12424;
    wire N__12421;
    wire N__12420;
    wire N__12419;
    wire N__12418;
    wire N__12417;
    wire N__12414;
    wire N__12411;
    wire N__12408;
    wire N__12405;
    wire N__12402;
    wire N__12399;
    wire N__12394;
    wire N__12391;
    wire N__12388;
    wire N__12385;
    wire N__12382;
    wire N__12381;
    wire N__12378;
    wire N__12375;
    wire N__12372;
    wire N__12369;
    wire N__12368;
    wire N__12367;
    wire N__12366;
    wire N__12363;
    wire N__12360;
    wire N__12351;
    wire N__12340;
    wire N__12337;
    wire N__12330;
    wire N__12327;
    wire N__12326;
    wire N__12325;
    wire N__12324;
    wire N__12321;
    wire N__12320;
    wire N__12317;
    wire N__12314;
    wire N__12313;
    wire N__12312;
    wire N__12309;
    wire N__12304;
    wire N__12299;
    wire N__12298;
    wire N__12297;
    wire N__12296;
    wire N__12293;
    wire N__12290;
    wire N__12283;
    wire N__12278;
    wire N__12273;
    wire N__12268;
    wire N__12265;
    wire N__12262;
    wire N__12259;
    wire N__12254;
    wire N__12251;
    wire N__12246;
    wire N__12241;
    wire N__12236;
    wire N__12233;
    wire N__12224;
    wire N__12219;
    wire N__12216;
    wire N__12211;
    wire N__12208;
    wire N__12203;
    wire N__12200;
    wire N__12195;
    wire N__12192;
    wire N__12191;
    wire N__12190;
    wire N__12189;
    wire N__12188;
    wire N__12187;
    wire N__12186;
    wire N__12185;
    wire N__12184;
    wire N__12183;
    wire N__12182;
    wire N__12181;
    wire N__12180;
    wire N__12179;
    wire N__12178;
    wire N__12177;
    wire N__12176;
    wire N__12175;
    wire N__12172;
    wire N__12171;
    wire N__12170;
    wire N__12169;
    wire N__12168;
    wire N__12167;
    wire N__12166;
    wire N__12165;
    wire N__12164;
    wire N__12163;
    wire N__12162;
    wire N__12161;
    wire N__12160;
    wire N__12159;
    wire N__12156;
    wire N__12153;
    wire N__12150;
    wire N__12147;
    wire N__12144;
    wire N__12141;
    wire N__12130;
    wire N__12125;
    wire N__12118;
    wire N__12115;
    wire N__12112;
    wire N__12105;
    wire N__12102;
    wire N__12099;
    wire N__12096;
    wire N__12093;
    wire N__12090;
    wire N__12085;
    wire N__12082;
    wire N__12077;
    wire N__12074;
    wire N__12071;
    wire N__12068;
    wire N__12065;
    wire N__12062;
    wire N__12059;
    wire N__12056;
    wire N__12053;
    wire N__12050;
    wire N__12047;
    wire N__12044;
    wire N__12041;
    wire N__12038;
    wire N__12035;
    wire N__12032;
    wire N__12029;
    wire N__12026;
    wire N__12023;
    wire N__12022;
    wire N__12021;
    wire N__12018;
    wire N__12015;
    wire N__12014;
    wire N__12013;
    wire N__12012;
    wire N__12011;
    wire N__12010;
    wire N__12009;
    wire N__12008;
    wire N__12007;
    wire N__11946;
    wire N__11943;
    wire N__11940;
    wire N__11939;
    wire N__11936;
    wire N__11933;
    wire N__11928;
    wire N__11925;
    wire N__11922;
    wire N__11919;
    wire N__11916;
    wire N__11913;
    wire N__11910;
    wire N__11907;
    wire N__11904;
    wire N__11901;
    wire N__11898;
    wire N__11895;
    wire N__11892;
    wire N__11889;
    wire N__11886;
    wire N__11883;
    wire N__11882;
    wire N__11879;
    wire N__11876;
    wire N__11871;
    wire N__11868;
    wire N__11865;
    wire N__11864;
    wire N__11861;
    wire N__11858;
    wire N__11853;
    wire N__11852;
    wire N__11849;
    wire N__11846;
    wire N__11841;
    wire N__11838;
    wire N__11835;
    wire N__11832;
    wire N__11829;
    wire N__11826;
    wire N__11823;
    wire N__11822;
    wire N__11819;
    wire N__11818;
    wire N__11815;
    wire N__11812;
    wire N__11809;
    wire N__11806;
    wire N__11799;
    wire N__11796;
    wire N__11795;
    wire N__11792;
    wire N__11789;
    wire N__11784;
    wire N__11781;
    wire N__11778;
    wire N__11775;
    wire N__11772;
    wire N__11769;
    wire N__11766;
    wire N__11763;
    wire N__11760;
    wire N__11757;
    wire N__11754;
    wire N__11753;
    wire N__11750;
    wire N__11749;
    wire N__11746;
    wire N__11745;
    wire N__11744;
    wire N__11741;
    wire N__11738;
    wire N__11735;
    wire N__11732;
    wire N__11729;
    wire N__11718;
    wire N__11715;
    wire N__11712;
    wire N__11709;
    wire N__11706;
    wire N__11703;
    wire N__11702;
    wire N__11699;
    wire N__11696;
    wire N__11691;
    wire N__11688;
    wire N__11685;
    wire N__11684;
    wire N__11681;
    wire N__11678;
    wire N__11673;
    wire N__11670;
    wire N__11667;
    wire N__11664;
    wire N__11661;
    wire N__11660;
    wire N__11659;
    wire N__11656;
    wire N__11653;
    wire N__11650;
    wire N__11645;
    wire N__11642;
    wire N__11637;
    wire N__11634;
    wire N__11631;
    wire N__11628;
    wire N__11627;
    wire N__11624;
    wire N__11621;
    wire N__11620;
    wire N__11617;
    wire N__11614;
    wire N__11611;
    wire N__11604;
    wire N__11601;
    wire N__11598;
    wire N__11597;
    wire N__11594;
    wire N__11591;
    wire N__11586;
    wire N__11583;
    wire N__11580;
    wire N__11579;
    wire N__11578;
    wire N__11577;
    wire N__11576;
    wire N__11575;
    wire N__11570;
    wire N__11567;
    wire N__11564;
    wire N__11559;
    wire N__11556;
    wire N__11547;
    wire N__11544;
    wire N__11543;
    wire N__11540;
    wire N__11537;
    wire N__11536;
    wire N__11533;
    wire N__11530;
    wire N__11527;
    wire N__11520;
    wire N__11517;
    wire N__11516;
    wire N__11513;
    wire N__11510;
    wire N__11507;
    wire N__11504;
    wire N__11499;
    wire N__11496;
    wire N__11495;
    wire N__11494;
    wire N__11491;
    wire N__11488;
    wire N__11487;
    wire N__11486;
    wire N__11483;
    wire N__11480;
    wire N__11477;
    wire N__11476;
    wire N__11473;
    wire N__11470;
    wire N__11467;
    wire N__11462;
    wire N__11459;
    wire N__11448;
    wire N__11445;
    wire N__11444;
    wire N__11443;
    wire N__11440;
    wire N__11437;
    wire N__11434;
    wire N__11431;
    wire N__11428;
    wire N__11421;
    wire N__11418;
    wire N__11415;
    wire N__11412;
    wire N__11411;
    wire N__11406;
    wire N__11403;
    wire N__11402;
    wire N__11399;
    wire N__11396;
    wire N__11393;
    wire N__11390;
    wire N__11387;
    wire N__11384;
    wire N__11379;
    wire N__11376;
    wire N__11373;
    wire N__11370;
    wire N__11367;
    wire N__11364;
    wire N__11363;
    wire N__11362;
    wire N__11361;
    wire N__11360;
    wire N__11357;
    wire N__11354;
    wire N__11347;
    wire N__11340;
    wire N__11339;
    wire N__11338;
    wire N__11337;
    wire N__11336;
    wire N__11335;
    wire N__11332;
    wire N__11329;
    wire N__11324;
    wire N__11315;
    wire N__11310;
    wire N__11309;
    wire N__11306;
    wire N__11303;
    wire N__11298;
    wire N__11295;
    wire N__11292;
    wire N__11289;
    wire N__11288;
    wire N__11287;
    wire N__11284;
    wire N__11281;
    wire N__11278;
    wire N__11275;
    wire N__11272;
    wire N__11269;
    wire N__11266;
    wire N__11261;
    wire N__11256;
    wire N__11253;
    wire N__11250;
    wire N__11247;
    wire N__11244;
    wire N__11243;
    wire N__11242;
    wire N__11241;
    wire N__11238;
    wire N__11235;
    wire N__11232;
    wire N__11229;
    wire N__11226;
    wire N__11223;
    wire N__11218;
    wire N__11215;
    wire N__11212;
    wire N__11209;
    wire N__11202;
    wire N__11199;
    wire N__11196;
    wire N__11193;
    wire N__11190;
    wire N__11187;
    wire N__11184;
    wire N__11181;
    wire N__11178;
    wire N__11175;
    wire N__11172;
    wire N__11171;
    wire N__11168;
    wire N__11165;
    wire N__11162;
    wire N__11157;
    wire N__11156;
    wire N__11153;
    wire N__11150;
    wire N__11147;
    wire N__11144;
    wire N__11139;
    wire N__11136;
    wire N__11135;
    wire N__11132;
    wire N__11129;
    wire N__11126;
    wire N__11121;
    wire N__11118;
    wire N__11115;
    wire N__11112;
    wire N__11109;
    wire N__11106;
    wire N__11103;
    wire N__11100;
    wire N__11097;
    wire N__11094;
    wire N__11091;
    wire N__11088;
    wire N__11085;
    wire N__11082;
    wire N__11079;
    wire N__11078;
    wire N__11075;
    wire N__11072;
    wire N__11069;
    wire N__11064;
    wire N__11061;
    wire N__11060;
    wire N__11059;
    wire N__11056;
    wire N__11055;
    wire N__11054;
    wire N__11053;
    wire N__11052;
    wire N__11051;
    wire N__11042;
    wire N__11033;
    wire N__11030;
    wire N__11025;
    wire N__11022;
    wire N__11019;
    wire N__11016;
    wire N__11013;
    wire N__11010;
    wire N__11007;
    wire N__11004;
    wire N__11001;
    wire N__10998;
    wire N__10995;
    wire N__10992;
    wire N__10989;
    wire N__10986;
    wire N__10983;
    wire N__10980;
    wire N__10977;
    wire N__10974;
    wire N__10971;
    wire N__10968;
    wire N__10965;
    wire N__10962;
    wire N__10961;
    wire N__10958;
    wire N__10955;
    wire N__10952;
    wire N__10949;
    wire N__10948;
    wire N__10943;
    wire N__10940;
    wire N__10935;
    wire N__10932;
    wire N__10929;
    wire N__10926;
    wire N__10923;
    wire N__10920;
    wire N__10917;
    wire N__10914;
    wire N__10911;
    wire N__10908;
    wire N__10905;
    wire N__10902;
    wire N__10899;
    wire N__10896;
    wire N__10893;
    wire N__10890;
    wire N__10889;
    wire N__10886;
    wire N__10883;
    wire N__10882;
    wire N__10879;
    wire N__10876;
    wire N__10873;
    wire N__10870;
    wire N__10867;
    wire N__10864;
    wire N__10857;
    wire N__10854;
    wire N__10853;
    wire N__10852;
    wire N__10849;
    wire N__10846;
    wire N__10843;
    wire N__10840;
    wire N__10837;
    wire N__10834;
    wire N__10827;
    wire N__10824;
    wire N__10821;
    wire N__10818;
    wire N__10815;
    wire N__10812;
    wire N__10809;
    wire N__10806;
    wire N__10803;
    wire N__10800;
    wire N__10797;
    wire N__10794;
    wire N__10791;
    wire N__10790;
    wire N__10787;
    wire N__10784;
    wire N__10779;
    wire N__10776;
    wire N__10773;
    wire N__10770;
    wire N__10767;
    wire N__10766;
    wire N__10763;
    wire N__10762;
    wire N__10759;
    wire N__10756;
    wire N__10753;
    wire N__10750;
    wire N__10743;
    wire N__10742;
    wire N__10737;
    wire N__10734;
    wire N__10731;
    wire N__10728;
    wire N__10725;
    wire N__10724;
    wire N__10721;
    wire N__10720;
    wire N__10717;
    wire N__10714;
    wire N__10711;
    wire N__10708;
    wire N__10701;
    wire N__10700;
    wire N__10695;
    wire N__10692;
    wire N__10689;
    wire N__10686;
    wire N__10685;
    wire N__10680;
    wire N__10677;
    wire N__10674;
    wire N__10673;
    wire N__10668;
    wire N__10665;
    wire N__10662;
    wire N__10659;
    wire N__10656;
    wire N__10653;
    wire N__10650;
    wire N__10647;
    wire N__10644;
    wire N__10641;
    wire N__10638;
    wire N__10635;
    wire N__10632;
    wire N__10629;
    wire N__10626;
    wire N__10623;
    wire N__10620;
    wire N__10617;
    wire N__10614;
    wire N__10611;
    wire N__10608;
    wire N__10605;
    wire N__10602;
    wire N__10599;
    wire N__10596;
    wire N__10593;
    wire N__10590;
    wire N__10587;
    wire N__10584;
    wire N__10581;
    wire N__10578;
    wire N__10575;
    wire N__10572;
    wire N__10569;
    wire N__10566;
    wire N__10563;
    wire N__10560;
    wire N__10557;
    wire N__10554;
    wire N__10551;
    wire N__10548;
    wire N__10547;
    wire N__10546;
    wire N__10545;
    wire N__10544;
    wire N__10543;
    wire N__10540;
    wire N__10539;
    wire N__10538;
    wire N__10537;
    wire N__10536;
    wire N__10535;
    wire N__10534;
    wire N__10533;
    wire N__10530;
    wire N__10527;
    wire N__10526;
    wire N__10523;
    wire N__10516;
    wire N__10513;
    wire N__10510;
    wire N__10509;
    wire N__10504;
    wire N__10503;
    wire N__10502;
    wire N__10501;
    wire N__10500;
    wire N__10499;
    wire N__10498;
    wire N__10495;
    wire N__10492;
    wire N__10491;
    wire N__10490;
    wire N__10481;
    wire N__10476;
    wire N__10475;
    wire N__10472;
    wire N__10469;
    wire N__10468;
    wire N__10465;
    wire N__10462;
    wire N__10453;
    wire N__10450;
    wire N__10447;
    wire N__10440;
    wire N__10437;
    wire N__10434;
    wire N__10431;
    wire N__10428;
    wire N__10423;
    wire N__10420;
    wire N__10417;
    wire N__10412;
    wire N__10389;
    wire N__10386;
    wire N__10383;
    wire N__10380;
    wire N__10377;
    wire N__10376;
    wire N__10373;
    wire N__10370;
    wire N__10365;
    wire N__10362;
    wire N__10359;
    wire N__10358;
    wire N__10355;
    wire N__10352;
    wire N__10347;
    wire N__10346;
    wire N__10341;
    wire N__10338;
    wire N__10335;
    wire N__10332;
    wire N__10329;
    wire N__10326;
    wire N__10323;
    wire N__10320;
    wire N__10317;
    wire N__10316;
    wire N__10313;
    wire N__10308;
    wire N__10305;
    wire N__10302;
    wire N__10299;
    wire N__10296;
    wire N__10293;
    wire N__10290;
    wire N__10287;
    wire N__10284;
    wire N__10281;
    wire N__10280;
    wire N__10277;
    wire N__10274;
    wire N__10273;
    wire N__10268;
    wire N__10265;
    wire N__10264;
    wire N__10263;
    wire N__10260;
    wire N__10257;
    wire N__10254;
    wire N__10251;
    wire N__10242;
    wire N__10239;
    wire N__10236;
    wire N__10233;
    wire N__10230;
    wire N__10229;
    wire N__10226;
    wire N__10223;
    wire N__10222;
    wire N__10221;
    wire N__10220;
    wire N__10217;
    wire N__10214;
    wire N__10211;
    wire N__10208;
    wire N__10205;
    wire N__10194;
    wire N__10191;
    wire N__10188;
    wire N__10187;
    wire N__10184;
    wire N__10183;
    wire N__10180;
    wire N__10177;
    wire N__10174;
    wire N__10171;
    wire N__10170;
    wire N__10169;
    wire N__10166;
    wire N__10163;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10143;
    wire N__10140;
    wire N__10137;
    wire N__10136;
    wire N__10133;
    wire N__10130;
    wire N__10129;
    wire N__10126;
    wire N__10123;
    wire N__10120;
    wire N__10119;
    wire N__10118;
    wire N__10115;
    wire N__10112;
    wire N__10109;
    wire N__10106;
    wire N__10103;
    wire N__10092;
    wire N__10089;
    wire N__10086;
    wire N__10083;
    wire N__10082;
    wire N__10079;
    wire N__10076;
    wire N__10073;
    wire N__10070;
    wire N__10067;
    wire N__10064;
    wire N__10059;
    wire N__10058;
    wire N__10055;
    wire N__10054;
    wire N__10051;
    wire N__10048;
    wire N__10045;
    wire N__10044;
    wire N__10037;
    wire N__10034;
    wire N__10031;
    wire N__10028;
    wire N__10023;
    wire N__10020;
    wire N__10017;
    wire N__10014;
    wire N__10013;
    wire N__10012;
    wire N__10009;
    wire N__10006;
    wire N__10003;
    wire N__10000;
    wire N__9997;
    wire N__9994;
    wire N__9989;
    wire N__9988;
    wire N__9985;
    wire N__9982;
    wire N__9979;
    wire N__9972;
    wire N__9969;
    wire N__9966;
    wire N__9965;
    wire N__9964;
    wire N__9963;
    wire N__9962;
    wire N__9961;
    wire N__9960;
    wire N__9959;
    wire N__9958;
    wire N__9955;
    wire N__9954;
    wire N__9953;
    wire N__9950;
    wire N__9947;
    wire N__9946;
    wire N__9945;
    wire N__9934;
    wire N__9927;
    wire N__9918;
    wire N__9917;
    wire N__9914;
    wire N__9913;
    wire N__9912;
    wire N__9911;
    wire N__9910;
    wire N__9909;
    wire N__9908;
    wire N__9905;
    wire N__9900;
    wire N__9895;
    wire N__9892;
    wire N__9887;
    wire N__9884;
    wire N__9879;
    wire N__9872;
    wire N__9869;
    wire N__9858;
    wire N__9855;
    wire N__9852;
    wire N__9849;
    wire N__9846;
    wire N__9845;
    wire N__9842;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9828;
    wire N__9827;
    wire N__9824;
    wire N__9821;
    wire N__9818;
    wire N__9815;
    wire N__9814;
    wire N__9811;
    wire N__9808;
    wire N__9805;
    wire N__9798;
    wire N__9795;
    wire N__9792;
    wire N__9789;
    wire N__9786;
    wire N__9783;
    wire N__9780;
    wire N__9777;
    wire N__9774;
    wire N__9773;
    wire N__9772;
    wire N__9769;
    wire N__9766;
    wire N__9763;
    wire N__9760;
    wire N__9757;
    wire N__9754;
    wire N__9751;
    wire N__9748;
    wire N__9745;
    wire N__9742;
    wire N__9735;
    wire N__9732;
    wire N__9729;
    wire N__9726;
    wire N__9725;
    wire N__9722;
    wire N__9719;
    wire N__9718;
    wire N__9717;
    wire N__9714;
    wire N__9711;
    wire N__9708;
    wire N__9705;
    wire N__9704;
    wire N__9701;
    wire N__9698;
    wire N__9695;
    wire N__9692;
    wire N__9689;
    wire N__9678;
    wire N__9675;
    wire N__9672;
    wire N__9669;
    wire N__9666;
    wire N__9665;
    wire N__9662;
    wire N__9659;
    wire N__9658;
    wire N__9653;
    wire N__9650;
    wire N__9649;
    wire N__9648;
    wire N__9645;
    wire N__9642;
    wire N__9639;
    wire N__9636;
    wire N__9627;
    wire N__9624;
    wire N__9621;
    wire N__9618;
    wire N__9615;
    wire N__9614;
    wire N__9611;
    wire N__9608;
    wire N__9607;
    wire N__9606;
    wire N__9605;
    wire N__9602;
    wire N__9599;
    wire N__9596;
    wire N__9593;
    wire N__9590;
    wire N__9579;
    wire N__9578;
    wire N__9575;
    wire N__9572;
    wire N__9567;
    wire N__9564;
    wire N__9561;
    wire N__9558;
    wire N__9555;
    wire N__9554;
    wire N__9551;
    wire N__9548;
    wire N__9543;
    wire N__9542;
    wire N__9539;
    wire N__9536;
    wire N__9531;
    wire N__9528;
    wire N__9527;
    wire N__9526;
    wire N__9525;
    wire N__9524;
    wire N__9521;
    wire N__9516;
    wire N__9511;
    wire N__9504;
    wire N__9503;
    wire N__9502;
    wire N__9499;
    wire N__9494;
    wire N__9491;
    wire N__9488;
    wire N__9485;
    wire N__9482;
    wire N__9479;
    wire N__9476;
    wire N__9473;
    wire N__9470;
    wire N__9467;
    wire N__9462;
    wire N__9461;
    wire N__9460;
    wire N__9455;
    wire N__9454;
    wire N__9453;
    wire N__9450;
    wire N__9447;
    wire N__9442;
    wire N__9435;
    wire N__9432;
    wire N__9429;
    wire N__9426;
    wire N__9423;
    wire N__9420;
    wire N__9417;
    wire N__9414;
    wire N__9413;
    wire N__9412;
    wire N__9411;
    wire N__9408;
    wire N__9401;
    wire N__9400;
    wire N__9399;
    wire N__9398;
    wire N__9397;
    wire N__9396;
    wire N__9395;
    wire N__9394;
    wire N__9393;
    wire N__9390;
    wire N__9387;
    wire N__9382;
    wire N__9381;
    wire N__9374;
    wire N__9367;
    wire N__9360;
    wire N__9357;
    wire N__9348;
    wire N__9345;
    wire N__9342;
    wire N__9339;
    wire N__9336;
    wire N__9333;
    wire N__9330;
    wire N__9327;
    wire N__9324;
    wire N__9321;
    wire N__9318;
    wire N__9315;
    wire N__9312;
    wire N__9309;
    wire N__9306;
    wire N__9303;
    wire N__9302;
    wire N__9301;
    wire N__9300;
    wire N__9299;
    wire N__9298;
    wire N__9297;
    wire N__9296;
    wire N__9295;
    wire N__9292;
    wire N__9287;
    wire N__9282;
    wire N__9279;
    wire N__9274;
    wire N__9271;
    wire N__9268;
    wire N__9263;
    wire N__9252;
    wire N__9249;
    wire N__9246;
    wire N__9243;
    wire N__9240;
    wire N__9239;
    wire N__9236;
    wire N__9235;
    wire N__9232;
    wire N__9229;
    wire N__9226;
    wire N__9219;
    wire N__9216;
    wire N__9213;
    wire N__9212;
    wire N__9211;
    wire N__9210;
    wire N__9207;
    wire N__9204;
    wire N__9201;
    wire N__9198;
    wire N__9195;
    wire N__9192;
    wire N__9183;
    wire N__9182;
    wire N__9179;
    wire N__9178;
    wire N__9177;
    wire N__9174;
    wire N__9173;
    wire N__9168;
    wire N__9165;
    wire N__9162;
    wire N__9159;
    wire N__9156;
    wire N__9149;
    wire N__9144;
    wire N__9141;
    wire N__9140;
    wire N__9139;
    wire N__9136;
    wire N__9131;
    wire N__9126;
    wire N__9123;
    wire N__9120;
    wire N__9119;
    wire N__9116;
    wire N__9111;
    wire N__9108;
    wire N__9107;
    wire N__9106;
    wire N__9103;
    wire N__9102;
    wire N__9101;
    wire N__9100;
    wire N__9099;
    wire N__9096;
    wire N__9093;
    wire N__9090;
    wire N__9083;
    wire N__9080;
    wire N__9069;
    wire N__9068;
    wire N__9067;
    wire N__9064;
    wire N__9061;
    wire N__9060;
    wire N__9059;
    wire N__9058;
    wire N__9055;
    wire N__9050;
    wire N__9043;
    wire N__9036;
    wire N__9033;
    wire N__9030;
    wire N__9029;
    wire N__9026;
    wire N__9023;
    wire N__9020;
    wire N__9017;
    wire N__9014;
    wire N__9011;
    wire N__9008;
    wire N__9005;
    wire N__9002;
    wire N__8999;
    wire N__8998;
    wire N__8995;
    wire N__8992;
    wire N__8989;
    wire N__8982;
    wire N__8979;
    wire N__8976;
    wire N__8973;
    wire N__8972;
    wire N__8969;
    wire N__8966;
    wire N__8963;
    wire N__8960;
    wire N__8955;
    wire N__8954;
    wire N__8953;
    wire N__8952;
    wire N__8951;
    wire N__8950;
    wire N__8947;
    wire N__8944;
    wire N__8939;
    wire N__8936;
    wire N__8933;
    wire N__8930;
    wire N__8927;
    wire N__8924;
    wire N__8921;
    wire N__8910;
    wire N__8909;
    wire N__8908;
    wire N__8905;
    wire N__8904;
    wire N__8903;
    wire N__8900;
    wire N__8895;
    wire N__8894;
    wire N__8891;
    wire N__8888;
    wire N__8883;
    wire N__8880;
    wire N__8871;
    wire N__8870;
    wire N__8869;
    wire N__8868;
    wire N__8867;
    wire N__8866;
    wire N__8863;
    wire N__8858;
    wire N__8855;
    wire N__8852;
    wire N__8849;
    wire N__8844;
    wire N__8841;
    wire N__8832;
    wire N__8831;
    wire N__8830;
    wire N__8829;
    wire N__8826;
    wire N__8821;
    wire N__8820;
    wire N__8817;
    wire N__8814;
    wire N__8811;
    wire N__8808;
    wire N__8799;
    wire N__8798;
    wire N__8795;
    wire N__8794;
    wire N__8793;
    wire N__8790;
    wire N__8789;
    wire N__8786;
    wire N__8781;
    wire N__8778;
    wire N__8775;
    wire N__8772;
    wire N__8769;
    wire N__8764;
    wire N__8757;
    wire N__8754;
    wire N__8753;
    wire N__8750;
    wire N__8749;
    wire N__8748;
    wire N__8747;
    wire N__8744;
    wire N__8739;
    wire N__8738;
    wire N__8735;
    wire N__8732;
    wire N__8729;
    wire N__8726;
    wire N__8723;
    wire N__8712;
    wire N__8709;
    wire N__8706;
    wire N__8703;
    wire N__8700;
    wire N__8697;
    wire N__8694;
    wire N__8693;
    wire N__8692;
    wire N__8691;
    wire N__8690;
    wire N__8689;
    wire N__8688;
    wire N__8683;
    wire N__8680;
    wire N__8675;
    wire N__8670;
    wire N__8667;
    wire N__8658;
    wire N__8655;
    wire N__8652;
    wire N__8649;
    wire N__8646;
    wire N__8643;
    wire N__8640;
    wire N__8637;
    wire N__8634;
    wire N__8631;
    wire N__8628;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8620;
    wire N__8617;
    wire N__8614;
    wire N__8611;
    wire N__8604;
    wire N__8601;
    wire N__8598;
    wire N__8595;
    wire N__8592;
    wire N__8589;
    wire N__8586;
    wire N__8583;
    wire N__8580;
    wire N__8577;
    wire N__8574;
    wire N__8571;
    wire N__8568;
    wire N__8565;
    wire N__8562;
    wire N__8559;
    wire N__8556;
    wire N__8553;
    wire N__8550;
    wire N__8547;
    wire N__8544;
    wire N__8541;
    wire N__8538;
    wire N__8537;
    wire N__8536;
    wire N__8535;
    wire N__8534;
    wire N__8533;
    wire N__8532;
    wire N__8531;
    wire N__8528;
    wire N__8525;
    wire N__8524;
    wire N__8521;
    wire N__8520;
    wire N__8517;
    wire N__8516;
    wire N__8513;
    wire N__8512;
    wire N__8509;
    wire N__8508;
    wire N__8505;
    wire N__8504;
    wire N__8503;
    wire N__8502;
    wire N__8501;
    wire N__8500;
    wire N__8499;
    wire N__8498;
    wire N__8497;
    wire N__8484;
    wire N__8469;
    wire N__8468;
    wire N__8467;
    wire N__8464;
    wire N__8463;
    wire N__8460;
    wire N__8459;
    wire N__8456;
    wire N__8455;
    wire N__8452;
    wire N__8451;
    wire N__8450;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8440;
    wire N__8439;
    wire N__8436;
    wire N__8435;
    wire N__8430;
    wire N__8427;
    wire N__8410;
    wire N__8407;
    wire N__8392;
    wire N__8389;
    wire N__8388;
    wire N__8381;
    wire N__8376;
    wire N__8373;
    wire N__8370;
    wire N__8365;
    wire N__8362;
    wire N__8359;
    wire N__8352;
    wire N__8351;
    wire N__8350;
    wire N__8349;
    wire N__8348;
    wire N__8345;
    wire N__8342;
    wire N__8341;
    wire N__8340;
    wire N__8337;
    wire N__8336;
    wire N__8335;
    wire N__8334;
    wire N__8333;
    wire N__8330;
    wire N__8329;
    wire N__8322;
    wire N__8321;
    wire N__8320;
    wire N__8319;
    wire N__8318;
    wire N__8317;
    wire N__8316;
    wire N__8315;
    wire N__8312;
    wire N__8309;
    wire N__8306;
    wire N__8303;
    wire N__8302;
    wire N__8301;
    wire N__8298;
    wire N__8293;
    wire N__8288;
    wire N__8287;
    wire N__8286;
    wire N__8285;
    wire N__8284;
    wire N__8283;
    wire N__8282;
    wire N__8281;
    wire N__8280;
    wire N__8279;
    wire N__8278;
    wire N__8275;
    wire N__8270;
    wire N__8265;
    wire N__8256;
    wire N__8253;
    wire N__8248;
    wire N__8245;
    wire N__8242;
    wire N__8235;
    wire N__8220;
    wire N__8217;
    wire N__8212;
    wire N__8207;
    wire N__8202;
    wire N__8199;
    wire N__8194;
    wire N__8183;
    wire N__8178;
    wire N__8171;
    wire N__8166;
    wire N__8163;
    wire N__8160;
    wire N__8157;
    wire N__8154;
    wire N__8151;
    wire N__8148;
    wire N__8147;
    wire N__8146;
    wire N__8145;
    wire N__8144;
    wire N__8141;
    wire N__8140;
    wire N__8139;
    wire N__8138;
    wire N__8137;
    wire N__8134;
    wire N__8131;
    wire N__8128;
    wire N__8125;
    wire N__8124;
    wire N__8123;
    wire N__8122;
    wire N__8121;
    wire N__8120;
    wire N__8119;
    wire N__8116;
    wire N__8115;
    wire N__8114;
    wire N__8111;
    wire N__8096;
    wire N__8091;
    wire N__8088;
    wire N__8085;
    wire N__8082;
    wire N__8079;
    wire N__8078;
    wire N__8077;
    wire N__8074;
    wire N__8071;
    wire N__8070;
    wire N__8065;
    wire N__8060;
    wire N__8047;
    wire N__8042;
    wire N__8041;
    wire N__8040;
    wire N__8037;
    wire N__8034;
    wire N__8031;
    wire N__8026;
    wire N__8021;
    wire N__8010;
    wire N__8009;
    wire N__8006;
    wire N__8003;
    wire N__8002;
    wire N__7999;
    wire N__7996;
    wire N__7993;
    wire N__7988;
    wire N__7983;
    wire N__7980;
    wire N__7977;
    wire N__7974;
    wire N__7971;
    wire N__7968;
    wire N__7965;
    wire N__7962;
    wire N__7959;
    wire N__7958;
    wire N__7955;
    wire N__7952;
    wire N__7947;
    wire N__7944;
    wire N__7941;
    wire N__7938;
    wire N__7935;
    wire N__7932;
    wire N__7929;
    wire N__7926;
    wire N__7923;
    wire N__7920;
    wire N__7917;
    wire N__7914;
    wire N__7911;
    wire N__7908;
    wire N__7905;
    wire N__7902;
    wire N__7899;
    wire N__7896;
    wire N__7893;
    wire N__7892;
    wire N__7891;
    wire N__7886;
    wire N__7883;
    wire N__7880;
    wire N__7875;
    wire N__7872;
    wire N__7869;
    wire N__7866;
    wire N__7863;
    wire N__7860;
    wire N__7857;
    wire N__7854;
    wire N__7851;
    wire N__7848;
    wire N__7845;
    wire N__7842;
    wire N__7839;
    wire N__7836;
    wire N__7833;
    wire N__7832;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7812;
    wire N__7809;
    wire N__7806;
    wire N__7805;
    wire N__7804;
    wire N__7803;
    wire N__7802;
    wire N__7801;
    wire N__7800;
    wire N__7795;
    wire N__7790;
    wire N__7783;
    wire N__7776;
    wire N__7775;
    wire N__7772;
    wire N__7769;
    wire N__7766;
    wire N__7761;
    wire N__7760;
    wire N__7759;
    wire N__7756;
    wire N__7755;
    wire N__7752;
    wire N__7751;
    wire N__7748;
    wire N__7747;
    wire N__7746;
    wire N__7743;
    wire N__7740;
    wire N__7735;
    wire N__7728;
    wire N__7719;
    wire N__7718;
    wire N__7717;
    wire N__7716;
    wire N__7715;
    wire N__7714;
    wire N__7713;
    wire N__7710;
    wire N__7705;
    wire N__7696;
    wire N__7689;
    wire N__7686;
    wire N__7683;
    wire N__7680;
    wire N__7677;
    wire N__7674;
    wire N__7671;
    wire N__7668;
    wire N__7667;
    wire N__7664;
    wire N__7661;
    wire N__7658;
    wire N__7655;
    wire N__7650;
    wire N__7647;
    wire N__7646;
    wire N__7643;
    wire N__7640;
    wire N__7635;
    wire N__7634;
    wire N__7631;
    wire N__7628;
    wire N__7623;
    wire N__7620;
    wire N__7617;
    wire N__7616;
    wire N__7613;
    wire N__7612;
    wire N__7609;
    wire N__7606;
    wire N__7603;
    wire N__7600;
    wire N__7593;
    wire N__7590;
    wire N__7587;
    wire N__7584;
    wire N__7583;
    wire N__7580;
    wire N__7577;
    wire N__7574;
    wire N__7571;
    wire N__7568;
    wire N__7565;
    wire N__7560;
    wire N__7557;
    wire N__7554;
    wire N__7551;
    wire N__7548;
    wire N__7547;
    wire N__7544;
    wire N__7541;
    wire N__7538;
    wire N__7535;
    wire N__7530;
    wire N__7527;
    wire N__7524;
    wire N__7521;
    wire N__7518;
    wire N__7515;
    wire N__7512;
    wire N__7509;
    wire N__7506;
    wire N__7503;
    wire N__7500;
    wire N__7499;
    wire N__7496;
    wire N__7495;
    wire N__7492;
    wire N__7489;
    wire N__7486;
    wire N__7483;
    wire N__7478;
    wire N__7475;
    wire N__7472;
    wire N__7469;
    wire N__7466;
    wire N__7461;
    wire N__7458;
    wire N__7457;
    wire N__7456;
    wire N__7455;
    wire N__7454;
    wire N__7453;
    wire N__7450;
    wire N__7447;
    wire N__7440;
    wire N__7437;
    wire N__7428;
    wire N__7427;
    wire N__7424;
    wire N__7421;
    wire N__7416;
    wire N__7415;
    wire N__7414;
    wire N__7413;
    wire N__7412;
    wire N__7407;
    wire N__7406;
    wire N__7403;
    wire N__7398;
    wire N__7395;
    wire N__7392;
    wire N__7391;
    wire N__7390;
    wire N__7387;
    wire N__7380;
    wire N__7375;
    wire N__7368;
    wire N__7365;
    wire N__7364;
    wire N__7363;
    wire N__7362;
    wire N__7361;
    wire N__7360;
    wire N__7359;
    wire N__7358;
    wire N__7355;
    wire N__7350;
    wire N__7349;
    wire N__7348;
    wire N__7341;
    wire N__7336;
    wire N__7333;
    wire N__7330;
    wire N__7325;
    wire N__7320;
    wire N__7317;
    wire N__7308;
    wire N__7307;
    wire N__7306;
    wire N__7303;
    wire N__7300;
    wire N__7297;
    wire N__7294;
    wire N__7289;
    wire N__7288;
    wire N__7287;
    wire N__7286;
    wire N__7285;
    wire N__7284;
    wire N__7283;
    wire N__7282;
    wire N__7281;
    wire N__7280;
    wire N__7277;
    wire N__7274;
    wire N__7267;
    wire N__7262;
    wire N__7253;
    wire N__7242;
    wire N__7239;
    wire N__7236;
    wire N__7235;
    wire N__7230;
    wire N__7227;
    wire N__7226;
    wire N__7221;
    wire N__7218;
    wire N__7215;
    wire N__7212;
    wire N__7209;
    wire N__7206;
    wire N__7203;
    wire N__7200;
    wire N__7199;
    wire N__7196;
    wire N__7193;
    wire N__7188;
    wire N__7187;
    wire N__7184;
    wire N__7181;
    wire N__7176;
    wire N__7173;
    wire N__7172;
    wire N__7169;
    wire N__7166;
    wire N__7161;
    wire N__7160;
    wire N__7157;
    wire N__7154;
    wire N__7149;
    wire N__7148;
    wire N__7145;
    wire N__7142;
    wire N__7137;
    wire N__7134;
    wire N__7133;
    wire N__7130;
    wire N__7129;
    wire N__7126;
    wire N__7123;
    wire N__7120;
    wire N__7113;
    wire N__7110;
    wire N__7107;
    wire N__7106;
    wire N__7103;
    wire N__7100;
    wire N__7095;
    wire N__7092;
    wire N__7089;
    wire N__7086;
    wire N__7085;
    wire N__7082;
    wire N__7081;
    wire N__7080;
    wire N__7075;
    wire N__7072;
    wire N__7069;
    wire N__7064;
    wire N__7061;
    wire N__7058;
    wire N__7057;
    wire N__7054;
    wire N__7051;
    wire N__7048;
    wire N__7041;
    wire N__7038;
    wire N__7035;
    wire N__7034;
    wire N__7031;
    wire N__7028;
    wire N__7027;
    wire N__7024;
    wire N__7019;
    wire N__7018;
    wire N__7017;
    wire N__7016;
    wire N__7015;
    wire N__7012;
    wire N__7009;
    wire N__7002;
    wire N__6999;
    wire N__6992;
    wire N__6989;
    wire N__6986;
    wire N__6981;
    wire N__6980;
    wire N__6977;
    wire N__6974;
    wire N__6971;
    wire N__6966;
    wire N__6965;
    wire N__6964;
    wire N__6961;
    wire N__6956;
    wire N__6951;
    wire N__6948;
    wire N__6945;
    wire N__6944;
    wire N__6943;
    wire N__6942;
    wire N__6939;
    wire N__6934;
    wire N__6931;
    wire N__6924;
    wire N__6923;
    wire N__6922;
    wire N__6921;
    wire N__6918;
    wire N__6913;
    wire N__6910;
    wire N__6903;
    wire N__6900;
    wire N__6899;
    wire N__6896;
    wire N__6893;
    wire N__6888;
    wire N__6887;
    wire N__6884;
    wire N__6881;
    wire N__6876;
    wire N__6875;
    wire N__6872;
    wire N__6869;
    wire N__6864;
    wire N__6861;
    wire N__6860;
    wire N__6857;
    wire N__6854;
    wire N__6851;
    wire N__6846;
    wire N__6843;
    wire N__6842;
    wire N__6839;
    wire N__6836;
    wire N__6831;
    wire N__6828;
    wire N__6825;
    wire N__6824;
    wire N__6821;
    wire N__6818;
    wire N__6813;
    wire N__6812;
    wire N__6809;
    wire N__6806;
    wire N__6801;
    wire N__6798;
    wire N__6797;
    wire N__6794;
    wire N__6791;
    wire N__6788;
    wire N__6783;
    wire N__6780;
    wire N__6779;
    wire N__6776;
    wire N__6773;
    wire N__6768;
    wire N__6765;
    wire N__6764;
    wire N__6763;
    wire N__6760;
    wire N__6757;
    wire N__6756;
    wire N__6753;
    wire N__6748;
    wire N__6745;
    wire N__6738;
    wire N__6735;
    wire N__6732;
    wire N__6729;
    wire N__6728;
    wire N__6725;
    wire N__6722;
    wire N__6717;
    wire N__6714;
    wire N__6711;
    wire N__6708;
    wire N__6707;
    wire N__6704;
    wire N__6701;
    wire N__6696;
    wire N__6693;
    wire N__6690;
    wire N__6689;
    wire N__6686;
    wire N__6683;
    wire N__6678;
    wire N__6675;
    wire N__6672;
    wire N__6669;
    wire N__6666;
    wire N__6663;
    wire N__6660;
    wire N__6657;
    wire N__6654;
    wire N__6651;
    wire N__6648;
    wire N__6645;
    wire N__6644;
    wire N__6641;
    wire N__6638;
    wire N__6633;
    wire N__6632;
    wire N__6629;
    wire N__6624;
    wire N__6621;
    wire N__6618;
    wire N__6615;
    wire N__6614;
    wire N__6613;
    wire N__6612;
    wire N__6611;
    wire N__6610;
    wire N__6609;
    wire N__6604;
    wire N__6601;
    wire N__6600;
    wire N__6597;
    wire N__6596;
    wire N__6595;
    wire N__6592;
    wire N__6589;
    wire N__6586;
    wire N__6583;
    wire N__6578;
    wire N__6571;
    wire N__6568;
    wire N__6565;
    wire N__6552;
    wire N__6551;
    wire N__6550;
    wire N__6549;
    wire N__6548;
    wire N__6547;
    wire N__6546;
    wire N__6545;
    wire N__6538;
    wire N__6533;
    wire N__6528;
    wire N__6525;
    wire N__6524;
    wire N__6523;
    wire N__6522;
    wire N__6519;
    wire N__6512;
    wire N__6507;
    wire N__6504;
    wire N__6497;
    wire N__6492;
    wire N__6489;
    wire N__6486;
    wire N__6483;
    wire N__6480;
    wire N__6477;
    wire N__6474;
    wire N__6471;
    wire N__6470;
    wire N__6467;
    wire N__6464;
    wire N__6459;
    wire N__6456;
    wire N__6453;
    wire N__6450;
    wire N__6447;
    wire N__6444;
    wire N__6443;
    wire N__6440;
    wire N__6437;
    wire N__6432;
    wire N__6429;
    wire N__6426;
    wire N__6423;
    wire N__6420;
    wire N__6417;
    wire N__6416;
    wire N__6413;
    wire N__6412;
    wire N__6411;
    wire N__6408;
    wire N__6401;
    wire N__6396;
    wire N__6395;
    wire N__6394;
    wire N__6393;
    wire N__6386;
    wire N__6385;
    wire N__6384;
    wire N__6381;
    wire N__6378;
    wire N__6371;
    wire N__6366;
    wire N__6365;
    wire N__6364;
    wire N__6363;
    wire N__6360;
    wire N__6355;
    wire N__6352;
    wire N__6351;
    wire N__6346;
    wire N__6341;
    wire N__6336;
    wire N__6335;
    wire N__6334;
    wire N__6333;
    wire N__6332;
    wire N__6327;
    wire N__6320;
    wire N__6315;
    wire N__6314;
    wire N__6313;
    wire N__6312;
    wire N__6309;
    wire N__6306;
    wire N__6305;
    wire N__6302;
    wire N__6293;
    wire N__6288;
    wire N__6285;
    wire N__6282;
    wire N__6279;
    wire N__6276;
    wire N__6273;
    wire N__6270;
    wire N__6267;
    wire N__6266;
    wire N__6265;
    wire N__6262;
    wire N__6255;
    wire N__6252;
    wire N__6249;
    wire N__6246;
    wire N__6245;
    wire N__6244;
    wire N__6243;
    wire N__6234;
    wire N__6231;
    wire N__6228;
    wire N__6225;
    wire N__6222;
    wire N__6219;
    wire N__6216;
    wire N__6213;
    wire N__6210;
    wire N__6207;
    wire N__6204;
    wire N__6201;
    wire N__6198;
    wire N__6195;
    wire N__6192;
    wire N__6189;
    wire N__6186;
    wire N__6183;
    wire N__6180;
    wire N__6177;
    wire N__6176;
    wire N__6175;
    wire N__6172;
    wire N__6169;
    wire N__6166;
    wire N__6163;
    wire N__6156;
    wire N__6153;
    wire N__6150;
    wire N__6147;
    wire N__6146;
    wire N__6143;
    wire N__6142;
    wire N__6139;
    wire N__6136;
    wire N__6133;
    wire N__6126;
    wire N__6123;
    wire N__6120;
    wire N__6119;
    wire N__6118;
    wire N__6115;
    wire N__6112;
    wire N__6109;
    wire N__6102;
    wire N__6099;
    wire N__6096;
    wire N__6093;
    wire N__6092;
    wire N__6089;
    wire N__6088;
    wire N__6085;
    wire N__6082;
    wire N__6079;
    wire N__6072;
    wire N__6069;
    wire N__6066;
    wire N__6063;
    wire N__6060;
    wire N__6057;
    wire N__6054;
    wire N__6053;
    wire N__6052;
    wire N__6051;
    wire N__6050;
    wire N__6047;
    wire N__6044;
    wire N__6037;
    wire N__6030;
    wire N__6029;
    wire N__6028;
    wire N__6027;
    wire N__6026;
    wire N__6025;
    wire N__6024;
    wire N__6023;
    wire N__6020;
    wire N__6015;
    wire N__6012;
    wire N__6009;
    wire N__6004;
    wire N__6001;
    wire N__5996;
    wire N__5985;
    wire N__5982;
    wire N__5981;
    wire N__5980;
    wire N__5979;
    wire N__5978;
    wire N__5977;
    wire N__5976;
    wire N__5973;
    wire N__5970;
    wire N__5965;
    wire N__5958;
    wire N__5949;
    wire N__5948;
    wire N__5947;
    wire N__5944;
    wire N__5941;
    wire N__5938;
    wire N__5931;
    wire N__5930;
    wire N__5927;
    wire N__5924;
    wire N__5919;
    wire N__5916;
    wire N__5915;
    wire N__5912;
    wire N__5911;
    wire N__5908;
    wire N__5905;
    wire N__5902;
    wire N__5895;
    wire N__5894;
    wire N__5891;
    wire N__5890;
    wire N__5887;
    wire N__5884;
    wire N__5881;
    wire N__5874;
    wire N__5871;
    wire N__5868;
    wire N__5867;
    wire N__5864;
    wire N__5861;
    wire N__5858;
    wire N__5855;
    wire N__5850;
    wire N__5847;
    wire N__5844;
    wire N__5841;
    wire N__5838;
    wire N__5835;
    wire N__5834;
    wire N__5833;
    wire N__5826;
    wire N__5823;
    wire N__5820;
    wire N__5817;
    wire N__5814;
    wire N__5811;
    wire N__5810;
    wire N__5809;
    wire N__5806;
    wire N__5805;
    wire N__5802;
    wire N__5795;
    wire N__5790;
    wire N__5787;
    wire N__5784;
    wire N__5781;
    wire N__5778;
    wire N__5775;
    wire N__5772;
    wire N__5769;
    wire N__5766;
    wire N__5763;
    wire N__5760;
    wire N__5759;
    wire N__5754;
    wire N__5751;
    wire N__5748;
    wire N__5745;
    wire N__5742;
    wire N__5741;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5731;
    wire N__5724;
    wire N__5721;
    wire N__5718;
    wire N__5715;
    wire N__5714;
    wire N__5711;
    wire N__5710;
    wire N__5707;
    wire N__5704;
    wire N__5701;
    wire N__5694;
    wire N__5691;
    wire N__5688;
    wire N__5685;
    wire N__5684;
    wire N__5683;
    wire N__5680;
    wire N__5677;
    wire N__5674;
    wire N__5667;
    wire N__5664;
    wire N__5661;
    wire N__5658;
    wire N__5657;
    wire N__5654;
    wire N__5653;
    wire N__5650;
    wire N__5647;
    wire N__5644;
    wire N__5637;
    wire N__5634;
    wire N__5631;
    wire N__5628;
    wire N__5627;
    wire N__5626;
    wire N__5623;
    wire N__5620;
    wire N__5617;
    wire N__5610;
    wire N__5607;
    wire N__5604;
    wire N__5601;
    wire N__5600;
    wire N__5599;
    wire N__5596;
    wire N__5593;
    wire N__5590;
    wire N__5587;
    wire N__5584;
    wire N__5577;
    wire N__5574;
    wire N__5571;
    wire N__5568;
    wire N__5565;
    wire N__5562;
    wire N__5559;
    wire N__5556;
    wire N__5553;
    wire N__5550;
    wire N__5547;
    wire N__5544;
    wire N__5541;
    wire N__5538;
    wire N__5535;
    wire N__5532;
    wire N__5529;
    wire N__5526;
    wire N__5523;
    wire N__5520;
    wire N__5517;
    wire N__5514;
    wire N__5511;
    wire N__5508;
    wire N__5505;
    wire N__5502;
    wire N__5499;
    wire N__5496;
    wire N__5493;
    wire N__5490;
    wire N__5487;
    wire N__5484;
    wire N__5481;
    wire N__5478;
    wire N__5475;
    wire N__5472;
    wire N__5469;
    wire N__5466;
    wire N__5463;
    wire N__5460;
    wire N__5457;
    wire N__5454;
    wire N__5451;
    wire N__5448;
    wire N__5445;
    wire N__5442;
    wire N__5439;
    wire N__5436;
    wire N__5433;
    wire N__5430;
    wire N__5427;
    wire N__5424;
    wire N__5421;
    wire N__5418;
    wire N__5415;
    wire N__5412;
    wire N__5409;
    wire N__5406;
    wire N__5403;
    wire N__5400;
    wire N__5397;
    wire N__5394;
    wire N__5391;
    wire N__5388;
    wire N__5385;
    wire N__5382;
    wire N__5379;
    wire N__5376;
    wire N__5373;
    wire N__5370;
    wire N__5367;
    wire N__5364;
    wire N__5361;
    wire BTN_N_c;
    wire wTxRdData_3;
    wire wTxRdData_5;
    wire wTxRdData_2;
    wire wTxRdData_6;
    wire wTxRdData_7;
    wire wTxRdData_0;
    wire VCCG0;
    wire wTxRdData_4;
    wire wTxRdData_1;
    wire GNDG0;
    wire \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_3_cascade_ ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_11 ;
    wire bfn_10_16_0_;
    wire \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0 ;
    wire \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_awe3_cascade_ ;
    wire \DUT.fifo_rx_inst.un1_i11_i_cascade_ ;
    wire \DUT.fifo_rx_inst.un1_i11_i ;
    wire bfn_11_11_0_;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_0 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_1 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_3 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_2 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_3 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_4 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_5 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_7 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_6 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_7 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_8 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO ;
    wire bfn_11_12_0_;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_9 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_8 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_10 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_9 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_11 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_10 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_12 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_11 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_12 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_13 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_14 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_15 ;
    wire bfn_11_13_0_;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_16 ;
    wire \DUT.uart_inst0.recv_stateZ0Z_4 ;
    wire \DUT.uart_inst0.recv_state_ns_0_0_0_cascade_ ;
    wire \DUT.uart_inst0.N_50 ;
    wire \DUT.uart_inst0.recv_state_srsts_1_3_cascade_ ;
    wire \DUT.uart_inst0.recv_stateZ0Z_3 ;
    wire \DUT.fifo_rx_inst.N_88_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoCount_RNIK3G92Z0Z_1 ;
    wire \DUT.fifo_rx_inst.rFifoCountZ0Z_1 ;
    wire \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1Z0Z_0_cascade_ ;
    wire \DUT.fifo_rx_inst.N_97_cascade_ ;
    wire \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0 ;
    wire \DUT.fifo_rx_inst.N_97 ;
    wire \DUT.fifo_rx_inst.rFifoCountZ0Z_0 ;
    wire \DUT.wRcvd ;
    wire \DUT.fifo_rx_inst.rFifoCountZ0Z_2 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ1Z_1 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_3 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_2 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_1 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_9_cascade_ ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_15_cascade_ ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_17 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_12 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_13 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_14 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_15 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_16 ;
    wire \DUT.uart_inst0.N_46_cascade_ ;
    wire \DUT.uart_inst0.rx_countdown_3_0 ;
    wire \DUT.uart_inst0.rx_countdown_RNI8KQG9Z0Z_0_cascade_ ;
    wire \DUT.uart_inst0.rx_countdown_8_i_o2_2_2_cascade_ ;
    wire \DUT.uart_inst0.N_42_cascade_ ;
    wire bfn_12_14_0_;
    wire \DUT.uart_inst0.tx_clk_divider_cry_0 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_1 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_2 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_3 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_4 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_5 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_6 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_7 ;
    wire bfn_12_15_0_;
    wire \DUT.uart_inst0.tx_clk_divider_cry_8 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_9 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_10 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_11 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_12 ;
    wire \DUT.uart_inst0.N_12_cascade_ ;
    wire \DUT.uart_inst0.N_7_0_cascade_ ;
    wire \DUT.uart_inst0.rx_bits_remainingZ0Z_3 ;
    wire \DUT.uart_inst0.m5_0_1_cascade_ ;
    wire \DUT.uart_inst0.N_6_cascade_ ;
    wire \DUT.uart_inst0.rx_bits_remainingZ0Z_2 ;
    wire \DUT.fifo_rx_inst.un1_i11_2_i ;
    wire \DUT.fifo_rx_inst.un1_i11_2_i_cascade_ ;
    wire \DUT.fifo_rx_inst.N_88 ;
    wire \DUT.fifo_rx_inst.rWritePtrZ0Z_0 ;
    wire \DUT.fifo_rx_inst.rWritePtrZ0Z_1 ;
    wire \DUT.fifo_rx_inst.N_85 ;
    wire \DUT.uart_inst0.rx_bits_remainingZ0Z_1 ;
    wire \DUT.uart_inst0.m5_1_cascade_ ;
    wire \DUT.uart_inst0.N_6_0 ;
    wire wPllLocked_i;
    wire \DUT.uart_inst0.rx_clk_divider_1_5 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_5 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_6 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_6 ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_3 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_0_c_RNOZ0 ;
    wire bfn_13_12_0_;
    wire \DUT.uart_inst0.rx_countdownZ0Z_1 ;
    wire \DUT.uart_inst0.rx_countdown_RNICSMA4Z0Z_1 ;
    wire \DUT.uart_inst0.rx_countdown_3_1 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_0 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_1 ;
    wire \DUT.uart_inst0.rx_countdownZ1Z_3 ;
    wire \DUT.uart_inst0.rx_countdown_RNIEUMA4Z0Z_3 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_2 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_3 ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_5 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_4 ;
    wire \DUT.uart_inst0.rx_countdown_3_5 ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_4 ;
    wire \DUT.uart_inst0.rx_countdown_RNIFVMA4Z0Z_4 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_15 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_14 ;
    wire \DUT.uart_inst0.rx_countdown_RNIDTMA4Z0Z_2 ;
    wire \DUT.uart_inst0.N_47 ;
    wire \DUT.uart_inst0.N_68 ;
    wire \DUT.uart_inst0.recv_stateZ0Z_5 ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_2 ;
    wire \DUT.uart_inst0.rx_countdown_3_2 ;
    wire \DUT.uart_inst0.rx_countdown_3_3 ;
    wire \DUT.uart_inst0.rx_countdown_3_4 ;
    wire \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa_0_a2_0_a2_1_cascade_ ;
    wire \DUT.uart_inst0.rx_countdown_8_i_o2_2_2 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_12 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_7 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_13 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_6 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_8_cascade_ ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_4 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_3 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_5 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_2 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_9_cascade_ ;
    wire \DUT.uart_inst0.tx_countdown_3_0_cascade_ ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_11 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_10 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_9 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_8 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_1 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_7_cascade_ ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_0 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_10_cascade_ ;
    wire \DUT.uart_inst0.tx_clk_divider_1_sqmuxa_1_0_cascade_ ;
    wire \DUT.uart_inst0.tx_clk_divider_1_sqmuxa_1_i ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_5 ;
    wire \DUT.uart_inst0.g0_0_1_cascade_ ;
    wire \DUT.uart_inst0.rx_bits_remainingZ0Z_0 ;
    wire \DUT.uart_inst0.N_62_4 ;
    wire \DUT.uart_inst0.recv_stateZ0Z_1 ;
    wire \DUT.uart_inst0.recv_state_srsts_1_2_cascade_ ;
    wire \DUT.uart_inst0.N_42 ;
    wire \DUT.uart_inst0.recv_stateZ0Z_2 ;
    wire \DUT.uart_inst0.m5_0_0 ;
    wire \DUT.fifo_rx_inst.rFifoDataro_0 ;
    wire \DUT.fifo_rx_inst.rFifoDataro_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_7 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_6 ;
    wire \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa ;
    wire \DUT.uart_inst0.tx_bits_remaining_RNI5UON8Z0Z_3_cascade_ ;
    wire \DUT.uart_inst0.N_109_cascade_ ;
    wire \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIKK41CZ0_cascade_ ;
    wire \DUT.uart_inst0.N_109 ;
    wire \DUT.uart_inst0.tx_state_ns_i_i_a3_1_0 ;
    wire \DUT.uart_inst0.N_82 ;
    wire \DUT.uart_inst0.tx_countdown_3_cry_0_c_RNOZ0 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_3 ;
    wire bfn_14_14_0_;
    wire \DUT.uart_inst0.tx_countdown_3_cry_0 ;
    wire \DUT.uart_inst0.tx_countdown_RNI5L692Z0Z_2 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_2 ;
    wire \DUT.uart_inst0.tx_countdown_3_cry_1 ;
    wire \DUT.uart_inst0.tx_countdown_3_cry_2 ;
    wire \DUT.uart_inst0.tx_countdown_RNI7N692Z0Z_4 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_4 ;
    wire \DUT.uart_inst0.tx_countdown_3_cry_3 ;
    wire \DUT.uart_inst0.tx_countdown_3_axb_5 ;
    wire \DUT.uart_inst0.tx_countdown_3_cry_4 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_1 ;
    wire \DUT.uart_inst0.tx_countdown_RNI4K692Z0Z_1 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_10 ;
    wire \DUT.uart_inst0.tx_countdownZ1Z_3 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_8 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_9 ;
    wire \DUT.uart_inst0.tx_countdown_RNI6M692Z0Z_3 ;
    wire bfn_14_15_0_;
    wire \DUT.uart_inst0.un1_tx_bits_remaining_cry_0 ;
    wire \DUT.uart_inst0.un1_tx_bits_remaining_cry_1 ;
    wire \DUT.uart_inst0.un1_tx_bits_remaining_cry_2 ;
    wire P1A3_c;
    wire N_100_i;
    wire \DUT.fifo_rx_inst.rTxByte_52_1 ;
    wire \DUT.fifo_rx_inst.rTxByte_52_0_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1Z0Z_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_2 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_2 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_6 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_7 ;
    wire \DUT.fifo_rx_inst.rFifoData_awe1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_4 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_4 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_5 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_5 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_3 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_3 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_6 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_3 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_5 ;
    wire CONSTANT_ONE_NET;
    wire P1A1_c;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO ;
    wire \DUT.uart_inst0.recv_stateZ0Z_0 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_4 ;
    wire \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_3 ;
    wire \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_3_cascade_ ;
    wire P1A7_c;
    wire \DUT.uart_inst0.N_112 ;
    wire \DUT.uart_inst0.tx_out_6_iv_0_a3_1_1_cascade_ ;
    wire \DUT.uart_inst0.tx_out_6_iv_0_a3_1_sx_cascade_ ;
    wire \DUT.uart_inst0.N_113 ;
    wire \DUT.uart_inst0.tx_countdown_7_i_a3_0_sx_3_cascade_ ;
    wire \DUT.uart_inst0.N_116 ;
    wire \DUT.uart_inst0.N_76_i ;
    wire \DUT.uart_inst0.tx_countdown_3_2 ;
    wire \DUT.uart_inst0.tx_countdown_3_4 ;
    wire \DUT.uart_inst0.tx_countdown_3_1 ;
    wire \DUT.uart_inst0.tx_countdown_3_3 ;
    wire \DUT.uart_inst0.tx_countdown_3_0 ;
    wire \DUT.uart_inst0.N_77_cascade_ ;
    wire \DUT.uart_inst0.tx_countdown_3_5 ;
    wire \DUT.uart_inst0.tx_state_RNI9DTT5Z0Z_0_cascade_ ;
    wire \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIMJ5ECZ0 ;
    wire \DUT.uart_inst0.N_99_cascade_ ;
    wire \DUT.uart_inst0.un1_tx_bits_remaining_cry_0_c_RNOZ0 ;
    wire \DUT.tx_state_1 ;
    wire \DUT.uart_inst0.N_77 ;
    wire \DUT.uart_inst0.tx_bits_remaining_RNO_0Z0Z_3 ;
    wire \DUT.uart_inst0.tx_bits_remaining_RNIAIE4LZ0Z_1 ;
    wire \DUT.uart_inst0.tx_bits_remainingZ0Z_1 ;
    wire \DUT.uart_inst0.tx_bits_remainingZ0Z_0 ;
    wire \DUT.uart_inst0.N_124 ;
    wire \DUT.uart_inst0.tx_bits_remainingZ0Z_2 ;
    wire \DUT.uart_inst0.tx_bits_remaining_RNIBJE4LZ0Z_2 ;
    wire \DUT.uart_inst0.tx_bits_remainingZ0Z_3 ;
    wire \DUT.uart_inst0.N_96 ;
    wire \DUT.uart_inst0.N_99 ;
    wire \DUT.uart_inst0.un1_tx_bits_remaining_axb_3 ;
    wire P1A4_c;
    wire \DUT.fifo_rx_inst.rFifoDataro_3 ;
    wire \fifo_inst.ft2232h_inst.rFifoStateZ0Z_1 ;
    wire \fifo_inst.ft2232h_inst.N_103 ;
    wire \fifo_inst.ft2232h_inst.rFifoStateZ0Z_2 ;
    wire \DUT.fifo_rx_inst.rFifoDataro_2 ;
    wire \fifo_inst.ft2232h_inst.rFifoStateZ0Z_0 ;
    wire iTxE_n_c;
    wire iRxF_n_c;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_0 ;
    wire \DUT.fifo_rx_inst.rReadPtrZ0Z_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_7 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1 ;
    wire \DUT.fifo_rx_inst.rReadPtrZ0Z_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2 ;
    wire N_100_i_0;
    wire rFifoDatarff_0_RNIHJV05;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_2 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_4 ;
    wire \DUT.fifo_rx_inst.rFifoData_awe3 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_0 ;
    wire \DUT.wRxByte_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_1 ;
    wire \DUT.wRxByte_2 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_2 ;
    wire \DUT.wRxByte_3 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_3 ;
    wire \DUT.wRxByte_4 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_4 ;
    wire \DUT.wRxByte_5 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_5 ;
    wire \DUT.wRxByte_6 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_6 ;
    wire \DUT.wRxByte_7 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_7 ;
    wire \DUT.fifo_rx_inst.rFifoData_awe2 ;
    wire \DUT.wRxByte_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_awe0 ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddr_0_2 ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_1_1_cascade_ ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIZ0Z_1 ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddr_0_1 ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIZ0Z_1_cascade_ ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_1 ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_1_cascade_ ;
    wire \DUT.uart_inst0.tx_dataZ0Z_0 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_1 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_3 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_2 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_4 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_7 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_6 ;
    wire \DUT.tx_state_0 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_5 ;
    wire \DUT.uart_inst0.N_71_i ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_ ;
    wire \DUT.rFifoDatarx_4 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_4 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_ ;
    wire \DUT.rFifoDatarx_6 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_4 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_6 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_6 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_4 ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddr_0_7 ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddr_0_4 ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddr_0_6 ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_1_1 ;
    wire bfn_17_10_0_;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_2 ;
    wire \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1_c_RNI5GZ0Z02 ;
    wire \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1 ;
    wire \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2 ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_4 ;
    wire \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_3_c_RNI7KZ0Z22 ;
    wire \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_3 ;
    wire \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_4 ;
    wire \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_5_c_RNI9OZ0Z42 ;
    wire \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_5 ;
    wire \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_6_c_RNIAQZ0Z52 ;
    wire \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_6 ;
    wire \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_7 ;
    wire \fifo_inst.ft2232h_inst.rFifoState_RNIG8PKZ0Z_4 ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_7 ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_6 ;
    wire \fifo_inst.tx_fifo_inst.un15_rRamRdAddr_5 ;
    wire \fifo_inst.tx_fifo_inst.un15_rRamRdAddr_cascade_ ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddr_0_0 ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddr_rst_cascade_ ;
    wire bfn_17_12_0_;
    wire \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1 ;
    wire \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_3 ;
    wire \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIJ4MZ0Z4 ;
    wire \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2 ;
    wire \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3 ;
    wire \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_4 ;
    wire \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5 ;
    wire \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_7 ;
    wire \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6 ;
    wire \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_7 ;
    wire \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_8 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_3 ;
    wire \DUT.rFifoDatarx_3 ;
    wire \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_4 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_7 ;
    wire \DUT.rFifoDatarx_7 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_5 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_5 ;
    wire \DUT.rFifoDatarx_5 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1_cascade_ ;
    wire \DUT.rFifoDatarx_1 ;
    wire \DUT.fifo_tx_inst.rFifoDataro_0 ;
    wire \DUT.fifo_tx_inst.rFifoDataror_1_0_cascade_ ;
    wire \DUT.rFifoDataror_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_0 ;
    wire \DUT.rFifoDatarxZ0Z_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_5 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_3 ;
    wire rTxByteZ0Z_4;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_4 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_6 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_7 ;
    wire \DUT.fifo_tx_inst.rFifoDataro_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_awe2 ;
    wire \DUT.fifo_tx_inst.rFifoData_awe2_cascade_ ;
    wire \DUT.fifo_tx_inst.rFifoDataro_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_awe3_cascade_ ;
    wire \DUT.fifo_tx_inst.un1_i11_i ;
    wire \DUT.fifo_tx_inst.un1_i11_i_cascade_ ;
    wire \DUT.fifo_tx_inst.rWritePtrZ0Z_1 ;
    wire \DUT.fifo_tx_inst.rWritePtrZ0Z_0 ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddr_rst_7 ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddr_0_8 ;
    wire \fifo_inst.rTxRdEn_RNIS0VN ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddr_rst_4 ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddr_0_5 ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_5 ;
    wire \fifo_inst.tx_fifo_inst.un18_rRamWrAddr_4 ;
    wire \fifo_inst.tx_fifo_inst.un18_rRamWrAddr ;
    wire \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_2 ;
    wire \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI6IZ0Z12 ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddr_0_3 ;
    wire \fifo_inst.rTxRdEn_fast ;
    wire \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI20CZ0Z4_cascade_ ;
    wire \fifo_inst.tx_fifo_inst.un15_rRamRdAddr ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_3 ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_0 ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_3_cascade_ ;
    wire \fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_8 ;
    wire \fifo_inst.tx_fifo_inst.un15_rRamRdAddr_4 ;
    wire \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNII2LZ0Z4 ;
    wire \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_6 ;
    wire \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNIJQZ0Z47 ;
    wire \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_7 ;
    wire \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIK6NZ0Z4 ;
    wire \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_4 ;
    wire \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_5 ;
    wire \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_2 ;
    wire \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_4_cascade_ ;
    wire \fifo_inst.tx_fifo_inst.un18_rRamWrAddr_5 ;
    wire \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_1 ;
    wire \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_1_cascade_ ;
    wire \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_0 ;
    wire \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIZ0 ;
    wire \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIZ0_cascade_ ;
    wire \fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7 ;
    wire \DUT.fifo_tx_inst.N_101_cascade_ ;
    wire wPllLocked;
    wire \DUT.fifo_tx_inst.un1_i11_2_i_cascade_ ;
    wire wPllLocked_g;
    wire \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNIIOZ0Z37 ;
    wire \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_6 ;
    wire \DUT.fifo_tx_inst.N_101 ;
    wire \DUT.fifo_tx_inst.un1_i11_2_i ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_3 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_7 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0 ;
    wire rTxByteZ0Z_0;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_0 ;
    wire rTxByteZ0Z_1;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_1 ;
    wire \DUT.fifo_tx_inst.rReadPtrZ0Z_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_ ;
    wire \DUT.fifo_tx_inst.rReadPtrZ0Z_1 ;
    wire \DUT.rFifoDatarx_2 ;
    wire rTxByteZ0Z_2;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_2 ;
    wire rTxByteZ0Z_6;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_6 ;
    wire rTxByteZ0Z_7;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_7 ;
    wire rTxByteZ0Z_3;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_3 ;
    wire \DUT.fifo_tx_inst.N_105 ;
    wire \DUT.N_93_cascade_ ;
    wire \DUT.fifo_tx_inst.N_98_cascade_ ;
    wire \DUT.fifo_tx_inst.N_86 ;
    wire \DUT.N_93 ;
    wire \DUT.rTransmitZ0 ;
    wire rRxReadZ0;
    wire \DUT.fifo_tx_inst.N_98 ;
    wire \fifo_inst.ft2232h_inst.rFifoStateZ0Z_3 ;
    wire rTxByteZ0Z_5;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_5 ;
    wire \DUT.fifo_tx_inst.rFifoData_awe1 ;
    wire \fifo_inst.ft2232h_inst.rFifoStatec_0 ;
    wire \fifo_inst.ft2232h_inst.rFifoStateZ0Z_4 ;
    wire \fifo_inst.wTxRdEn ;
    wire rTxBusReady;
    wire \DUT.fifo_tx_inst.rFifoCountZ0Z_0 ;
    wire \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0 ;
    wire bfn_20_17_0_;
    wire \DUT.fifo_tx_inst.rFifoCount_RNIBPFMZ0Z_1 ;
    wire \DUT.fifo_tx_inst.rFifoCountZ0Z_1 ;
    wire \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0 ;
    wire \DUT.fifo_tx_inst.un1_rFifoCount_1_axb_2 ;
    wire \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1 ;
    wire \DUT.fifo_tx_inst.rFifoCountZ0Z_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_awe3 ;
    wire \DUT.fifo_tx_inst.rFifoDataro_3 ;
    wire _gnd_net_;
    wire clk_48mhz_0;
    wire wPllLocked_i_g;

    defparam \fifo_inst.tx_fifo_inst.ram512x8_inst_physical .WRITE_MODE=1;
    defparam \fifo_inst.tx_fifo_inst.ram512x8_inst_physical .READ_MODE=1;
    SB_RAM40_4K \fifo_inst.tx_fifo_inst.ram512x8_inst_physical  (
            .RDATA({dangling_wire_0,wTxRdData_7,dangling_wire_1,wTxRdData_6,dangling_wire_2,wTxRdData_5,dangling_wire_3,wTxRdData_4,dangling_wire_4,wTxRdData_3,dangling_wire_5,wTxRdData_2,dangling_wire_6,wTxRdData_1,dangling_wire_7,wTxRdData_0}),
            .RADDR({dangling_wire_8,dangling_wire_9,N__11445,N__10890,N__10857,N__11667,N__10728,N__11520,N__10773,N__10335,N__11499}),
            .WADDR({dangling_wire_10,dangling_wire_11,N__10965,N__11871,N__11403,N__11829,N__11841,N__8658,N__11799,N__11709,N__11760}),
            .MASK({dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27}),
            .WDATA({dangling_wire_28,dangling_wire_29,dangling_wire_30,N__8388,dangling_wire_31,dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,N__12167}),
            .RCLKE(),
            .RCLK(N__13500),
            .RE(N__13853),
            .WCLKE(),
            .WCLK(N__13499),
            .WE(N__12168));
    defparam \top_pll_inst.top_pll_inst_pll .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \top_pll_inst.top_pll_inst_pll .TEST_MODE=1'b0;
    defparam \top_pll_inst.top_pll_inst_pll .SHIFTREG_DIV_MODE=2'b00;
    defparam \top_pll_inst.top_pll_inst_pll .PLLOUT_SELECT="GENCLK";
    defparam \top_pll_inst.top_pll_inst_pll .FILTER_RANGE=3'b001;
    defparam \top_pll_inst.top_pll_inst_pll .FEEDBACK_PATH="SIMPLE";
    defparam \top_pll_inst.top_pll_inst_pll .FDA_RELATIVE=4'b0000;
    defparam \top_pll_inst.top_pll_inst_pll .FDA_FEEDBACK=4'b0000;
    defparam \top_pll_inst.top_pll_inst_pll .ENABLE_ICEGATE=1'b0;
    defparam \top_pll_inst.top_pll_inst_pll .DIVR=4'b0000;
    defparam \top_pll_inst.top_pll_inst_pll .DIVQ=3'b100;
    defparam \top_pll_inst.top_pll_inst_pll .DIVF=7'b0111111;
    defparam \top_pll_inst.top_pll_inst_pll .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    PLL40 \top_pll_inst.top_pll_inst_pll  (
            .PLLOUTGLOBAL(clk_48mhz_0),
            .SDI(GNDG0),
            .BYPASS(GNDG0),
            .RESETB(N__5433),
            .PLLOUTCORE(),
            .LOCK(\PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO ),
            .SDO(),
            .SCLK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .EXTFEEDBACK(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLIN(N__14220));
    IO_PAD \top_pll_inst.top_pll_inst_iopad  (
            .OE(VCCG0),
            .DIN(),
            .DOUT(N__14220),
            .PACKAGEPIN(iClk));
    IO_PAD P1A8_obuft_iopad (
            .OE(N__14206),
            .DIN(N__14205),
            .DOUT(N__14204),
            .PACKAGEPIN(P1A8));
    defparam P1A8_obuft_preio.NEG_TRIGGER=1'b0;
    defparam P1A8_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO P1A8_obuft_preio (
            .PADOEN(N__14206),
            .PADOUT(N__14205),
            .PADIN(N__14204),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_1_iopad (
            .OE(N__14197),
            .DIN(N__14196),
            .DOUT(N__14195),
            .PACKAGEPIN(ioFifoData[1]));
    defparam ioFifoData_obuft_1_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_1_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_1_preio (
            .PADOEN(N__14197),
            .PADOUT(N__14196),
            .PADIN(N__14195),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__13765),
            .DIN0(),
            .DOUT0(N__5502),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_4_iopad (
            .OE(N__14188),
            .DIN(N__14187),
            .DOUT(N__14186),
            .PACKAGEPIN(ioFifoData[4]));
    defparam ioFifoData_obuft_4_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_4_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_4_preio (
            .PADOEN(N__14188),
            .PADOUT(N__14187),
            .PADIN(N__14186),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__13749),
            .DIN0(),
            .DOUT0(N__5514),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A2_obuft_iopad (
            .OE(N__14179),
            .DIN(N__14178),
            .DOUT(N__14177),
            .PACKAGEPIN(P1A2));
    defparam P1A2_obuft_preio.NEG_TRIGGER=1'b0;
    defparam P1A2_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO P1A2_obuft_preio (
            .PADOEN(N__14179),
            .PADOUT(N__14178),
            .PADIN(N__14177),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A4_obuf_iopad (
            .OE(N__14170),
            .DIN(N__14169),
            .DOUT(N__14168),
            .PACKAGEPIN(P1A4));
    defparam P1A4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO P1A4_obuf_preio (
            .PADOEN(N__14170),
            .PADOUT(N__14169),
            .PADIN(N__14168),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9030),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_0_iopad (
            .OE(N__14161),
            .DIN(N__14160),
            .DOUT(N__14159),
            .PACKAGEPIN(ioFifoData[0]));
    defparam ioFifoData_obuft_0_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_0_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_0_preio (
            .PADOEN(N__14161),
            .PADOUT(N__14160),
            .PADIN(N__14159),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__13770),
            .DIN0(),
            .DOUT0(N__5454),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD oRx_n_obuf_iopad (
            .OE(N__14152),
            .DIN(N__14151),
            .DOUT(N__14150),
            .PACKAGEPIN(oRx_n));
    defparam oRx_n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam oRx_n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO oRx_n_obuf_preio (
            .PADOEN(N__14152),
            .PADOUT(N__14151),
            .PADIN(N__14150),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7667),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_7_iopad (
            .OE(N__14143),
            .DIN(N__14142),
            .DOUT(N__14141),
            .PACKAGEPIN(ioFifoData[7]));
    defparam ioFifoData_obuft_7_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_7_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_7_preio (
            .PADOEN(N__14143),
            .PADOUT(N__14142),
            .PADIN(N__14141),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__13763),
            .DIN0(),
            .DOUT0(N__5469),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD iRxF_n_ibuf_iopad (
            .OE(N__14134),
            .DIN(N__14133),
            .DOUT(N__14132),
            .PACKAGEPIN(iRxF_n));
    defparam iRxF_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam iRxF_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO iRxF_n_ibuf_preio (
            .PADOEN(N__14134),
            .PADOUT(N__14133),
            .PADIN(N__14132),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(iRxF_n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A3_obuf_iopad (
            .OE(N__14125),
            .DIN(N__14124),
            .DOUT(N__14123),
            .PACKAGEPIN(P1A3));
    defparam P1A3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO P1A3_obuf_preio (
            .PADOEN(N__14125),
            .PADOUT(N__14124),
            .PADIN(N__14123),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7674),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A7_obuf_iopad (
            .OE(N__14116),
            .DIN(N__14115),
            .DOUT(N__14114),
            .PACKAGEPIN(P1A7));
    defparam P1A7_obuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A7_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO P1A7_obuf_preio (
            .PADOEN(N__14116),
            .PADOUT(N__14115),
            .PADIN(N__14114),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8640),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BTN_N_ibuf_iopad (
            .OE(N__14107),
            .DIN(N__14106),
            .DOUT(N__14105),
            .PACKAGEPIN(BTN_N));
    defparam BTN_N_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam BTN_N_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO BTN_N_ibuf_preio (
            .PADOEN(N__14107),
            .PADOUT(N__14106),
            .PADIN(N__14105),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(BTN_N_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_3_iopad (
            .OE(N__14098),
            .DIN(N__14097),
            .DOUT(N__14096),
            .PACKAGEPIN(ioFifoData[3]));
    defparam ioFifoData_obuft_3_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_3_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_3_preio (
            .PADOEN(N__14098),
            .PADOUT(N__14097),
            .PADIN(N__14096),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__13729),
            .DIN0(),
            .DOUT0(N__5418),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_6_iopad (
            .OE(N__14089),
            .DIN(N__14088),
            .DOUT(N__14087),
            .PACKAGEPIN(ioFifoData[6]));
    defparam ioFifoData_obuft_6_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_6_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_6_preio (
            .PADOEN(N__14089),
            .PADOUT(N__14088),
            .PADIN(N__14087),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__13762),
            .DIN0(),
            .DOUT0(N__5370),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_5_iopad (
            .OE(N__14080),
            .DIN(N__14079),
            .DOUT(N__14078),
            .PACKAGEPIN(ioFifoData[5]));
    defparam ioFifoData_obuft_5_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_5_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_5_preio (
            .PADOEN(N__14080),
            .PADOUT(N__14079),
            .PADIN(N__14078),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__13764),
            .DIN0(),
            .DOUT0(N__5400),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD oTx_n_obuf_iopad (
            .OE(N__14071),
            .DIN(N__14070),
            .DOUT(N__14069),
            .PACKAGEPIN(oTx_n));
    defparam oTx_n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam oTx_n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO oTx_n_obuf_preio (
            .PADOEN(N__14071),
            .PADOUT(N__14070),
            .PADIN(N__14069),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9029),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD iTxE_n_ibuf_iopad (
            .OE(N__14062),
            .DIN(N__14061),
            .DOUT(N__14060),
            .PACKAGEPIN(iTxE_n));
    defparam iTxE_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam iTxE_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO iTxE_n_ibuf_preio (
            .PADOEN(N__14062),
            .PADOUT(N__14061),
            .PADIN(N__14060),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(iTxE_n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_2_iopad (
            .OE(N__14053),
            .DIN(N__14052),
            .DOUT(N__14051),
            .PACKAGEPIN(ioFifoData[2]));
    defparam ioFifoData_obuft_2_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_2_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_2_preio (
            .PADOEN(N__14053),
            .PADOUT(N__14052),
            .PADIN(N__14051),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__13769),
            .DIN0(),
            .DOUT0(N__5388),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A1_ibuf_iopad (
            .OE(N__14044),
            .DIN(N__14043),
            .DOUT(N__14042),
            .PACKAGEPIN(P1A1));
    defparam P1A1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO P1A1_ibuf_preio (
            .PADOEN(N__14044),
            .PADOUT(N__14043),
            .PADIN(N__14042),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(P1A1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A9_obuft_iopad (
            .OE(N__14035),
            .DIN(N__14034),
            .DOUT(N__14033),
            .PACKAGEPIN(P1A9));
    defparam P1A9_obuft_preio.NEG_TRIGGER=1'b0;
    defparam P1A9_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO P1A9_obuft_preio (
            .PADOEN(N__14035),
            .PADOUT(N__14034),
            .PADIN(N__14033),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__3332 (
            .O(N__14016),
            .I(N__14013));
    LocalMux I__3331 (
            .O(N__14013),
            .I(N__14009));
    InMux I__3330 (
            .O(N__14012),
            .I(N__14006));
    Span4Mux_v I__3329 (
            .O(N__14009),
            .I(N__14001));
    LocalMux I__3328 (
            .O(N__14006),
            .I(N__13998));
    InMux I__3327 (
            .O(N__14005),
            .I(N__13995));
    InMux I__3326 (
            .O(N__14004),
            .I(N__13992));
    Span4Mux_h I__3325 (
            .O(N__14001),
            .I(N__13987));
    Span4Mux_v I__3324 (
            .O(N__13998),
            .I(N__13987));
    LocalMux I__3323 (
            .O(N__13995),
            .I(N__13982));
    LocalMux I__3322 (
            .O(N__13992),
            .I(N__13982));
    Span4Mux_v I__3321 (
            .O(N__13987),
            .I(N__13979));
    Span4Mux_h I__3320 (
            .O(N__13982),
            .I(N__13976));
    Odrv4 I__3319 (
            .O(N__13979),
            .I(rTxByteZ0Z_5));
    Odrv4 I__3318 (
            .O(N__13976),
            .I(rTxByteZ0Z_5));
    InMux I__3317 (
            .O(N__13971),
            .I(N__13968));
    LocalMux I__3316 (
            .O(N__13968),
            .I(N__13965));
    Odrv4 I__3315 (
            .O(N__13965),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_5 ));
    CEMux I__3314 (
            .O(N__13962),
            .I(N__13958));
    CEMux I__3313 (
            .O(N__13961),
            .I(N__13955));
    LocalMux I__3312 (
            .O(N__13958),
            .I(N__13949));
    LocalMux I__3311 (
            .O(N__13955),
            .I(N__13949));
    CEMux I__3310 (
            .O(N__13954),
            .I(N__13946));
    Span4Mux_h I__3309 (
            .O(N__13949),
            .I(N__13942));
    LocalMux I__3308 (
            .O(N__13946),
            .I(N__13939));
    InMux I__3307 (
            .O(N__13945),
            .I(N__13936));
    Odrv4 I__3306 (
            .O(N__13942),
            .I(\DUT.fifo_tx_inst.rFifoData_awe1 ));
    Odrv4 I__3305 (
            .O(N__13939),
            .I(\DUT.fifo_tx_inst.rFifoData_awe1 ));
    LocalMux I__3304 (
            .O(N__13936),
            .I(\DUT.fifo_tx_inst.rFifoData_awe1 ));
    InMux I__3303 (
            .O(N__13929),
            .I(N__13926));
    LocalMux I__3302 (
            .O(N__13926),
            .I(N__13923));
    Odrv12 I__3301 (
            .O(N__13923),
            .I(\fifo_inst.ft2232h_inst.rFifoStatec_0 ));
    InMux I__3300 (
            .O(N__13920),
            .I(N__13914));
    InMux I__3299 (
            .O(N__13919),
            .I(N__13914));
    LocalMux I__3298 (
            .O(N__13914),
            .I(N__13908));
    InMux I__3297 (
            .O(N__13913),
            .I(N__13904));
    InMux I__3296 (
            .O(N__13912),
            .I(N__13899));
    InMux I__3295 (
            .O(N__13911),
            .I(N__13899));
    Span4Mux_v I__3294 (
            .O(N__13908),
            .I(N__13895));
    InMux I__3293 (
            .O(N__13907),
            .I(N__13892));
    LocalMux I__3292 (
            .O(N__13904),
            .I(N__13887));
    LocalMux I__3291 (
            .O(N__13899),
            .I(N__13887));
    InMux I__3290 (
            .O(N__13898),
            .I(N__13884));
    Span4Mux_h I__3289 (
            .O(N__13895),
            .I(N__13877));
    LocalMux I__3288 (
            .O(N__13892),
            .I(N__13877));
    Span4Mux_h I__3287 (
            .O(N__13887),
            .I(N__13877));
    LocalMux I__3286 (
            .O(N__13884),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_4 ));
    Odrv4 I__3285 (
            .O(N__13877),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_4 ));
    CascadeMux I__3284 (
            .O(N__13872),
            .I(N__13867));
    CascadeMux I__3283 (
            .O(N__13871),
            .I(N__13864));
    CascadeMux I__3282 (
            .O(N__13870),
            .I(N__13860));
    InMux I__3281 (
            .O(N__13867),
            .I(N__13855));
    InMux I__3280 (
            .O(N__13864),
            .I(N__13855));
    InMux I__3279 (
            .O(N__13863),
            .I(N__13850));
    InMux I__3278 (
            .O(N__13860),
            .I(N__13847));
    LocalMux I__3277 (
            .O(N__13855),
            .I(N__13844));
    InMux I__3276 (
            .O(N__13854),
            .I(N__13840));
    SRMux I__3275 (
            .O(N__13853),
            .I(N__13835));
    LocalMux I__3274 (
            .O(N__13850),
            .I(N__13830));
    LocalMux I__3273 (
            .O(N__13847),
            .I(N__13830));
    Span4Mux_h I__3272 (
            .O(N__13844),
            .I(N__13823));
    InMux I__3271 (
            .O(N__13843),
            .I(N__13820));
    LocalMux I__3270 (
            .O(N__13840),
            .I(N__13817));
    CascadeMux I__3269 (
            .O(N__13839),
            .I(N__13814));
    CascadeMux I__3268 (
            .O(N__13838),
            .I(N__13811));
    LocalMux I__3267 (
            .O(N__13835),
            .I(N__13808));
    Span4Mux_v I__3266 (
            .O(N__13830),
            .I(N__13805));
    InMux I__3265 (
            .O(N__13829),
            .I(N__13796));
    InMux I__3264 (
            .O(N__13828),
            .I(N__13796));
    InMux I__3263 (
            .O(N__13827),
            .I(N__13796));
    InMux I__3262 (
            .O(N__13826),
            .I(N__13796));
    Span4Mux_v I__3261 (
            .O(N__13823),
            .I(N__13791));
    LocalMux I__3260 (
            .O(N__13820),
            .I(N__13791));
    Span4Mux_h I__3259 (
            .O(N__13817),
            .I(N__13788));
    InMux I__3258 (
            .O(N__13814),
            .I(N__13783));
    InMux I__3257 (
            .O(N__13811),
            .I(N__13783));
    Odrv4 I__3256 (
            .O(N__13808),
            .I(\fifo_inst.wTxRdEn ));
    Odrv4 I__3255 (
            .O(N__13805),
            .I(\fifo_inst.wTxRdEn ));
    LocalMux I__3254 (
            .O(N__13796),
            .I(\fifo_inst.wTxRdEn ));
    Odrv4 I__3253 (
            .O(N__13791),
            .I(\fifo_inst.wTxRdEn ));
    Odrv4 I__3252 (
            .O(N__13788),
            .I(\fifo_inst.wTxRdEn ));
    LocalMux I__3251 (
            .O(N__13783),
            .I(\fifo_inst.wTxRdEn ));
    IoInMux I__3250 (
            .O(N__13770),
            .I(N__13766));
    IoInMux I__3249 (
            .O(N__13769),
            .I(N__13759));
    LocalMux I__3248 (
            .O(N__13766),
            .I(N__13756));
    IoInMux I__3247 (
            .O(N__13765),
            .I(N__13753));
    IoInMux I__3246 (
            .O(N__13764),
            .I(N__13750));
    IoInMux I__3245 (
            .O(N__13763),
            .I(N__13746));
    IoInMux I__3244 (
            .O(N__13762),
            .I(N__13743));
    LocalMux I__3243 (
            .O(N__13759),
            .I(N__13740));
    IoSpan4Mux I__3242 (
            .O(N__13756),
            .I(N__13733));
    LocalMux I__3241 (
            .O(N__13753),
            .I(N__13733));
    LocalMux I__3240 (
            .O(N__13750),
            .I(N__13733));
    IoInMux I__3239 (
            .O(N__13749),
            .I(N__13730));
    LocalMux I__3238 (
            .O(N__13746),
            .I(N__13724));
    LocalMux I__3237 (
            .O(N__13743),
            .I(N__13724));
    IoSpan4Mux I__3236 (
            .O(N__13740),
            .I(N__13719));
    IoSpan4Mux I__3235 (
            .O(N__13733),
            .I(N__13719));
    LocalMux I__3234 (
            .O(N__13730),
            .I(N__13716));
    IoInMux I__3233 (
            .O(N__13729),
            .I(N__13713));
    Span4Mux_s3_v I__3232 (
            .O(N__13724),
            .I(N__13710));
    Span4Mux_s2_v I__3231 (
            .O(N__13719),
            .I(N__13705));
    Span4Mux_s2_v I__3230 (
            .O(N__13716),
            .I(N__13705));
    LocalMux I__3229 (
            .O(N__13713),
            .I(N__13702));
    Span4Mux_v I__3228 (
            .O(N__13710),
            .I(N__13699));
    Span4Mux_v I__3227 (
            .O(N__13705),
            .I(N__13696));
    Span12Mux_s2_v I__3226 (
            .O(N__13702),
            .I(N__13693));
    Span4Mux_v I__3225 (
            .O(N__13699),
            .I(N__13690));
    Span4Mux_v I__3224 (
            .O(N__13696),
            .I(N__13687));
    Span12Mux_v I__3223 (
            .O(N__13693),
            .I(N__13683));
    Span4Mux_v I__3222 (
            .O(N__13690),
            .I(N__13678));
    Span4Mux_v I__3221 (
            .O(N__13687),
            .I(N__13678));
    InMux I__3220 (
            .O(N__13686),
            .I(N__13675));
    Odrv12 I__3219 (
            .O(N__13683),
            .I(rTxBusReady));
    Odrv4 I__3218 (
            .O(N__13678),
            .I(rTxBusReady));
    LocalMux I__3217 (
            .O(N__13675),
            .I(rTxBusReady));
    InMux I__3216 (
            .O(N__13668),
            .I(N__13664));
    CascadeMux I__3215 (
            .O(N__13667),
            .I(N__13661));
    LocalMux I__3214 (
            .O(N__13664),
            .I(N__13658));
    InMux I__3213 (
            .O(N__13661),
            .I(N__13653));
    Span4Mux_h I__3212 (
            .O(N__13658),
            .I(N__13650));
    InMux I__3211 (
            .O(N__13657),
            .I(N__13645));
    InMux I__3210 (
            .O(N__13656),
            .I(N__13645));
    LocalMux I__3209 (
            .O(N__13653),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_0 ));
    Odrv4 I__3208 (
            .O(N__13650),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_0 ));
    LocalMux I__3207 (
            .O(N__13645),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_0 ));
    CascadeMux I__3206 (
            .O(N__13638),
            .I(N__13635));
    InMux I__3205 (
            .O(N__13635),
            .I(N__13632));
    LocalMux I__3204 (
            .O(N__13632),
            .I(N__13629));
    Odrv4 I__3203 (
            .O(N__13629),
            .I(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0 ));
    CascadeMux I__3202 (
            .O(N__13626),
            .I(N__13623));
    InMux I__3201 (
            .O(N__13623),
            .I(N__13620));
    LocalMux I__3200 (
            .O(N__13620),
            .I(N__13617));
    Odrv4 I__3199 (
            .O(N__13617),
            .I(\DUT.fifo_tx_inst.rFifoCount_RNIBPFMZ0Z_1 ));
    CascadeMux I__3198 (
            .O(N__13614),
            .I(N__13611));
    InMux I__3197 (
            .O(N__13611),
            .I(N__13604));
    InMux I__3196 (
            .O(N__13610),
            .I(N__13604));
    InMux I__3195 (
            .O(N__13609),
            .I(N__13601));
    LocalMux I__3194 (
            .O(N__13604),
            .I(N__13598));
    LocalMux I__3193 (
            .O(N__13601),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_1 ));
    Odrv4 I__3192 (
            .O(N__13598),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_1 ));
    InMux I__3191 (
            .O(N__13593),
            .I(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0 ));
    InMux I__3190 (
            .O(N__13590),
            .I(N__13587));
    LocalMux I__3189 (
            .O(N__13587),
            .I(N__13584));
    Odrv12 I__3188 (
            .O(N__13584),
            .I(\DUT.fifo_tx_inst.un1_rFifoCount_1_axb_2 ));
    InMux I__3187 (
            .O(N__13581),
            .I(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1 ));
    InMux I__3186 (
            .O(N__13578),
            .I(N__13574));
    CascadeMux I__3185 (
            .O(N__13577),
            .I(N__13570));
    LocalMux I__3184 (
            .O(N__13574),
            .I(N__13564));
    InMux I__3183 (
            .O(N__13573),
            .I(N__13561));
    InMux I__3182 (
            .O(N__13570),
            .I(N__13552));
    InMux I__3181 (
            .O(N__13569),
            .I(N__13552));
    InMux I__3180 (
            .O(N__13568),
            .I(N__13552));
    InMux I__3179 (
            .O(N__13567),
            .I(N__13552));
    Span4Mux_h I__3178 (
            .O(N__13564),
            .I(N__13549));
    LocalMux I__3177 (
            .O(N__13561),
            .I(N__13544));
    LocalMux I__3176 (
            .O(N__13552),
            .I(N__13544));
    Odrv4 I__3175 (
            .O(N__13549),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_2 ));
    Odrv4 I__3174 (
            .O(N__13544),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_2 ));
    InMux I__3173 (
            .O(N__13539),
            .I(N__13535));
    CEMux I__3172 (
            .O(N__13538),
            .I(N__13532));
    LocalMux I__3171 (
            .O(N__13535),
            .I(N__13529));
    LocalMux I__3170 (
            .O(N__13532),
            .I(N__13526));
    Span4Mux_h I__3169 (
            .O(N__13529),
            .I(N__13523));
    Odrv4 I__3168 (
            .O(N__13526),
            .I(\DUT.fifo_tx_inst.rFifoData_awe3 ));
    Odrv4 I__3167 (
            .O(N__13523),
            .I(\DUT.fifo_tx_inst.rFifoData_awe3 ));
    InMux I__3166 (
            .O(N__13518),
            .I(N__13515));
    LocalMux I__3165 (
            .O(N__13515),
            .I(N__13511));
    InMux I__3164 (
            .O(N__13514),
            .I(N__13508));
    Span4Mux_h I__3163 (
            .O(N__13511),
            .I(N__13505));
    LocalMux I__3162 (
            .O(N__13508),
            .I(\DUT.fifo_tx_inst.rFifoDataro_3 ));
    Odrv4 I__3161 (
            .O(N__13505),
            .I(\DUT.fifo_tx_inst.rFifoDataro_3 ));
    ClkMux I__3160 (
            .O(N__13500),
            .I(N__13296));
    ClkMux I__3159 (
            .O(N__13499),
            .I(N__13296));
    ClkMux I__3158 (
            .O(N__13498),
            .I(N__13296));
    ClkMux I__3157 (
            .O(N__13497),
            .I(N__13296));
    ClkMux I__3156 (
            .O(N__13496),
            .I(N__13296));
    ClkMux I__3155 (
            .O(N__13495),
            .I(N__13296));
    ClkMux I__3154 (
            .O(N__13494),
            .I(N__13296));
    ClkMux I__3153 (
            .O(N__13493),
            .I(N__13296));
    ClkMux I__3152 (
            .O(N__13492),
            .I(N__13296));
    ClkMux I__3151 (
            .O(N__13491),
            .I(N__13296));
    ClkMux I__3150 (
            .O(N__13490),
            .I(N__13296));
    ClkMux I__3149 (
            .O(N__13489),
            .I(N__13296));
    ClkMux I__3148 (
            .O(N__13488),
            .I(N__13296));
    ClkMux I__3147 (
            .O(N__13487),
            .I(N__13296));
    ClkMux I__3146 (
            .O(N__13486),
            .I(N__13296));
    ClkMux I__3145 (
            .O(N__13485),
            .I(N__13296));
    ClkMux I__3144 (
            .O(N__13484),
            .I(N__13296));
    ClkMux I__3143 (
            .O(N__13483),
            .I(N__13296));
    ClkMux I__3142 (
            .O(N__13482),
            .I(N__13296));
    ClkMux I__3141 (
            .O(N__13481),
            .I(N__13296));
    ClkMux I__3140 (
            .O(N__13480),
            .I(N__13296));
    ClkMux I__3139 (
            .O(N__13479),
            .I(N__13296));
    ClkMux I__3138 (
            .O(N__13478),
            .I(N__13296));
    ClkMux I__3137 (
            .O(N__13477),
            .I(N__13296));
    ClkMux I__3136 (
            .O(N__13476),
            .I(N__13296));
    ClkMux I__3135 (
            .O(N__13475),
            .I(N__13296));
    ClkMux I__3134 (
            .O(N__13474),
            .I(N__13296));
    ClkMux I__3133 (
            .O(N__13473),
            .I(N__13296));
    ClkMux I__3132 (
            .O(N__13472),
            .I(N__13296));
    ClkMux I__3131 (
            .O(N__13471),
            .I(N__13296));
    ClkMux I__3130 (
            .O(N__13470),
            .I(N__13296));
    ClkMux I__3129 (
            .O(N__13469),
            .I(N__13296));
    ClkMux I__3128 (
            .O(N__13468),
            .I(N__13296));
    ClkMux I__3127 (
            .O(N__13467),
            .I(N__13296));
    ClkMux I__3126 (
            .O(N__13466),
            .I(N__13296));
    ClkMux I__3125 (
            .O(N__13465),
            .I(N__13296));
    ClkMux I__3124 (
            .O(N__13464),
            .I(N__13296));
    ClkMux I__3123 (
            .O(N__13463),
            .I(N__13296));
    ClkMux I__3122 (
            .O(N__13462),
            .I(N__13296));
    ClkMux I__3121 (
            .O(N__13461),
            .I(N__13296));
    ClkMux I__3120 (
            .O(N__13460),
            .I(N__13296));
    ClkMux I__3119 (
            .O(N__13459),
            .I(N__13296));
    ClkMux I__3118 (
            .O(N__13458),
            .I(N__13296));
    ClkMux I__3117 (
            .O(N__13457),
            .I(N__13296));
    ClkMux I__3116 (
            .O(N__13456),
            .I(N__13296));
    ClkMux I__3115 (
            .O(N__13455),
            .I(N__13296));
    ClkMux I__3114 (
            .O(N__13454),
            .I(N__13296));
    ClkMux I__3113 (
            .O(N__13453),
            .I(N__13296));
    ClkMux I__3112 (
            .O(N__13452),
            .I(N__13296));
    ClkMux I__3111 (
            .O(N__13451),
            .I(N__13296));
    ClkMux I__3110 (
            .O(N__13450),
            .I(N__13296));
    ClkMux I__3109 (
            .O(N__13449),
            .I(N__13296));
    ClkMux I__3108 (
            .O(N__13448),
            .I(N__13296));
    ClkMux I__3107 (
            .O(N__13447),
            .I(N__13296));
    ClkMux I__3106 (
            .O(N__13446),
            .I(N__13296));
    ClkMux I__3105 (
            .O(N__13445),
            .I(N__13296));
    ClkMux I__3104 (
            .O(N__13444),
            .I(N__13296));
    ClkMux I__3103 (
            .O(N__13443),
            .I(N__13296));
    ClkMux I__3102 (
            .O(N__13442),
            .I(N__13296));
    ClkMux I__3101 (
            .O(N__13441),
            .I(N__13296));
    ClkMux I__3100 (
            .O(N__13440),
            .I(N__13296));
    ClkMux I__3099 (
            .O(N__13439),
            .I(N__13296));
    ClkMux I__3098 (
            .O(N__13438),
            .I(N__13296));
    ClkMux I__3097 (
            .O(N__13437),
            .I(N__13296));
    ClkMux I__3096 (
            .O(N__13436),
            .I(N__13296));
    ClkMux I__3095 (
            .O(N__13435),
            .I(N__13296));
    ClkMux I__3094 (
            .O(N__13434),
            .I(N__13296));
    ClkMux I__3093 (
            .O(N__13433),
            .I(N__13296));
    GlobalMux I__3092 (
            .O(N__13296),
            .I(clk_48mhz_0));
    SRMux I__3091 (
            .O(N__13293),
            .I(N__13245));
    SRMux I__3090 (
            .O(N__13292),
            .I(N__13245));
    SRMux I__3089 (
            .O(N__13291),
            .I(N__13245));
    SRMux I__3088 (
            .O(N__13290),
            .I(N__13245));
    SRMux I__3087 (
            .O(N__13289),
            .I(N__13245));
    SRMux I__3086 (
            .O(N__13288),
            .I(N__13245));
    SRMux I__3085 (
            .O(N__13287),
            .I(N__13245));
    SRMux I__3084 (
            .O(N__13286),
            .I(N__13245));
    SRMux I__3083 (
            .O(N__13285),
            .I(N__13245));
    SRMux I__3082 (
            .O(N__13284),
            .I(N__13245));
    SRMux I__3081 (
            .O(N__13283),
            .I(N__13245));
    SRMux I__3080 (
            .O(N__13282),
            .I(N__13245));
    SRMux I__3079 (
            .O(N__13281),
            .I(N__13245));
    SRMux I__3078 (
            .O(N__13280),
            .I(N__13245));
    SRMux I__3077 (
            .O(N__13279),
            .I(N__13245));
    SRMux I__3076 (
            .O(N__13278),
            .I(N__13245));
    GlobalMux I__3075 (
            .O(N__13245),
            .I(N__13242));
    gio2CtrlBuf I__3074 (
            .O(N__13242),
            .I(wPllLocked_i_g));
    InMux I__3073 (
            .O(N__13239),
            .I(N__13235));
    InMux I__3072 (
            .O(N__13238),
            .I(N__13232));
    LocalMux I__3071 (
            .O(N__13235),
            .I(N__13228));
    LocalMux I__3070 (
            .O(N__13232),
            .I(N__13225));
    InMux I__3069 (
            .O(N__13231),
            .I(N__13222));
    Span4Mux_v I__3068 (
            .O(N__13228),
            .I(N__13214));
    Span4Mux_v I__3067 (
            .O(N__13225),
            .I(N__13214));
    LocalMux I__3066 (
            .O(N__13222),
            .I(N__13214));
    InMux I__3065 (
            .O(N__13221),
            .I(N__13211));
    Span4Mux_h I__3064 (
            .O(N__13214),
            .I(N__13208));
    LocalMux I__3063 (
            .O(N__13211),
            .I(N__13205));
    Span4Mux_v I__3062 (
            .O(N__13208),
            .I(N__13202));
    Span4Mux_v I__3061 (
            .O(N__13205),
            .I(N__13199));
    Odrv4 I__3060 (
            .O(N__13202),
            .I(rTxByteZ0Z_3));
    Odrv4 I__3059 (
            .O(N__13199),
            .I(rTxByteZ0Z_3));
    InMux I__3058 (
            .O(N__13194),
            .I(N__13191));
    LocalMux I__3057 (
            .O(N__13191),
            .I(N__13188));
    Odrv4 I__3056 (
            .O(N__13188),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_3 ));
    CEMux I__3055 (
            .O(N__13185),
            .I(N__13182));
    LocalMux I__3054 (
            .O(N__13182),
            .I(N__13178));
    CEMux I__3053 (
            .O(N__13181),
            .I(N__13175));
    Span4Mux_h I__3052 (
            .O(N__13178),
            .I(N__13168));
    LocalMux I__3051 (
            .O(N__13175),
            .I(N__13168));
    CEMux I__3050 (
            .O(N__13174),
            .I(N__13165));
    InMux I__3049 (
            .O(N__13173),
            .I(N__13162));
    Span4Mux_h I__3048 (
            .O(N__13168),
            .I(N__13159));
    LocalMux I__3047 (
            .O(N__13165),
            .I(N__13156));
    LocalMux I__3046 (
            .O(N__13162),
            .I(N__13153));
    Odrv4 I__3045 (
            .O(N__13159),
            .I(\DUT.fifo_tx_inst.N_105 ));
    Odrv12 I__3044 (
            .O(N__13156),
            .I(\DUT.fifo_tx_inst.N_105 ));
    Odrv4 I__3043 (
            .O(N__13153),
            .I(\DUT.fifo_tx_inst.N_105 ));
    CascadeMux I__3042 (
            .O(N__13146),
            .I(\DUT.N_93_cascade_ ));
    CascadeMux I__3041 (
            .O(N__13143),
            .I(\DUT.fifo_tx_inst.N_98_cascade_ ));
    InMux I__3040 (
            .O(N__13140),
            .I(N__13131));
    InMux I__3039 (
            .O(N__13139),
            .I(N__13131));
    InMux I__3038 (
            .O(N__13138),
            .I(N__13124));
    InMux I__3037 (
            .O(N__13137),
            .I(N__13124));
    InMux I__3036 (
            .O(N__13136),
            .I(N__13124));
    LocalMux I__3035 (
            .O(N__13131),
            .I(\DUT.fifo_tx_inst.N_86 ));
    LocalMux I__3034 (
            .O(N__13124),
            .I(\DUT.fifo_tx_inst.N_86 ));
    InMux I__3033 (
            .O(N__13119),
            .I(N__13116));
    LocalMux I__3032 (
            .O(N__13116),
            .I(N__13111));
    InMux I__3031 (
            .O(N__13115),
            .I(N__13104));
    InMux I__3030 (
            .O(N__13114),
            .I(N__13104));
    Span12Mux_v I__3029 (
            .O(N__13111),
            .I(N__13101));
    InMux I__3028 (
            .O(N__13110),
            .I(N__13098));
    InMux I__3027 (
            .O(N__13109),
            .I(N__13095));
    LocalMux I__3026 (
            .O(N__13104),
            .I(N__13092));
    Odrv12 I__3025 (
            .O(N__13101),
            .I(\DUT.N_93 ));
    LocalMux I__3024 (
            .O(N__13098),
            .I(\DUT.N_93 ));
    LocalMux I__3023 (
            .O(N__13095),
            .I(\DUT.N_93 ));
    Odrv12 I__3022 (
            .O(N__13092),
            .I(\DUT.N_93 ));
    InMux I__3021 (
            .O(N__13083),
            .I(N__13073));
    InMux I__3020 (
            .O(N__13082),
            .I(N__13073));
    InMux I__3019 (
            .O(N__13081),
            .I(N__13066));
    InMux I__3018 (
            .O(N__13080),
            .I(N__13066));
    InMux I__3017 (
            .O(N__13079),
            .I(N__13066));
    CascadeMux I__3016 (
            .O(N__13078),
            .I(N__13062));
    LocalMux I__3015 (
            .O(N__13073),
            .I(N__13059));
    LocalMux I__3014 (
            .O(N__13066),
            .I(N__13056));
    CascadeMux I__3013 (
            .O(N__13065),
            .I(N__13053));
    InMux I__3012 (
            .O(N__13062),
            .I(N__13049));
    Span4Mux_v I__3011 (
            .O(N__13059),
            .I(N__13044));
    Span4Mux_v I__3010 (
            .O(N__13056),
            .I(N__13044));
    InMux I__3009 (
            .O(N__13053),
            .I(N__13041));
    InMux I__3008 (
            .O(N__13052),
            .I(N__13038));
    LocalMux I__3007 (
            .O(N__13049),
            .I(N__13029));
    Span4Mux_h I__3006 (
            .O(N__13044),
            .I(N__13029));
    LocalMux I__3005 (
            .O(N__13041),
            .I(N__13029));
    LocalMux I__3004 (
            .O(N__13038),
            .I(N__13029));
    Odrv4 I__3003 (
            .O(N__13029),
            .I(\DUT.rTransmitZ0 ));
    InMux I__3002 (
            .O(N__13026),
            .I(N__13023));
    LocalMux I__3001 (
            .O(N__13023),
            .I(N__13012));
    InMux I__3000 (
            .O(N__13022),
            .I(N__13009));
    InMux I__2999 (
            .O(N__13021),
            .I(N__13000));
    InMux I__2998 (
            .O(N__13020),
            .I(N__13000));
    InMux I__2997 (
            .O(N__13019),
            .I(N__13000));
    InMux I__2996 (
            .O(N__13018),
            .I(N__13000));
    InMux I__2995 (
            .O(N__13017),
            .I(N__12997));
    InMux I__2994 (
            .O(N__13016),
            .I(N__12992));
    InMux I__2993 (
            .O(N__13015),
            .I(N__12992));
    Span4Mux_v I__2992 (
            .O(N__13012),
            .I(N__12983));
    LocalMux I__2991 (
            .O(N__13009),
            .I(N__12983));
    LocalMux I__2990 (
            .O(N__13000),
            .I(N__12983));
    LocalMux I__2989 (
            .O(N__12997),
            .I(N__12983));
    LocalMux I__2988 (
            .O(N__12992),
            .I(N__12980));
    Span4Mux_h I__2987 (
            .O(N__12983),
            .I(N__12977));
    Odrv12 I__2986 (
            .O(N__12980),
            .I(rRxReadZ0));
    Odrv4 I__2985 (
            .O(N__12977),
            .I(rRxReadZ0));
    InMux I__2984 (
            .O(N__12972),
            .I(N__12969));
    LocalMux I__2983 (
            .O(N__12969),
            .I(\DUT.fifo_tx_inst.N_98 ));
    InMux I__2982 (
            .O(N__12966),
            .I(N__12963));
    LocalMux I__2981 (
            .O(N__12963),
            .I(N__12960));
    Span4Mux_h I__2980 (
            .O(N__12960),
            .I(N__12956));
    InMux I__2979 (
            .O(N__12959),
            .I(N__12953));
    Span4Mux_h I__2978 (
            .O(N__12956),
            .I(N__12950));
    LocalMux I__2977 (
            .O(N__12953),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_3 ));
    Odrv4 I__2976 (
            .O(N__12950),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_3 ));
    InMux I__2975 (
            .O(N__12945),
            .I(N__12942));
    LocalMux I__2974 (
            .O(N__12942),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_0 ));
    InMux I__2973 (
            .O(N__12939),
            .I(N__12936));
    LocalMux I__2972 (
            .O(N__12936),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0 ));
    InMux I__2971 (
            .O(N__12933),
            .I(N__12930));
    LocalMux I__2970 (
            .O(N__12930),
            .I(N__12925));
    InMux I__2969 (
            .O(N__12929),
            .I(N__12922));
    InMux I__2968 (
            .O(N__12928),
            .I(N__12919));
    Span4Mux_v I__2967 (
            .O(N__12925),
            .I(N__12911));
    LocalMux I__2966 (
            .O(N__12922),
            .I(N__12911));
    LocalMux I__2965 (
            .O(N__12919),
            .I(N__12911));
    InMux I__2964 (
            .O(N__12918),
            .I(N__12908));
    Span4Mux_h I__2963 (
            .O(N__12911),
            .I(N__12905));
    LocalMux I__2962 (
            .O(N__12908),
            .I(N__12902));
    Odrv4 I__2961 (
            .O(N__12905),
            .I(rTxByteZ0Z_0));
    Odrv4 I__2960 (
            .O(N__12902),
            .I(rTxByteZ0Z_0));
    InMux I__2959 (
            .O(N__12897),
            .I(N__12894));
    LocalMux I__2958 (
            .O(N__12894),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_0 ));
    InMux I__2957 (
            .O(N__12891),
            .I(N__12888));
    LocalMux I__2956 (
            .O(N__12888),
            .I(N__12883));
    InMux I__2955 (
            .O(N__12887),
            .I(N__12880));
    InMux I__2954 (
            .O(N__12886),
            .I(N__12877));
    Span4Mux_v I__2953 (
            .O(N__12883),
            .I(N__12869));
    LocalMux I__2952 (
            .O(N__12880),
            .I(N__12869));
    LocalMux I__2951 (
            .O(N__12877),
            .I(N__12869));
    InMux I__2950 (
            .O(N__12876),
            .I(N__12866));
    Span4Mux_h I__2949 (
            .O(N__12869),
            .I(N__12863));
    LocalMux I__2948 (
            .O(N__12866),
            .I(N__12860));
    Odrv4 I__2947 (
            .O(N__12863),
            .I(rTxByteZ0Z_1));
    Odrv4 I__2946 (
            .O(N__12860),
            .I(rTxByteZ0Z_1));
    InMux I__2945 (
            .O(N__12855),
            .I(N__12852));
    LocalMux I__2944 (
            .O(N__12852),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_1 ));
    InMux I__2943 (
            .O(N__12849),
            .I(N__12840));
    InMux I__2942 (
            .O(N__12848),
            .I(N__12840));
    InMux I__2941 (
            .O(N__12847),
            .I(N__12829));
    InMux I__2940 (
            .O(N__12846),
            .I(N__12829));
    InMux I__2939 (
            .O(N__12845),
            .I(N__12826));
    LocalMux I__2938 (
            .O(N__12840),
            .I(N__12823));
    InMux I__2937 (
            .O(N__12839),
            .I(N__12820));
    InMux I__2936 (
            .O(N__12838),
            .I(N__12817));
    InMux I__2935 (
            .O(N__12837),
            .I(N__12810));
    InMux I__2934 (
            .O(N__12836),
            .I(N__12810));
    InMux I__2933 (
            .O(N__12835),
            .I(N__12810));
    InMux I__2932 (
            .O(N__12834),
            .I(N__12807));
    LocalMux I__2931 (
            .O(N__12829),
            .I(N__12800));
    LocalMux I__2930 (
            .O(N__12826),
            .I(N__12800));
    Span4Mux_v I__2929 (
            .O(N__12823),
            .I(N__12800));
    LocalMux I__2928 (
            .O(N__12820),
            .I(N__12795));
    LocalMux I__2927 (
            .O(N__12817),
            .I(N__12795));
    LocalMux I__2926 (
            .O(N__12810),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__2925 (
            .O(N__12807),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    Odrv4 I__2924 (
            .O(N__12800),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    Odrv4 I__2923 (
            .O(N__12795),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    InMux I__2922 (
            .O(N__12786),
            .I(N__12783));
    LocalMux I__2921 (
            .O(N__12783),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_2 ));
    InMux I__2920 (
            .O(N__12780),
            .I(N__12777));
    LocalMux I__2919 (
            .O(N__12777),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_2 ));
    InMux I__2918 (
            .O(N__12774),
            .I(N__12771));
    LocalMux I__2917 (
            .O(N__12771),
            .I(N__12768));
    Span4Mux_h I__2916 (
            .O(N__12768),
            .I(N__12765));
    Odrv4 I__2915 (
            .O(N__12765),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_2 ));
    CascadeMux I__2914 (
            .O(N__12762),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_ ));
    CascadeMux I__2913 (
            .O(N__12759),
            .I(N__12753));
    CascadeMux I__2912 (
            .O(N__12758),
            .I(N__12750));
    InMux I__2911 (
            .O(N__12757),
            .I(N__12736));
    InMux I__2910 (
            .O(N__12756),
            .I(N__12736));
    InMux I__2909 (
            .O(N__12753),
            .I(N__12736));
    InMux I__2908 (
            .O(N__12750),
            .I(N__12736));
    CascadeMux I__2907 (
            .O(N__12749),
            .I(N__12731));
    CascadeMux I__2906 (
            .O(N__12748),
            .I(N__12727));
    CascadeMux I__2905 (
            .O(N__12747),
            .I(N__12717));
    CascadeMux I__2904 (
            .O(N__12746),
            .I(N__12714));
    CascadeMux I__2903 (
            .O(N__12745),
            .I(N__12710));
    LocalMux I__2902 (
            .O(N__12736),
            .I(N__12707));
    InMux I__2901 (
            .O(N__12735),
            .I(N__12700));
    InMux I__2900 (
            .O(N__12734),
            .I(N__12700));
    InMux I__2899 (
            .O(N__12731),
            .I(N__12700));
    InMux I__2898 (
            .O(N__12730),
            .I(N__12697));
    InMux I__2897 (
            .O(N__12727),
            .I(N__12694));
    InMux I__2896 (
            .O(N__12726),
            .I(N__12687));
    InMux I__2895 (
            .O(N__12725),
            .I(N__12687));
    InMux I__2894 (
            .O(N__12724),
            .I(N__12687));
    InMux I__2893 (
            .O(N__12723),
            .I(N__12674));
    InMux I__2892 (
            .O(N__12722),
            .I(N__12674));
    InMux I__2891 (
            .O(N__12721),
            .I(N__12674));
    InMux I__2890 (
            .O(N__12720),
            .I(N__12674));
    InMux I__2889 (
            .O(N__12717),
            .I(N__12674));
    InMux I__2888 (
            .O(N__12714),
            .I(N__12674));
    InMux I__2887 (
            .O(N__12713),
            .I(N__12669));
    InMux I__2886 (
            .O(N__12710),
            .I(N__12669));
    Span4Mux_h I__2885 (
            .O(N__12707),
            .I(N__12666));
    LocalMux I__2884 (
            .O(N__12700),
            .I(N__12663));
    LocalMux I__2883 (
            .O(N__12697),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__2882 (
            .O(N__12694),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__2881 (
            .O(N__12687),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__2880 (
            .O(N__12674),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__2879 (
            .O(N__12669),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    Odrv4 I__2878 (
            .O(N__12666),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    Odrv4 I__2877 (
            .O(N__12663),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    InMux I__2876 (
            .O(N__12648),
            .I(N__12645));
    LocalMux I__2875 (
            .O(N__12645),
            .I(N__12642));
    Span4Mux_h I__2874 (
            .O(N__12642),
            .I(N__12639));
    Odrv4 I__2873 (
            .O(N__12639),
            .I(\DUT.rFifoDatarx_2 ));
    InMux I__2872 (
            .O(N__12636),
            .I(N__12632));
    InMux I__2871 (
            .O(N__12635),
            .I(N__12628));
    LocalMux I__2870 (
            .O(N__12632),
            .I(N__12625));
    InMux I__2869 (
            .O(N__12631),
            .I(N__12622));
    LocalMux I__2868 (
            .O(N__12628),
            .I(N__12619));
    Span4Mux_v I__2867 (
            .O(N__12625),
            .I(N__12614));
    LocalMux I__2866 (
            .O(N__12622),
            .I(N__12614));
    Span4Mux_h I__2865 (
            .O(N__12619),
            .I(N__12610));
    Span4Mux_h I__2864 (
            .O(N__12614),
            .I(N__12607));
    InMux I__2863 (
            .O(N__12613),
            .I(N__12604));
    Odrv4 I__2862 (
            .O(N__12610),
            .I(rTxByteZ0Z_2));
    Odrv4 I__2861 (
            .O(N__12607),
            .I(rTxByteZ0Z_2));
    LocalMux I__2860 (
            .O(N__12604),
            .I(rTxByteZ0Z_2));
    CascadeMux I__2859 (
            .O(N__12597),
            .I(N__12594));
    InMux I__2858 (
            .O(N__12594),
            .I(N__12591));
    LocalMux I__2857 (
            .O(N__12591),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_2 ));
    InMux I__2856 (
            .O(N__12588),
            .I(N__12585));
    LocalMux I__2855 (
            .O(N__12585),
            .I(N__12579));
    InMux I__2854 (
            .O(N__12584),
            .I(N__12576));
    InMux I__2853 (
            .O(N__12583),
            .I(N__12573));
    InMux I__2852 (
            .O(N__12582),
            .I(N__12570));
    Span4Mux_h I__2851 (
            .O(N__12579),
            .I(N__12567));
    LocalMux I__2850 (
            .O(N__12576),
            .I(N__12562));
    LocalMux I__2849 (
            .O(N__12573),
            .I(N__12562));
    LocalMux I__2848 (
            .O(N__12570),
            .I(N__12559));
    Span4Mux_v I__2847 (
            .O(N__12567),
            .I(N__12556));
    Span4Mux_h I__2846 (
            .O(N__12562),
            .I(N__12553));
    Span4Mux_h I__2845 (
            .O(N__12559),
            .I(N__12550));
    Odrv4 I__2844 (
            .O(N__12556),
            .I(rTxByteZ0Z_6));
    Odrv4 I__2843 (
            .O(N__12553),
            .I(rTxByteZ0Z_6));
    Odrv4 I__2842 (
            .O(N__12550),
            .I(rTxByteZ0Z_6));
    InMux I__2841 (
            .O(N__12543),
            .I(N__12540));
    LocalMux I__2840 (
            .O(N__12540),
            .I(N__12537));
    Span4Mux_v I__2839 (
            .O(N__12537),
            .I(N__12534));
    Odrv4 I__2838 (
            .O(N__12534),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_6 ));
    InMux I__2837 (
            .O(N__12531),
            .I(N__12526));
    InMux I__2836 (
            .O(N__12530),
            .I(N__12523));
    InMux I__2835 (
            .O(N__12529),
            .I(N__12519));
    LocalMux I__2834 (
            .O(N__12526),
            .I(N__12514));
    LocalMux I__2833 (
            .O(N__12523),
            .I(N__12514));
    InMux I__2832 (
            .O(N__12522),
            .I(N__12511));
    LocalMux I__2831 (
            .O(N__12519),
            .I(N__12508));
    Span4Mux_v I__2830 (
            .O(N__12514),
            .I(N__12505));
    LocalMux I__2829 (
            .O(N__12511),
            .I(N__12502));
    Span4Mux_h I__2828 (
            .O(N__12508),
            .I(N__12499));
    Odrv4 I__2827 (
            .O(N__12505),
            .I(rTxByteZ0Z_7));
    Odrv4 I__2826 (
            .O(N__12502),
            .I(rTxByteZ0Z_7));
    Odrv4 I__2825 (
            .O(N__12499),
            .I(rTxByteZ0Z_7));
    InMux I__2824 (
            .O(N__12492),
            .I(N__12489));
    LocalMux I__2823 (
            .O(N__12489),
            .I(N__12486));
    Odrv4 I__2822 (
            .O(N__12486),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_7 ));
    CascadeMux I__2821 (
            .O(N__12483),
            .I(\DUT.fifo_tx_inst.N_101_cascade_ ));
    CascadeMux I__2820 (
            .O(N__12480),
            .I(N__12473));
    CascadeMux I__2819 (
            .O(N__12479),
            .I(N__12470));
    CascadeMux I__2818 (
            .O(N__12478),
            .I(N__12467));
    CascadeMux I__2817 (
            .O(N__12477),
            .I(N__12464));
    CascadeMux I__2816 (
            .O(N__12476),
            .I(N__12457));
    InMux I__2815 (
            .O(N__12473),
            .I(N__12450));
    InMux I__2814 (
            .O(N__12470),
            .I(N__12437));
    InMux I__2813 (
            .O(N__12467),
            .I(N__12437));
    InMux I__2812 (
            .O(N__12464),
            .I(N__12437));
    InMux I__2811 (
            .O(N__12463),
            .I(N__12437));
    InMux I__2810 (
            .O(N__12462),
            .I(N__12437));
    InMux I__2809 (
            .O(N__12461),
            .I(N__12437));
    InMux I__2808 (
            .O(N__12460),
            .I(N__12432));
    InMux I__2807 (
            .O(N__12457),
            .I(N__12429));
    CascadeMux I__2806 (
            .O(N__12456),
            .I(N__12425));
    CascadeMux I__2805 (
            .O(N__12455),
            .I(N__12421));
    IoInMux I__2804 (
            .O(N__12454),
            .I(N__12414));
    InMux I__2803 (
            .O(N__12453),
            .I(N__12411));
    LocalMux I__2802 (
            .O(N__12450),
            .I(N__12408));
    LocalMux I__2801 (
            .O(N__12437),
            .I(N__12405));
    InMux I__2800 (
            .O(N__12436),
            .I(N__12402));
    InMux I__2799 (
            .O(N__12435),
            .I(N__12399));
    LocalMux I__2798 (
            .O(N__12432),
            .I(N__12394));
    LocalMux I__2797 (
            .O(N__12429),
            .I(N__12394));
    InMux I__2796 (
            .O(N__12428),
            .I(N__12391));
    InMux I__2795 (
            .O(N__12425),
            .I(N__12388));
    InMux I__2794 (
            .O(N__12424),
            .I(N__12385));
    InMux I__2793 (
            .O(N__12421),
            .I(N__12382));
    CascadeMux I__2792 (
            .O(N__12420),
            .I(N__12378));
    CascadeMux I__2791 (
            .O(N__12419),
            .I(N__12375));
    CascadeMux I__2790 (
            .O(N__12418),
            .I(N__12372));
    CascadeMux I__2789 (
            .O(N__12417),
            .I(N__12369));
    LocalMux I__2788 (
            .O(N__12414),
            .I(N__12363));
    LocalMux I__2787 (
            .O(N__12411),
            .I(N__12360));
    Span4Mux_v I__2786 (
            .O(N__12408),
            .I(N__12351));
    Span4Mux_v I__2785 (
            .O(N__12405),
            .I(N__12351));
    LocalMux I__2784 (
            .O(N__12402),
            .I(N__12351));
    LocalMux I__2783 (
            .O(N__12399),
            .I(N__12351));
    Span4Mux_h I__2782 (
            .O(N__12394),
            .I(N__12340));
    LocalMux I__2781 (
            .O(N__12391),
            .I(N__12340));
    LocalMux I__2780 (
            .O(N__12388),
            .I(N__12340));
    LocalMux I__2779 (
            .O(N__12385),
            .I(N__12340));
    LocalMux I__2778 (
            .O(N__12382),
            .I(N__12340));
    InMux I__2777 (
            .O(N__12381),
            .I(N__12337));
    InMux I__2776 (
            .O(N__12378),
            .I(N__12330));
    InMux I__2775 (
            .O(N__12375),
            .I(N__12330));
    InMux I__2774 (
            .O(N__12372),
            .I(N__12330));
    InMux I__2773 (
            .O(N__12369),
            .I(N__12327));
    CascadeMux I__2772 (
            .O(N__12368),
            .I(N__12321));
    InMux I__2771 (
            .O(N__12367),
            .I(N__12317));
    InMux I__2770 (
            .O(N__12366),
            .I(N__12314));
    Span4Mux_s1_v I__2769 (
            .O(N__12363),
            .I(N__12309));
    Span4Mux_v I__2768 (
            .O(N__12360),
            .I(N__12304));
    Span4Mux_v I__2767 (
            .O(N__12351),
            .I(N__12304));
    Span4Mux_v I__2766 (
            .O(N__12340),
            .I(N__12299));
    LocalMux I__2765 (
            .O(N__12337),
            .I(N__12299));
    LocalMux I__2764 (
            .O(N__12330),
            .I(N__12293));
    LocalMux I__2763 (
            .O(N__12327),
            .I(N__12290));
    InMux I__2762 (
            .O(N__12326),
            .I(N__12283));
    InMux I__2761 (
            .O(N__12325),
            .I(N__12283));
    InMux I__2760 (
            .O(N__12324),
            .I(N__12283));
    InMux I__2759 (
            .O(N__12321),
            .I(N__12278));
    InMux I__2758 (
            .O(N__12320),
            .I(N__12278));
    LocalMux I__2757 (
            .O(N__12317),
            .I(N__12273));
    LocalMux I__2756 (
            .O(N__12314),
            .I(N__12273));
    InMux I__2755 (
            .O(N__12313),
            .I(N__12268));
    InMux I__2754 (
            .O(N__12312),
            .I(N__12268));
    Sp12to4 I__2753 (
            .O(N__12309),
            .I(N__12265));
    Span4Mux_h I__2752 (
            .O(N__12304),
            .I(N__12262));
    Span4Mux_h I__2751 (
            .O(N__12299),
            .I(N__12259));
    InMux I__2750 (
            .O(N__12298),
            .I(N__12254));
    InMux I__2749 (
            .O(N__12297),
            .I(N__12254));
    InMux I__2748 (
            .O(N__12296),
            .I(N__12251));
    Span4Mux_v I__2747 (
            .O(N__12293),
            .I(N__12246));
    Span4Mux_v I__2746 (
            .O(N__12290),
            .I(N__12246));
    LocalMux I__2745 (
            .O(N__12283),
            .I(N__12241));
    LocalMux I__2744 (
            .O(N__12278),
            .I(N__12241));
    Sp12to4 I__2743 (
            .O(N__12273),
            .I(N__12236));
    LocalMux I__2742 (
            .O(N__12268),
            .I(N__12236));
    Span12Mux_h I__2741 (
            .O(N__12265),
            .I(N__12233));
    Sp12to4 I__2740 (
            .O(N__12262),
            .I(N__12224));
    Sp12to4 I__2739 (
            .O(N__12259),
            .I(N__12224));
    LocalMux I__2738 (
            .O(N__12254),
            .I(N__12224));
    LocalMux I__2737 (
            .O(N__12251),
            .I(N__12224));
    Span4Mux_h I__2736 (
            .O(N__12246),
            .I(N__12219));
    Span4Mux_v I__2735 (
            .O(N__12241),
            .I(N__12219));
    Span12Mux_v I__2734 (
            .O(N__12236),
            .I(N__12216));
    Span12Mux_v I__2733 (
            .O(N__12233),
            .I(N__12211));
    Span12Mux_h I__2732 (
            .O(N__12224),
            .I(N__12211));
    Sp12to4 I__2731 (
            .O(N__12219),
            .I(N__12208));
    Span12Mux_h I__2730 (
            .O(N__12216),
            .I(N__12203));
    Span12Mux_v I__2729 (
            .O(N__12211),
            .I(N__12203));
    Span12Mux_h I__2728 (
            .O(N__12208),
            .I(N__12200));
    Odrv12 I__2727 (
            .O(N__12203),
            .I(wPllLocked));
    Odrv12 I__2726 (
            .O(N__12200),
            .I(wPllLocked));
    CascadeMux I__2725 (
            .O(N__12195),
            .I(\DUT.fifo_tx_inst.un1_i11_2_i_cascade_ ));
    CascadeMux I__2724 (
            .O(N__12192),
            .I(N__12172));
    InMux I__2723 (
            .O(N__12191),
            .I(N__12156));
    InMux I__2722 (
            .O(N__12190),
            .I(N__12153));
    InMux I__2721 (
            .O(N__12189),
            .I(N__12150));
    InMux I__2720 (
            .O(N__12188),
            .I(N__12147));
    InMux I__2719 (
            .O(N__12187),
            .I(N__12144));
    InMux I__2718 (
            .O(N__12186),
            .I(N__12141));
    InMux I__2717 (
            .O(N__12185),
            .I(N__12130));
    InMux I__2716 (
            .O(N__12184),
            .I(N__12130));
    InMux I__2715 (
            .O(N__12183),
            .I(N__12130));
    InMux I__2714 (
            .O(N__12182),
            .I(N__12130));
    InMux I__2713 (
            .O(N__12181),
            .I(N__12130));
    InMux I__2712 (
            .O(N__12180),
            .I(N__12125));
    InMux I__2711 (
            .O(N__12179),
            .I(N__12125));
    InMux I__2710 (
            .O(N__12178),
            .I(N__12118));
    InMux I__2709 (
            .O(N__12177),
            .I(N__12118));
    InMux I__2708 (
            .O(N__12176),
            .I(N__12118));
    InMux I__2707 (
            .O(N__12175),
            .I(N__12115));
    InMux I__2706 (
            .O(N__12172),
            .I(N__12112));
    InMux I__2705 (
            .O(N__12171),
            .I(N__12105));
    InMux I__2704 (
            .O(N__12170),
            .I(N__12105));
    InMux I__2703 (
            .O(N__12169),
            .I(N__12105));
    SRMux I__2702 (
            .O(N__12168),
            .I(N__12102));
    InMux I__2701 (
            .O(N__12167),
            .I(N__12099));
    InMux I__2700 (
            .O(N__12166),
            .I(N__12096));
    InMux I__2699 (
            .O(N__12165),
            .I(N__12093));
    InMux I__2698 (
            .O(N__12164),
            .I(N__12090));
    InMux I__2697 (
            .O(N__12163),
            .I(N__12085));
    InMux I__2696 (
            .O(N__12162),
            .I(N__12085));
    InMux I__2695 (
            .O(N__12161),
            .I(N__12082));
    InMux I__2694 (
            .O(N__12160),
            .I(N__12077));
    InMux I__2693 (
            .O(N__12159),
            .I(N__12077));
    LocalMux I__2692 (
            .O(N__12156),
            .I(N__12074));
    LocalMux I__2691 (
            .O(N__12153),
            .I(N__12071));
    LocalMux I__2690 (
            .O(N__12150),
            .I(N__12068));
    LocalMux I__2689 (
            .O(N__12147),
            .I(N__12065));
    LocalMux I__2688 (
            .O(N__12144),
            .I(N__12062));
    LocalMux I__2687 (
            .O(N__12141),
            .I(N__12059));
    LocalMux I__2686 (
            .O(N__12130),
            .I(N__12056));
    LocalMux I__2685 (
            .O(N__12125),
            .I(N__12053));
    LocalMux I__2684 (
            .O(N__12118),
            .I(N__12050));
    LocalMux I__2683 (
            .O(N__12115),
            .I(N__12047));
    LocalMux I__2682 (
            .O(N__12112),
            .I(N__12044));
    LocalMux I__2681 (
            .O(N__12105),
            .I(N__12041));
    LocalMux I__2680 (
            .O(N__12102),
            .I(N__12038));
    LocalMux I__2679 (
            .O(N__12099),
            .I(N__12035));
    LocalMux I__2678 (
            .O(N__12096),
            .I(N__12032));
    LocalMux I__2677 (
            .O(N__12093),
            .I(N__12029));
    LocalMux I__2676 (
            .O(N__12090),
            .I(N__12026));
    LocalMux I__2675 (
            .O(N__12085),
            .I(N__12023));
    LocalMux I__2674 (
            .O(N__12082),
            .I(N__12018));
    LocalMux I__2673 (
            .O(N__12077),
            .I(N__12015));
    Glb2LocalMux I__2672 (
            .O(N__12074),
            .I(N__11946));
    Glb2LocalMux I__2671 (
            .O(N__12071),
            .I(N__11946));
    Glb2LocalMux I__2670 (
            .O(N__12068),
            .I(N__11946));
    Glb2LocalMux I__2669 (
            .O(N__12065),
            .I(N__11946));
    Glb2LocalMux I__2668 (
            .O(N__12062),
            .I(N__11946));
    Glb2LocalMux I__2667 (
            .O(N__12059),
            .I(N__11946));
    Glb2LocalMux I__2666 (
            .O(N__12056),
            .I(N__11946));
    Glb2LocalMux I__2665 (
            .O(N__12053),
            .I(N__11946));
    Glb2LocalMux I__2664 (
            .O(N__12050),
            .I(N__11946));
    Glb2LocalMux I__2663 (
            .O(N__12047),
            .I(N__11946));
    Glb2LocalMux I__2662 (
            .O(N__12044),
            .I(N__11946));
    Glb2LocalMux I__2661 (
            .O(N__12041),
            .I(N__11946));
    Glb2LocalMux I__2660 (
            .O(N__12038),
            .I(N__11946));
    Glb2LocalMux I__2659 (
            .O(N__12035),
            .I(N__11946));
    Glb2LocalMux I__2658 (
            .O(N__12032),
            .I(N__11946));
    Glb2LocalMux I__2657 (
            .O(N__12029),
            .I(N__11946));
    Glb2LocalMux I__2656 (
            .O(N__12026),
            .I(N__11946));
    Glb2LocalMux I__2655 (
            .O(N__12023),
            .I(N__11946));
    CEMux I__2654 (
            .O(N__12022),
            .I(N__11946));
    CEMux I__2653 (
            .O(N__12021),
            .I(N__11946));
    Glb2LocalMux I__2652 (
            .O(N__12018),
            .I(N__11946));
    Glb2LocalMux I__2651 (
            .O(N__12015),
            .I(N__11946));
    CEMux I__2650 (
            .O(N__12014),
            .I(N__11946));
    CEMux I__2649 (
            .O(N__12013),
            .I(N__11946));
    CEMux I__2648 (
            .O(N__12012),
            .I(N__11946));
    CEMux I__2647 (
            .O(N__12011),
            .I(N__11946));
    CEMux I__2646 (
            .O(N__12010),
            .I(N__11946));
    CEMux I__2645 (
            .O(N__12009),
            .I(N__11946));
    CEMux I__2644 (
            .O(N__12008),
            .I(N__11946));
    CEMux I__2643 (
            .O(N__12007),
            .I(N__11946));
    GlobalMux I__2642 (
            .O(N__11946),
            .I(N__11943));
    gio2CtrlBuf I__2641 (
            .O(N__11943),
            .I(wPllLocked_g));
    InMux I__2640 (
            .O(N__11940),
            .I(N__11936));
    InMux I__2639 (
            .O(N__11939),
            .I(N__11933));
    LocalMux I__2638 (
            .O(N__11936),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNIIOZ0Z37 ));
    LocalMux I__2637 (
            .O(N__11933),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNIIOZ0Z37 ));
    InMux I__2636 (
            .O(N__11928),
            .I(N__11925));
    LocalMux I__2635 (
            .O(N__11925),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_6 ));
    InMux I__2634 (
            .O(N__11922),
            .I(N__11919));
    LocalMux I__2633 (
            .O(N__11919),
            .I(\DUT.fifo_tx_inst.N_101 ));
    InMux I__2632 (
            .O(N__11916),
            .I(N__11913));
    LocalMux I__2631 (
            .O(N__11913),
            .I(\DUT.fifo_tx_inst.un1_i11_2_i ));
    InMux I__2630 (
            .O(N__11910),
            .I(N__11907));
    LocalMux I__2629 (
            .O(N__11907),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_1 ));
    CascadeMux I__2628 (
            .O(N__11904),
            .I(N__11901));
    InMux I__2627 (
            .O(N__11901),
            .I(N__11898));
    LocalMux I__2626 (
            .O(N__11898),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_3 ));
    InMux I__2625 (
            .O(N__11895),
            .I(N__11892));
    LocalMux I__2624 (
            .O(N__11892),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_7 ));
    InMux I__2623 (
            .O(N__11889),
            .I(N__11886));
    LocalMux I__2622 (
            .O(N__11886),
            .I(N__11883));
    Span4Mux_v I__2621 (
            .O(N__11883),
            .I(N__11879));
    InMux I__2620 (
            .O(N__11882),
            .I(N__11876));
    Odrv4 I__2619 (
            .O(N__11879),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNIJQZ0Z47 ));
    LocalMux I__2618 (
            .O(N__11876),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNIJQZ0Z47 ));
    CascadeMux I__2617 (
            .O(N__11871),
            .I(N__11868));
    InMux I__2616 (
            .O(N__11868),
            .I(N__11865));
    LocalMux I__2615 (
            .O(N__11865),
            .I(N__11861));
    InMux I__2614 (
            .O(N__11864),
            .I(N__11858));
    Odrv4 I__2613 (
            .O(N__11861),
            .I(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_7 ));
    LocalMux I__2612 (
            .O(N__11858),
            .I(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_7 ));
    InMux I__2611 (
            .O(N__11853),
            .I(N__11849));
    InMux I__2610 (
            .O(N__11852),
            .I(N__11846));
    LocalMux I__2609 (
            .O(N__11849),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIK6NZ0Z4 ));
    LocalMux I__2608 (
            .O(N__11846),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIK6NZ0Z4 ));
    CascadeMux I__2607 (
            .O(N__11841),
            .I(N__11838));
    InMux I__2606 (
            .O(N__11838),
            .I(N__11835));
    LocalMux I__2605 (
            .O(N__11835),
            .I(N__11832));
    Odrv4 I__2604 (
            .O(N__11832),
            .I(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_4 ));
    CascadeMux I__2603 (
            .O(N__11829),
            .I(N__11826));
    InMux I__2602 (
            .O(N__11826),
            .I(N__11823));
    LocalMux I__2601 (
            .O(N__11823),
            .I(N__11819));
    CascadeMux I__2600 (
            .O(N__11822),
            .I(N__11815));
    Span4Mux_v I__2599 (
            .O(N__11819),
            .I(N__11812));
    InMux I__2598 (
            .O(N__11818),
            .I(N__11809));
    InMux I__2597 (
            .O(N__11815),
            .I(N__11806));
    Odrv4 I__2596 (
            .O(N__11812),
            .I(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_5 ));
    LocalMux I__2595 (
            .O(N__11809),
            .I(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_5 ));
    LocalMux I__2594 (
            .O(N__11806),
            .I(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_5 ));
    CascadeMux I__2593 (
            .O(N__11799),
            .I(N__11796));
    InMux I__2592 (
            .O(N__11796),
            .I(N__11792));
    InMux I__2591 (
            .O(N__11795),
            .I(N__11789));
    LocalMux I__2590 (
            .O(N__11792),
            .I(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_2 ));
    LocalMux I__2589 (
            .O(N__11789),
            .I(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_2 ));
    CascadeMux I__2588 (
            .O(N__11784),
            .I(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_4_cascade_ ));
    InMux I__2587 (
            .O(N__11781),
            .I(N__11778));
    LocalMux I__2586 (
            .O(N__11778),
            .I(\fifo_inst.tx_fifo_inst.un18_rRamWrAddr_5 ));
    CascadeMux I__2585 (
            .O(N__11775),
            .I(N__11772));
    InMux I__2584 (
            .O(N__11772),
            .I(N__11769));
    LocalMux I__2583 (
            .O(N__11769),
            .I(N__11766));
    Odrv4 I__2582 (
            .O(N__11766),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_1 ));
    CascadeMux I__2581 (
            .O(N__11763),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_1_cascade_ ));
    CascadeMux I__2580 (
            .O(N__11760),
            .I(N__11757));
    InMux I__2579 (
            .O(N__11757),
            .I(N__11754));
    LocalMux I__2578 (
            .O(N__11754),
            .I(N__11750));
    InMux I__2577 (
            .O(N__11753),
            .I(N__11746));
    Span4Mux_v I__2576 (
            .O(N__11750),
            .I(N__11741));
    InMux I__2575 (
            .O(N__11749),
            .I(N__11738));
    LocalMux I__2574 (
            .O(N__11746),
            .I(N__11735));
    InMux I__2573 (
            .O(N__11745),
            .I(N__11732));
    InMux I__2572 (
            .O(N__11744),
            .I(N__11729));
    Odrv4 I__2571 (
            .O(N__11741),
            .I(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_0 ));
    LocalMux I__2570 (
            .O(N__11738),
            .I(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_0 ));
    Odrv4 I__2569 (
            .O(N__11735),
            .I(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_0 ));
    LocalMux I__2568 (
            .O(N__11732),
            .I(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_0 ));
    LocalMux I__2567 (
            .O(N__11729),
            .I(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_0 ));
    InMux I__2566 (
            .O(N__11718),
            .I(N__11715));
    LocalMux I__2565 (
            .O(N__11715),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIZ0 ));
    CascadeMux I__2564 (
            .O(N__11712),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIZ0_cascade_ ));
    CascadeMux I__2563 (
            .O(N__11709),
            .I(N__11706));
    InMux I__2562 (
            .O(N__11706),
            .I(N__11703));
    LocalMux I__2561 (
            .O(N__11703),
            .I(N__11699));
    InMux I__2560 (
            .O(N__11702),
            .I(N__11696));
    Odrv4 I__2559 (
            .O(N__11699),
            .I(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_1 ));
    LocalMux I__2558 (
            .O(N__11696),
            .I(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_1 ));
    InMux I__2557 (
            .O(N__11691),
            .I(N__11688));
    LocalMux I__2556 (
            .O(N__11688),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7 ));
    InMux I__2555 (
            .O(N__11685),
            .I(N__11681));
    InMux I__2554 (
            .O(N__11684),
            .I(N__11678));
    LocalMux I__2553 (
            .O(N__11681),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddr_rst_4 ));
    LocalMux I__2552 (
            .O(N__11678),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddr_rst_4 ));
    InMux I__2551 (
            .O(N__11673),
            .I(N__11670));
    LocalMux I__2550 (
            .O(N__11670),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddr_0_5 ));
    CascadeMux I__2549 (
            .O(N__11667),
            .I(N__11664));
    InMux I__2548 (
            .O(N__11664),
            .I(N__11661));
    LocalMux I__2547 (
            .O(N__11661),
            .I(N__11656));
    InMux I__2546 (
            .O(N__11660),
            .I(N__11653));
    CascadeMux I__2545 (
            .O(N__11659),
            .I(N__11650));
    Span4Mux_v I__2544 (
            .O(N__11656),
            .I(N__11645));
    LocalMux I__2543 (
            .O(N__11653),
            .I(N__11645));
    InMux I__2542 (
            .O(N__11650),
            .I(N__11642));
    Odrv4 I__2541 (
            .O(N__11645),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_5 ));
    LocalMux I__2540 (
            .O(N__11642),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_5 ));
    InMux I__2539 (
            .O(N__11637),
            .I(N__11634));
    LocalMux I__2538 (
            .O(N__11634),
            .I(N__11631));
    Odrv4 I__2537 (
            .O(N__11631),
            .I(\fifo_inst.tx_fifo_inst.un18_rRamWrAddr_4 ));
    InMux I__2536 (
            .O(N__11628),
            .I(N__11624));
    InMux I__2535 (
            .O(N__11627),
            .I(N__11621));
    LocalMux I__2534 (
            .O(N__11624),
            .I(N__11617));
    LocalMux I__2533 (
            .O(N__11621),
            .I(N__11614));
    InMux I__2532 (
            .O(N__11620),
            .I(N__11611));
    Odrv12 I__2531 (
            .O(N__11617),
            .I(\fifo_inst.tx_fifo_inst.un18_rRamWrAddr ));
    Odrv4 I__2530 (
            .O(N__11614),
            .I(\fifo_inst.tx_fifo_inst.un18_rRamWrAddr ));
    LocalMux I__2529 (
            .O(N__11611),
            .I(\fifo_inst.tx_fifo_inst.un18_rRamWrAddr ));
    InMux I__2528 (
            .O(N__11604),
            .I(N__11601));
    LocalMux I__2527 (
            .O(N__11601),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_2 ));
    InMux I__2526 (
            .O(N__11598),
            .I(N__11594));
    InMux I__2525 (
            .O(N__11597),
            .I(N__11591));
    LocalMux I__2524 (
            .O(N__11594),
            .I(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI6IZ0Z12 ));
    LocalMux I__2523 (
            .O(N__11591),
            .I(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI6IZ0Z12 ));
    InMux I__2522 (
            .O(N__11586),
            .I(N__11583));
    LocalMux I__2521 (
            .O(N__11583),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddr_0_3 ));
    InMux I__2520 (
            .O(N__11580),
            .I(N__11570));
    InMux I__2519 (
            .O(N__11579),
            .I(N__11570));
    InMux I__2518 (
            .O(N__11578),
            .I(N__11567));
    InMux I__2517 (
            .O(N__11577),
            .I(N__11564));
    InMux I__2516 (
            .O(N__11576),
            .I(N__11559));
    InMux I__2515 (
            .O(N__11575),
            .I(N__11559));
    LocalMux I__2514 (
            .O(N__11570),
            .I(N__11556));
    LocalMux I__2513 (
            .O(N__11567),
            .I(\fifo_inst.rTxRdEn_fast ));
    LocalMux I__2512 (
            .O(N__11564),
            .I(\fifo_inst.rTxRdEn_fast ));
    LocalMux I__2511 (
            .O(N__11559),
            .I(\fifo_inst.rTxRdEn_fast ));
    Odrv4 I__2510 (
            .O(N__11556),
            .I(\fifo_inst.rTxRdEn_fast ));
    CascadeMux I__2509 (
            .O(N__11547),
            .I(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI20CZ0Z4_cascade_ ));
    CascadeMux I__2508 (
            .O(N__11544),
            .I(N__11540));
    InMux I__2507 (
            .O(N__11543),
            .I(N__11537));
    InMux I__2506 (
            .O(N__11540),
            .I(N__11533));
    LocalMux I__2505 (
            .O(N__11537),
            .I(N__11530));
    InMux I__2504 (
            .O(N__11536),
            .I(N__11527));
    LocalMux I__2503 (
            .O(N__11533),
            .I(\fifo_inst.tx_fifo_inst.un15_rRamRdAddr ));
    Odrv4 I__2502 (
            .O(N__11530),
            .I(\fifo_inst.tx_fifo_inst.un15_rRamRdAddr ));
    LocalMux I__2501 (
            .O(N__11527),
            .I(\fifo_inst.tx_fifo_inst.un15_rRamRdAddr ));
    CascadeMux I__2500 (
            .O(N__11520),
            .I(N__11517));
    InMux I__2499 (
            .O(N__11517),
            .I(N__11513));
    CascadeMux I__2498 (
            .O(N__11516),
            .I(N__11510));
    LocalMux I__2497 (
            .O(N__11513),
            .I(N__11507));
    InMux I__2496 (
            .O(N__11510),
            .I(N__11504));
    Odrv4 I__2495 (
            .O(N__11507),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_3 ));
    LocalMux I__2494 (
            .O(N__11504),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_3 ));
    CascadeMux I__2493 (
            .O(N__11499),
            .I(N__11496));
    InMux I__2492 (
            .O(N__11496),
            .I(N__11491));
    CascadeMux I__2491 (
            .O(N__11495),
            .I(N__11488));
    InMux I__2490 (
            .O(N__11494),
            .I(N__11483));
    LocalMux I__2489 (
            .O(N__11491),
            .I(N__11480));
    InMux I__2488 (
            .O(N__11488),
            .I(N__11477));
    InMux I__2487 (
            .O(N__11487),
            .I(N__11473));
    InMux I__2486 (
            .O(N__11486),
            .I(N__11470));
    LocalMux I__2485 (
            .O(N__11483),
            .I(N__11467));
    Span4Mux_h I__2484 (
            .O(N__11480),
            .I(N__11462));
    LocalMux I__2483 (
            .O(N__11477),
            .I(N__11462));
    InMux I__2482 (
            .O(N__11476),
            .I(N__11459));
    LocalMux I__2481 (
            .O(N__11473),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_0 ));
    LocalMux I__2480 (
            .O(N__11470),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_0 ));
    Odrv4 I__2479 (
            .O(N__11467),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_0 ));
    Odrv4 I__2478 (
            .O(N__11462),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_0 ));
    LocalMux I__2477 (
            .O(N__11459),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_0 ));
    CascadeMux I__2476 (
            .O(N__11448),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_3_cascade_ ));
    CascadeMux I__2475 (
            .O(N__11445),
            .I(N__11440));
    InMux I__2474 (
            .O(N__11444),
            .I(N__11437));
    InMux I__2473 (
            .O(N__11443),
            .I(N__11434));
    InMux I__2472 (
            .O(N__11440),
            .I(N__11431));
    LocalMux I__2471 (
            .O(N__11437),
            .I(N__11428));
    LocalMux I__2470 (
            .O(N__11434),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_8 ));
    LocalMux I__2469 (
            .O(N__11431),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_8 ));
    Odrv4 I__2468 (
            .O(N__11428),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_8 ));
    CascadeMux I__2467 (
            .O(N__11421),
            .I(N__11418));
    InMux I__2466 (
            .O(N__11418),
            .I(N__11415));
    LocalMux I__2465 (
            .O(N__11415),
            .I(\fifo_inst.tx_fifo_inst.un15_rRamRdAddr_4 ));
    InMux I__2464 (
            .O(N__11412),
            .I(N__11406));
    InMux I__2463 (
            .O(N__11411),
            .I(N__11406));
    LocalMux I__2462 (
            .O(N__11406),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNII2LZ0Z4 ));
    CascadeMux I__2461 (
            .O(N__11403),
            .I(N__11399));
    CascadeMux I__2460 (
            .O(N__11402),
            .I(N__11396));
    InMux I__2459 (
            .O(N__11399),
            .I(N__11393));
    InMux I__2458 (
            .O(N__11396),
            .I(N__11390));
    LocalMux I__2457 (
            .O(N__11393),
            .I(N__11387));
    LocalMux I__2456 (
            .O(N__11390),
            .I(N__11384));
    Odrv4 I__2455 (
            .O(N__11387),
            .I(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_6 ));
    Odrv4 I__2454 (
            .O(N__11384),
            .I(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_6 ));
    CascadeMux I__2453 (
            .O(N__11379),
            .I(\DUT.fifo_tx_inst.rFifoData_awe3_cascade_ ));
    CascadeMux I__2452 (
            .O(N__11376),
            .I(N__11373));
    InMux I__2451 (
            .O(N__11373),
            .I(N__11370));
    LocalMux I__2450 (
            .O(N__11370),
            .I(\DUT.fifo_tx_inst.un1_i11_i ));
    CascadeMux I__2449 (
            .O(N__11367),
            .I(\DUT.fifo_tx_inst.un1_i11_i_cascade_ ));
    InMux I__2448 (
            .O(N__11364),
            .I(N__11357));
    InMux I__2447 (
            .O(N__11363),
            .I(N__11354));
    InMux I__2446 (
            .O(N__11362),
            .I(N__11347));
    InMux I__2445 (
            .O(N__11361),
            .I(N__11347));
    InMux I__2444 (
            .O(N__11360),
            .I(N__11347));
    LocalMux I__2443 (
            .O(N__11357),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_1 ));
    LocalMux I__2442 (
            .O(N__11354),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_1 ));
    LocalMux I__2441 (
            .O(N__11347),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_1 ));
    CascadeMux I__2440 (
            .O(N__11340),
            .I(N__11332));
    CascadeMux I__2439 (
            .O(N__11339),
            .I(N__11329));
    InMux I__2438 (
            .O(N__11338),
            .I(N__11324));
    InMux I__2437 (
            .O(N__11337),
            .I(N__11324));
    InMux I__2436 (
            .O(N__11336),
            .I(N__11315));
    InMux I__2435 (
            .O(N__11335),
            .I(N__11315));
    InMux I__2434 (
            .O(N__11332),
            .I(N__11315));
    InMux I__2433 (
            .O(N__11329),
            .I(N__11315));
    LocalMux I__2432 (
            .O(N__11324),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_0 ));
    LocalMux I__2431 (
            .O(N__11315),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_0 ));
    InMux I__2430 (
            .O(N__11310),
            .I(N__11306));
    InMux I__2429 (
            .O(N__11309),
            .I(N__11303));
    LocalMux I__2428 (
            .O(N__11306),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddr_rst_7 ));
    LocalMux I__2427 (
            .O(N__11303),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddr_rst_7 ));
    InMux I__2426 (
            .O(N__11298),
            .I(N__11295));
    LocalMux I__2425 (
            .O(N__11295),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddr_0_8 ));
    CEMux I__2424 (
            .O(N__11292),
            .I(N__11289));
    LocalMux I__2423 (
            .O(N__11289),
            .I(N__11284));
    CEMux I__2422 (
            .O(N__11288),
            .I(N__11281));
    CEMux I__2421 (
            .O(N__11287),
            .I(N__11278));
    Span4Mux_v I__2420 (
            .O(N__11284),
            .I(N__11275));
    LocalMux I__2419 (
            .O(N__11281),
            .I(N__11272));
    LocalMux I__2418 (
            .O(N__11278),
            .I(N__11269));
    Span4Mux_h I__2417 (
            .O(N__11275),
            .I(N__11266));
    Sp12to4 I__2416 (
            .O(N__11272),
            .I(N__11261));
    Sp12to4 I__2415 (
            .O(N__11269),
            .I(N__11261));
    Odrv4 I__2414 (
            .O(N__11266),
            .I(\fifo_inst.rTxRdEn_RNIS0VN ));
    Odrv12 I__2413 (
            .O(N__11261),
            .I(\fifo_inst.rTxRdEn_RNIS0VN ));
    InMux I__2412 (
            .O(N__11256),
            .I(N__11253));
    LocalMux I__2411 (
            .O(N__11253),
            .I(N__11250));
    Odrv4 I__2410 (
            .O(N__11250),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_3 ));
    InMux I__2409 (
            .O(N__11247),
            .I(N__11244));
    LocalMux I__2408 (
            .O(N__11244),
            .I(N__11238));
    InMux I__2407 (
            .O(N__11243),
            .I(N__11235));
    InMux I__2406 (
            .O(N__11242),
            .I(N__11232));
    InMux I__2405 (
            .O(N__11241),
            .I(N__11229));
    Span4Mux_h I__2404 (
            .O(N__11238),
            .I(N__11226));
    LocalMux I__2403 (
            .O(N__11235),
            .I(N__11223));
    LocalMux I__2402 (
            .O(N__11232),
            .I(N__11218));
    LocalMux I__2401 (
            .O(N__11229),
            .I(N__11218));
    Sp12to4 I__2400 (
            .O(N__11226),
            .I(N__11215));
    Span4Mux_h I__2399 (
            .O(N__11223),
            .I(N__11212));
    Span4Mux_h I__2398 (
            .O(N__11218),
            .I(N__11209));
    Odrv12 I__2397 (
            .O(N__11215),
            .I(rTxByteZ0Z_4));
    Odrv4 I__2396 (
            .O(N__11212),
            .I(rTxByteZ0Z_4));
    Odrv4 I__2395 (
            .O(N__11209),
            .I(rTxByteZ0Z_4));
    InMux I__2394 (
            .O(N__11202),
            .I(N__11199));
    LocalMux I__2393 (
            .O(N__11199),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_4 ));
    InMux I__2392 (
            .O(N__11196),
            .I(N__11193));
    LocalMux I__2391 (
            .O(N__11193),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_1 ));
    InMux I__2390 (
            .O(N__11190),
            .I(N__11187));
    LocalMux I__2389 (
            .O(N__11187),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_6 ));
    CascadeMux I__2388 (
            .O(N__11184),
            .I(N__11181));
    InMux I__2387 (
            .O(N__11181),
            .I(N__11178));
    LocalMux I__2386 (
            .O(N__11178),
            .I(N__11175));
    Odrv4 I__2385 (
            .O(N__11175),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_7 ));
    InMux I__2384 (
            .O(N__11172),
            .I(N__11168));
    InMux I__2383 (
            .O(N__11171),
            .I(N__11165));
    LocalMux I__2382 (
            .O(N__11168),
            .I(N__11162));
    LocalMux I__2381 (
            .O(N__11165),
            .I(\DUT.fifo_tx_inst.rFifoDataro_1 ));
    Odrv4 I__2380 (
            .O(N__11162),
            .I(\DUT.fifo_tx_inst.rFifoDataro_1 ));
    CEMux I__2379 (
            .O(N__11157),
            .I(N__11153));
    CEMux I__2378 (
            .O(N__11156),
            .I(N__11150));
    LocalMux I__2377 (
            .O(N__11153),
            .I(N__11147));
    LocalMux I__2376 (
            .O(N__11150),
            .I(N__11144));
    Odrv4 I__2375 (
            .O(N__11147),
            .I(\DUT.fifo_tx_inst.rFifoData_awe2 ));
    Odrv4 I__2374 (
            .O(N__11144),
            .I(\DUT.fifo_tx_inst.rFifoData_awe2 ));
    CascadeMux I__2373 (
            .O(N__11139),
            .I(\DUT.fifo_tx_inst.rFifoData_awe2_cascade_ ));
    InMux I__2372 (
            .O(N__11136),
            .I(N__11132));
    InMux I__2371 (
            .O(N__11135),
            .I(N__11129));
    LocalMux I__2370 (
            .O(N__11132),
            .I(N__11126));
    LocalMux I__2369 (
            .O(N__11129),
            .I(\DUT.fifo_tx_inst.rFifoDataro_2 ));
    Odrv4 I__2368 (
            .O(N__11126),
            .I(\DUT.fifo_tx_inst.rFifoDataro_2 ));
    CascadeMux I__2367 (
            .O(N__11121),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ));
    InMux I__2366 (
            .O(N__11118),
            .I(N__11115));
    LocalMux I__2365 (
            .O(N__11115),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_5 ));
    CascadeMux I__2364 (
            .O(N__11112),
            .I(N__11109));
    InMux I__2363 (
            .O(N__11109),
            .I(N__11106));
    LocalMux I__2362 (
            .O(N__11106),
            .I(\DUT.rFifoDatarx_5 ));
    InMux I__2361 (
            .O(N__11103),
            .I(N__11100));
    LocalMux I__2360 (
            .O(N__11100),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_1 ));
    CascadeMux I__2359 (
            .O(N__11097),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1_cascade_ ));
    CascadeMux I__2358 (
            .O(N__11094),
            .I(N__11091));
    InMux I__2357 (
            .O(N__11091),
            .I(N__11088));
    LocalMux I__2356 (
            .O(N__11088),
            .I(N__11085));
    Odrv4 I__2355 (
            .O(N__11085),
            .I(\DUT.rFifoDatarx_1 ));
    InMux I__2354 (
            .O(N__11082),
            .I(N__11079));
    LocalMux I__2353 (
            .O(N__11079),
            .I(N__11075));
    InMux I__2352 (
            .O(N__11078),
            .I(N__11072));
    Span4Mux_h I__2351 (
            .O(N__11075),
            .I(N__11069));
    LocalMux I__2350 (
            .O(N__11072),
            .I(\DUT.fifo_tx_inst.rFifoDataro_0 ));
    Odrv4 I__2349 (
            .O(N__11069),
            .I(\DUT.fifo_tx_inst.rFifoDataro_0 ));
    CascadeMux I__2348 (
            .O(N__11064),
            .I(\DUT.fifo_tx_inst.rFifoDataror_1_0_cascade_ ));
    CascadeMux I__2347 (
            .O(N__11061),
            .I(N__11056));
    InMux I__2346 (
            .O(N__11060),
            .I(N__11042));
    InMux I__2345 (
            .O(N__11059),
            .I(N__11042));
    InMux I__2344 (
            .O(N__11056),
            .I(N__11042));
    InMux I__2343 (
            .O(N__11055),
            .I(N__11042));
    InMux I__2342 (
            .O(N__11054),
            .I(N__11033));
    InMux I__2341 (
            .O(N__11053),
            .I(N__11033));
    InMux I__2340 (
            .O(N__11052),
            .I(N__11033));
    InMux I__2339 (
            .O(N__11051),
            .I(N__11033));
    LocalMux I__2338 (
            .O(N__11042),
            .I(N__11030));
    LocalMux I__2337 (
            .O(N__11033),
            .I(\DUT.rFifoDataror_0 ));
    Odrv4 I__2336 (
            .O(N__11030),
            .I(\DUT.rFifoDataror_0 ));
    InMux I__2335 (
            .O(N__11025),
            .I(N__11022));
    LocalMux I__2334 (
            .O(N__11022),
            .I(N__11019));
    Odrv4 I__2333 (
            .O(N__11019),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_0 ));
    InMux I__2332 (
            .O(N__11016),
            .I(N__11013));
    LocalMux I__2331 (
            .O(N__11013),
            .I(N__11010));
    Odrv4 I__2330 (
            .O(N__11010),
            .I(\DUT.rFifoDatarxZ0Z_0 ));
    CascadeMux I__2329 (
            .O(N__11007),
            .I(N__11004));
    InMux I__2328 (
            .O(N__11004),
            .I(N__11001));
    LocalMux I__2327 (
            .O(N__11001),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_0 ));
    InMux I__2326 (
            .O(N__10998),
            .I(N__10995));
    LocalMux I__2325 (
            .O(N__10995),
            .I(N__10992));
    Odrv4 I__2324 (
            .O(N__10992),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_5 ));
    InMux I__2323 (
            .O(N__10989),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_4 ));
    InMux I__2322 (
            .O(N__10986),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5 ));
    InMux I__2321 (
            .O(N__10983),
            .I(N__10980));
    LocalMux I__2320 (
            .O(N__10980),
            .I(N__10977));
    Span4Mux_v I__2319 (
            .O(N__10977),
            .I(N__10974));
    Odrv4 I__2318 (
            .O(N__10974),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_7 ));
    InMux I__2317 (
            .O(N__10971),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6 ));
    InMux I__2316 (
            .O(N__10968),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_7 ));
    CascadeMux I__2315 (
            .O(N__10965),
            .I(N__10962));
    InMux I__2314 (
            .O(N__10962),
            .I(N__10958));
    InMux I__2313 (
            .O(N__10961),
            .I(N__10955));
    LocalMux I__2312 (
            .O(N__10958),
            .I(N__10952));
    LocalMux I__2311 (
            .O(N__10955),
            .I(N__10949));
    Span4Mux_v I__2310 (
            .O(N__10952),
            .I(N__10943));
    Span4Mux_v I__2309 (
            .O(N__10949),
            .I(N__10943));
    InMux I__2308 (
            .O(N__10948),
            .I(N__10940));
    Odrv4 I__2307 (
            .O(N__10943),
            .I(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_8 ));
    LocalMux I__2306 (
            .O(N__10940),
            .I(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_8 ));
    CascadeMux I__2305 (
            .O(N__10935),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ));
    InMux I__2304 (
            .O(N__10932),
            .I(N__10929));
    LocalMux I__2303 (
            .O(N__10929),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_3 ));
    InMux I__2302 (
            .O(N__10926),
            .I(N__10923));
    LocalMux I__2301 (
            .O(N__10923),
            .I(\DUT.rFifoDatarx_3 ));
    InMux I__2300 (
            .O(N__10920),
            .I(N__10917));
    LocalMux I__2299 (
            .O(N__10917),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_4 ));
    InMux I__2298 (
            .O(N__10914),
            .I(N__10911));
    LocalMux I__2297 (
            .O(N__10911),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_7 ));
    InMux I__2296 (
            .O(N__10908),
            .I(N__10905));
    LocalMux I__2295 (
            .O(N__10905),
            .I(\DUT.rFifoDatarx_7 ));
    InMux I__2294 (
            .O(N__10902),
            .I(N__10899));
    LocalMux I__2293 (
            .O(N__10899),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_5 ));
    InMux I__2292 (
            .O(N__10896),
            .I(N__10893));
    LocalMux I__2291 (
            .O(N__10893),
            .I(\fifo_inst.ft2232h_inst.rFifoState_RNIG8PKZ0Z_4 ));
    CascadeMux I__2290 (
            .O(N__10890),
            .I(N__10886));
    InMux I__2289 (
            .O(N__10889),
            .I(N__10883));
    InMux I__2288 (
            .O(N__10886),
            .I(N__10879));
    LocalMux I__2287 (
            .O(N__10883),
            .I(N__10876));
    CascadeMux I__2286 (
            .O(N__10882),
            .I(N__10873));
    LocalMux I__2285 (
            .O(N__10879),
            .I(N__10870));
    Span4Mux_h I__2284 (
            .O(N__10876),
            .I(N__10867));
    InMux I__2283 (
            .O(N__10873),
            .I(N__10864));
    Odrv4 I__2282 (
            .O(N__10870),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_7 ));
    Odrv4 I__2281 (
            .O(N__10867),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_7 ));
    LocalMux I__2280 (
            .O(N__10864),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_7 ));
    CascadeMux I__2279 (
            .O(N__10857),
            .I(N__10854));
    InMux I__2278 (
            .O(N__10854),
            .I(N__10849));
    InMux I__2277 (
            .O(N__10853),
            .I(N__10846));
    CascadeMux I__2276 (
            .O(N__10852),
            .I(N__10843));
    LocalMux I__2275 (
            .O(N__10849),
            .I(N__10840));
    LocalMux I__2274 (
            .O(N__10846),
            .I(N__10837));
    InMux I__2273 (
            .O(N__10843),
            .I(N__10834));
    Odrv4 I__2272 (
            .O(N__10840),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_6 ));
    Odrv4 I__2271 (
            .O(N__10837),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_6 ));
    LocalMux I__2270 (
            .O(N__10834),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_6 ));
    InMux I__2269 (
            .O(N__10827),
            .I(N__10824));
    LocalMux I__2268 (
            .O(N__10824),
            .I(\fifo_inst.tx_fifo_inst.un15_rRamRdAddr_5 ));
    CascadeMux I__2267 (
            .O(N__10821),
            .I(\fifo_inst.tx_fifo_inst.un15_rRamRdAddr_cascade_ ));
    InMux I__2266 (
            .O(N__10818),
            .I(N__10815));
    LocalMux I__2265 (
            .O(N__10815),
            .I(N__10812));
    Odrv4 I__2264 (
            .O(N__10812),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddr_0_0 ));
    CascadeMux I__2263 (
            .O(N__10809),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddr_rst_cascade_ ));
    InMux I__2262 (
            .O(N__10806),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1 ));
    InMux I__2261 (
            .O(N__10803),
            .I(N__10800));
    LocalMux I__2260 (
            .O(N__10800),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_3 ));
    InMux I__2259 (
            .O(N__10797),
            .I(N__10794));
    LocalMux I__2258 (
            .O(N__10794),
            .I(N__10791));
    Span4Mux_v I__2257 (
            .O(N__10791),
            .I(N__10787));
    InMux I__2256 (
            .O(N__10790),
            .I(N__10784));
    Odrv4 I__2255 (
            .O(N__10787),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIJ4MZ0Z4 ));
    LocalMux I__2254 (
            .O(N__10784),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIJ4MZ0Z4 ));
    InMux I__2253 (
            .O(N__10779),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2 ));
    InMux I__2252 (
            .O(N__10776),
            .I(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3 ));
    CascadeMux I__2251 (
            .O(N__10773),
            .I(N__10770));
    InMux I__2250 (
            .O(N__10770),
            .I(N__10767));
    LocalMux I__2249 (
            .O(N__10767),
            .I(N__10763));
    CascadeMux I__2248 (
            .O(N__10766),
            .I(N__10759));
    Span4Mux_v I__2247 (
            .O(N__10763),
            .I(N__10756));
    InMux I__2246 (
            .O(N__10762),
            .I(N__10753));
    InMux I__2245 (
            .O(N__10759),
            .I(N__10750));
    Odrv4 I__2244 (
            .O(N__10756),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_2 ));
    LocalMux I__2243 (
            .O(N__10753),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_2 ));
    LocalMux I__2242 (
            .O(N__10750),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_2 ));
    InMux I__2241 (
            .O(N__10743),
            .I(N__10737));
    InMux I__2240 (
            .O(N__10742),
            .I(N__10737));
    LocalMux I__2239 (
            .O(N__10737),
            .I(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1_c_RNI5GZ0Z02 ));
    InMux I__2238 (
            .O(N__10734),
            .I(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1 ));
    InMux I__2237 (
            .O(N__10731),
            .I(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2 ));
    CascadeMux I__2236 (
            .O(N__10728),
            .I(N__10725));
    InMux I__2235 (
            .O(N__10725),
            .I(N__10721));
    InMux I__2234 (
            .O(N__10724),
            .I(N__10717));
    LocalMux I__2233 (
            .O(N__10721),
            .I(N__10714));
    InMux I__2232 (
            .O(N__10720),
            .I(N__10711));
    LocalMux I__2231 (
            .O(N__10717),
            .I(N__10708));
    Odrv4 I__2230 (
            .O(N__10714),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_4 ));
    LocalMux I__2229 (
            .O(N__10711),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_4 ));
    Odrv4 I__2228 (
            .O(N__10708),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_4 ));
    InMux I__2227 (
            .O(N__10701),
            .I(N__10695));
    InMux I__2226 (
            .O(N__10700),
            .I(N__10695));
    LocalMux I__2225 (
            .O(N__10695),
            .I(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_3_c_RNI7KZ0Z22 ));
    InMux I__2224 (
            .O(N__10692),
            .I(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_3 ));
    InMux I__2223 (
            .O(N__10689),
            .I(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_4 ));
    InMux I__2222 (
            .O(N__10686),
            .I(N__10680));
    InMux I__2221 (
            .O(N__10685),
            .I(N__10680));
    LocalMux I__2220 (
            .O(N__10680),
            .I(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_5_c_RNI9OZ0Z42 ));
    InMux I__2219 (
            .O(N__10677),
            .I(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_5 ));
    InMux I__2218 (
            .O(N__10674),
            .I(N__10668));
    InMux I__2217 (
            .O(N__10673),
            .I(N__10668));
    LocalMux I__2216 (
            .O(N__10668),
            .I(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_6_c_RNIAQZ0Z52 ));
    InMux I__2215 (
            .O(N__10665),
            .I(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_6 ));
    InMux I__2214 (
            .O(N__10662),
            .I(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_7 ));
    InMux I__2213 (
            .O(N__10659),
            .I(N__10656));
    LocalMux I__2212 (
            .O(N__10656),
            .I(N__10653));
    Odrv4 I__2211 (
            .O(N__10653),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_4 ));
    InMux I__2210 (
            .O(N__10650),
            .I(N__10647));
    LocalMux I__2209 (
            .O(N__10647),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddr_0_7 ));
    InMux I__2208 (
            .O(N__10644),
            .I(N__10641));
    LocalMux I__2207 (
            .O(N__10641),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddr_0_4 ));
    InMux I__2206 (
            .O(N__10638),
            .I(N__10635));
    LocalMux I__2205 (
            .O(N__10635),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddr_0_6 ));
    InMux I__2204 (
            .O(N__10632),
            .I(N__10629));
    LocalMux I__2203 (
            .O(N__10629),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_1_1 ));
    CascadeMux I__2202 (
            .O(N__10626),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_ ));
    CascadeMux I__2201 (
            .O(N__10623),
            .I(N__10620));
    InMux I__2200 (
            .O(N__10620),
            .I(N__10617));
    LocalMux I__2199 (
            .O(N__10617),
            .I(N__10614));
    Span4Mux_h I__2198 (
            .O(N__10614),
            .I(N__10611));
    Odrv4 I__2197 (
            .O(N__10611),
            .I(\DUT.rFifoDatarx_4 ));
    InMux I__2196 (
            .O(N__10608),
            .I(N__10605));
    LocalMux I__2195 (
            .O(N__10605),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_4 ));
    CascadeMux I__2194 (
            .O(N__10602),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_ ));
    InMux I__2193 (
            .O(N__10599),
            .I(N__10596));
    LocalMux I__2192 (
            .O(N__10596),
            .I(N__10593));
    Odrv12 I__2191 (
            .O(N__10593),
            .I(\DUT.rFifoDatarx_6 ));
    InMux I__2190 (
            .O(N__10590),
            .I(N__10587));
    LocalMux I__2189 (
            .O(N__10587),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_4 ));
    InMux I__2188 (
            .O(N__10584),
            .I(N__10581));
    LocalMux I__2187 (
            .O(N__10581),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_6 ));
    InMux I__2186 (
            .O(N__10578),
            .I(N__10575));
    LocalMux I__2185 (
            .O(N__10575),
            .I(N__10572));
    Odrv4 I__2184 (
            .O(N__10572),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_6 ));
    InMux I__2183 (
            .O(N__10569),
            .I(N__10566));
    LocalMux I__2182 (
            .O(N__10566),
            .I(N__10563));
    Odrv4 I__2181 (
            .O(N__10563),
            .I(\DUT.uart_inst0.tx_dataZ0Z_4 ));
    InMux I__2180 (
            .O(N__10560),
            .I(N__10557));
    LocalMux I__2179 (
            .O(N__10557),
            .I(\DUT.uart_inst0.tx_dataZ0Z_7 ));
    InMux I__2178 (
            .O(N__10554),
            .I(N__10551));
    LocalMux I__2177 (
            .O(N__10551),
            .I(\DUT.uart_inst0.tx_dataZ0Z_6 ));
    CascadeMux I__2176 (
            .O(N__10548),
            .I(N__10540));
    CascadeMux I__2175 (
            .O(N__10547),
            .I(N__10530));
    CascadeMux I__2174 (
            .O(N__10546),
            .I(N__10527));
    InMux I__2173 (
            .O(N__10545),
            .I(N__10523));
    InMux I__2172 (
            .O(N__10544),
            .I(N__10516));
    InMux I__2171 (
            .O(N__10543),
            .I(N__10516));
    InMux I__2170 (
            .O(N__10540),
            .I(N__10516));
    InMux I__2169 (
            .O(N__10539),
            .I(N__10513));
    InMux I__2168 (
            .O(N__10538),
            .I(N__10510));
    InMux I__2167 (
            .O(N__10537),
            .I(N__10504));
    InMux I__2166 (
            .O(N__10536),
            .I(N__10504));
    CascadeMux I__2165 (
            .O(N__10535),
            .I(N__10495));
    CascadeMux I__2164 (
            .O(N__10534),
            .I(N__10492));
    InMux I__2163 (
            .O(N__10533),
            .I(N__10481));
    InMux I__2162 (
            .O(N__10530),
            .I(N__10481));
    InMux I__2161 (
            .O(N__10527),
            .I(N__10481));
    InMux I__2160 (
            .O(N__10526),
            .I(N__10481));
    LocalMux I__2159 (
            .O(N__10523),
            .I(N__10476));
    LocalMux I__2158 (
            .O(N__10516),
            .I(N__10476));
    LocalMux I__2157 (
            .O(N__10513),
            .I(N__10472));
    LocalMux I__2156 (
            .O(N__10510),
            .I(N__10469));
    CascadeMux I__2155 (
            .O(N__10509),
            .I(N__10465));
    LocalMux I__2154 (
            .O(N__10504),
            .I(N__10462));
    InMux I__2153 (
            .O(N__10503),
            .I(N__10453));
    InMux I__2152 (
            .O(N__10502),
            .I(N__10453));
    InMux I__2151 (
            .O(N__10501),
            .I(N__10453));
    InMux I__2150 (
            .O(N__10500),
            .I(N__10453));
    InMux I__2149 (
            .O(N__10499),
            .I(N__10450));
    InMux I__2148 (
            .O(N__10498),
            .I(N__10447));
    InMux I__2147 (
            .O(N__10495),
            .I(N__10440));
    InMux I__2146 (
            .O(N__10492),
            .I(N__10440));
    InMux I__2145 (
            .O(N__10491),
            .I(N__10440));
    InMux I__2144 (
            .O(N__10490),
            .I(N__10437));
    LocalMux I__2143 (
            .O(N__10481),
            .I(N__10434));
    Span4Mux_v I__2142 (
            .O(N__10476),
            .I(N__10431));
    InMux I__2141 (
            .O(N__10475),
            .I(N__10428));
    Span4Mux_h I__2140 (
            .O(N__10472),
            .I(N__10423));
    Span4Mux_h I__2139 (
            .O(N__10469),
            .I(N__10423));
    InMux I__2138 (
            .O(N__10468),
            .I(N__10420));
    InMux I__2137 (
            .O(N__10465),
            .I(N__10417));
    Span4Mux_h I__2136 (
            .O(N__10462),
            .I(N__10412));
    LocalMux I__2135 (
            .O(N__10453),
            .I(N__10412));
    LocalMux I__2134 (
            .O(N__10450),
            .I(\DUT.tx_state_0 ));
    LocalMux I__2133 (
            .O(N__10447),
            .I(\DUT.tx_state_0 ));
    LocalMux I__2132 (
            .O(N__10440),
            .I(\DUT.tx_state_0 ));
    LocalMux I__2131 (
            .O(N__10437),
            .I(\DUT.tx_state_0 ));
    Odrv4 I__2130 (
            .O(N__10434),
            .I(\DUT.tx_state_0 ));
    Odrv4 I__2129 (
            .O(N__10431),
            .I(\DUT.tx_state_0 ));
    LocalMux I__2128 (
            .O(N__10428),
            .I(\DUT.tx_state_0 ));
    Odrv4 I__2127 (
            .O(N__10423),
            .I(\DUT.tx_state_0 ));
    LocalMux I__2126 (
            .O(N__10420),
            .I(\DUT.tx_state_0 ));
    LocalMux I__2125 (
            .O(N__10417),
            .I(\DUT.tx_state_0 ));
    Odrv4 I__2124 (
            .O(N__10412),
            .I(\DUT.tx_state_0 ));
    InMux I__2123 (
            .O(N__10389),
            .I(N__10386));
    LocalMux I__2122 (
            .O(N__10386),
            .I(\DUT.uart_inst0.tx_dataZ0Z_5 ));
    CEMux I__2121 (
            .O(N__10383),
            .I(N__10380));
    LocalMux I__2120 (
            .O(N__10380),
            .I(N__10377));
    Span4Mux_v I__2119 (
            .O(N__10377),
            .I(N__10373));
    CEMux I__2118 (
            .O(N__10376),
            .I(N__10370));
    Sp12to4 I__2117 (
            .O(N__10373),
            .I(N__10365));
    LocalMux I__2116 (
            .O(N__10370),
            .I(N__10365));
    Odrv12 I__2115 (
            .O(N__10365),
            .I(\DUT.uart_inst0.N_71_i ));
    CascadeMux I__2114 (
            .O(N__10362),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_1_1_cascade_ ));
    InMux I__2113 (
            .O(N__10359),
            .I(N__10355));
    InMux I__2112 (
            .O(N__10358),
            .I(N__10352));
    LocalMux I__2111 (
            .O(N__10355),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddr_RNIZ0Z_1 ));
    LocalMux I__2110 (
            .O(N__10352),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddr_RNIZ0Z_1 ));
    InMux I__2109 (
            .O(N__10347),
            .I(N__10341));
    InMux I__2108 (
            .O(N__10346),
            .I(N__10341));
    LocalMux I__2107 (
            .O(N__10341),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddr_0_1 ));
    CascadeMux I__2106 (
            .O(N__10338),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddr_RNIZ0Z_1_cascade_ ));
    CascadeMux I__2105 (
            .O(N__10335),
            .I(N__10332));
    InMux I__2104 (
            .O(N__10332),
            .I(N__10329));
    LocalMux I__2103 (
            .O(N__10329),
            .I(N__10326));
    Span4Mux_h I__2102 (
            .O(N__10326),
            .I(N__10323));
    Odrv4 I__2101 (
            .O(N__10323),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_1 ));
    CascadeMux I__2100 (
            .O(N__10320),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_1_cascade_ ));
    CascadeMux I__2099 (
            .O(N__10317),
            .I(N__10313));
    InMux I__2098 (
            .O(N__10316),
            .I(N__10308));
    InMux I__2097 (
            .O(N__10313),
            .I(N__10308));
    LocalMux I__2096 (
            .O(N__10308),
            .I(\DUT.uart_inst0.tx_dataZ0Z_0 ));
    InMux I__2095 (
            .O(N__10305),
            .I(N__10302));
    LocalMux I__2094 (
            .O(N__10302),
            .I(\DUT.uart_inst0.tx_dataZ0Z_1 ));
    InMux I__2093 (
            .O(N__10299),
            .I(N__10296));
    LocalMux I__2092 (
            .O(N__10296),
            .I(\DUT.uart_inst0.tx_dataZ0Z_3 ));
    InMux I__2091 (
            .O(N__10293),
            .I(N__10290));
    LocalMux I__2090 (
            .O(N__10290),
            .I(\DUT.uart_inst0.tx_dataZ0Z_2 ));
    InMux I__2089 (
            .O(N__10287),
            .I(N__10284));
    LocalMux I__2088 (
            .O(N__10284),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_3 ));
    InMux I__2087 (
            .O(N__10281),
            .I(N__10277));
    InMux I__2086 (
            .O(N__10280),
            .I(N__10274));
    LocalMux I__2085 (
            .O(N__10277),
            .I(N__10268));
    LocalMux I__2084 (
            .O(N__10274),
            .I(N__10268));
    InMux I__2083 (
            .O(N__10273),
            .I(N__10265));
    Span4Mux_h I__2082 (
            .O(N__10268),
            .I(N__10260));
    LocalMux I__2081 (
            .O(N__10265),
            .I(N__10257));
    InMux I__2080 (
            .O(N__10264),
            .I(N__10254));
    InMux I__2079 (
            .O(N__10263),
            .I(N__10251));
    Odrv4 I__2078 (
            .O(N__10260),
            .I(\DUT.wRxByte_4 ));
    Odrv4 I__2077 (
            .O(N__10257),
            .I(\DUT.wRxByte_4 ));
    LocalMux I__2076 (
            .O(N__10254),
            .I(\DUT.wRxByte_4 ));
    LocalMux I__2075 (
            .O(N__10251),
            .I(\DUT.wRxByte_4 ));
    InMux I__2074 (
            .O(N__10242),
            .I(N__10239));
    LocalMux I__2073 (
            .O(N__10239),
            .I(N__10236));
    Odrv4 I__2072 (
            .O(N__10236),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_4 ));
    InMux I__2071 (
            .O(N__10233),
            .I(N__10230));
    LocalMux I__2070 (
            .O(N__10230),
            .I(N__10226));
    InMux I__2069 (
            .O(N__10229),
            .I(N__10223));
    Span4Mux_h I__2068 (
            .O(N__10226),
            .I(N__10217));
    LocalMux I__2067 (
            .O(N__10223),
            .I(N__10214));
    InMux I__2066 (
            .O(N__10222),
            .I(N__10211));
    InMux I__2065 (
            .O(N__10221),
            .I(N__10208));
    InMux I__2064 (
            .O(N__10220),
            .I(N__10205));
    Odrv4 I__2063 (
            .O(N__10217),
            .I(\DUT.wRxByte_5 ));
    Odrv4 I__2062 (
            .O(N__10214),
            .I(\DUT.wRxByte_5 ));
    LocalMux I__2061 (
            .O(N__10211),
            .I(\DUT.wRxByte_5 ));
    LocalMux I__2060 (
            .O(N__10208),
            .I(\DUT.wRxByte_5 ));
    LocalMux I__2059 (
            .O(N__10205),
            .I(\DUT.wRxByte_5 ));
    InMux I__2058 (
            .O(N__10194),
            .I(N__10191));
    LocalMux I__2057 (
            .O(N__10191),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_5 ));
    InMux I__2056 (
            .O(N__10188),
            .I(N__10184));
    InMux I__2055 (
            .O(N__10187),
            .I(N__10180));
    LocalMux I__2054 (
            .O(N__10184),
            .I(N__10177));
    InMux I__2053 (
            .O(N__10183),
            .I(N__10174));
    LocalMux I__2052 (
            .O(N__10180),
            .I(N__10171));
    Span4Mux_h I__2051 (
            .O(N__10177),
            .I(N__10166));
    LocalMux I__2050 (
            .O(N__10174),
            .I(N__10163));
    Span4Mux_h I__2049 (
            .O(N__10171),
            .I(N__10160));
    InMux I__2048 (
            .O(N__10170),
            .I(N__10157));
    InMux I__2047 (
            .O(N__10169),
            .I(N__10154));
    Odrv4 I__2046 (
            .O(N__10166),
            .I(\DUT.wRxByte_6 ));
    Odrv4 I__2045 (
            .O(N__10163),
            .I(\DUT.wRxByte_6 ));
    Odrv4 I__2044 (
            .O(N__10160),
            .I(\DUT.wRxByte_6 ));
    LocalMux I__2043 (
            .O(N__10157),
            .I(\DUT.wRxByte_6 ));
    LocalMux I__2042 (
            .O(N__10154),
            .I(\DUT.wRxByte_6 ));
    InMux I__2041 (
            .O(N__10143),
            .I(N__10140));
    LocalMux I__2040 (
            .O(N__10140),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_6 ));
    InMux I__2039 (
            .O(N__10137),
            .I(N__10133));
    InMux I__2038 (
            .O(N__10136),
            .I(N__10130));
    LocalMux I__2037 (
            .O(N__10133),
            .I(N__10126));
    LocalMux I__2036 (
            .O(N__10130),
            .I(N__10123));
    InMux I__2035 (
            .O(N__10129),
            .I(N__10120));
    Span4Mux_v I__2034 (
            .O(N__10126),
            .I(N__10115));
    Span4Mux_h I__2033 (
            .O(N__10123),
            .I(N__10112));
    LocalMux I__2032 (
            .O(N__10120),
            .I(N__10109));
    InMux I__2031 (
            .O(N__10119),
            .I(N__10106));
    InMux I__2030 (
            .O(N__10118),
            .I(N__10103));
    Odrv4 I__2029 (
            .O(N__10115),
            .I(\DUT.wRxByte_7 ));
    Odrv4 I__2028 (
            .O(N__10112),
            .I(\DUT.wRxByte_7 ));
    Odrv4 I__2027 (
            .O(N__10109),
            .I(\DUT.wRxByte_7 ));
    LocalMux I__2026 (
            .O(N__10106),
            .I(\DUT.wRxByte_7 ));
    LocalMux I__2025 (
            .O(N__10103),
            .I(\DUT.wRxByte_7 ));
    InMux I__2024 (
            .O(N__10092),
            .I(N__10089));
    LocalMux I__2023 (
            .O(N__10089),
            .I(N__10086));
    Odrv4 I__2022 (
            .O(N__10086),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_7 ));
    CEMux I__2021 (
            .O(N__10083),
            .I(N__10079));
    InMux I__2020 (
            .O(N__10082),
            .I(N__10076));
    LocalMux I__2019 (
            .O(N__10079),
            .I(N__10073));
    LocalMux I__2018 (
            .O(N__10076),
            .I(N__10070));
    Span4Mux_h I__2017 (
            .O(N__10073),
            .I(N__10067));
    Span4Mux_h I__2016 (
            .O(N__10070),
            .I(N__10064));
    Odrv4 I__2015 (
            .O(N__10067),
            .I(\DUT.fifo_rx_inst.rFifoData_awe2 ));
    Odrv4 I__2014 (
            .O(N__10064),
            .I(\DUT.fifo_rx_inst.rFifoData_awe2 ));
    InMux I__2013 (
            .O(N__10059),
            .I(N__10055));
    InMux I__2012 (
            .O(N__10058),
            .I(N__10051));
    LocalMux I__2011 (
            .O(N__10055),
            .I(N__10048));
    InMux I__2010 (
            .O(N__10054),
            .I(N__10045));
    LocalMux I__2009 (
            .O(N__10051),
            .I(N__10037));
    Span4Mux_v I__2008 (
            .O(N__10048),
            .I(N__10037));
    LocalMux I__2007 (
            .O(N__10045),
            .I(N__10037));
    InMux I__2006 (
            .O(N__10044),
            .I(N__10034));
    Span4Mux_h I__2005 (
            .O(N__10037),
            .I(N__10031));
    LocalMux I__2004 (
            .O(N__10034),
            .I(N__10028));
    Odrv4 I__2003 (
            .O(N__10031),
            .I(\DUT.wRxByte_0 ));
    Odrv12 I__2002 (
            .O(N__10028),
            .I(\DUT.wRxByte_0 ));
    InMux I__2001 (
            .O(N__10023),
            .I(N__10020));
    LocalMux I__2000 (
            .O(N__10020),
            .I(N__10017));
    Odrv4 I__1999 (
            .O(N__10017),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_0 ));
    CEMux I__1998 (
            .O(N__10014),
            .I(N__10009));
    CEMux I__1997 (
            .O(N__10013),
            .I(N__10006));
    CEMux I__1996 (
            .O(N__10012),
            .I(N__10003));
    LocalMux I__1995 (
            .O(N__10009),
            .I(N__10000));
    LocalMux I__1994 (
            .O(N__10006),
            .I(N__9997));
    LocalMux I__1993 (
            .O(N__10003),
            .I(N__9994));
    Span4Mux_v I__1992 (
            .O(N__10000),
            .I(N__9989));
    Span4Mux_v I__1991 (
            .O(N__9997),
            .I(N__9989));
    Span4Mux_h I__1990 (
            .O(N__9994),
            .I(N__9985));
    Span4Mux_h I__1989 (
            .O(N__9989),
            .I(N__9982));
    InMux I__1988 (
            .O(N__9988),
            .I(N__9979));
    Odrv4 I__1987 (
            .O(N__9985),
            .I(\DUT.fifo_rx_inst.rFifoData_awe0 ));
    Odrv4 I__1986 (
            .O(N__9982),
            .I(\DUT.fifo_rx_inst.rFifoData_awe0 ));
    LocalMux I__1985 (
            .O(N__9979),
            .I(\DUT.fifo_rx_inst.rFifoData_awe0 ));
    InMux I__1984 (
            .O(N__9972),
            .I(N__9969));
    LocalMux I__1983 (
            .O(N__9969),
            .I(\fifo_inst.tx_fifo_inst.rRamRdAddr_0_2 ));
    CascadeMux I__1982 (
            .O(N__9966),
            .I(N__9955));
    CascadeMux I__1981 (
            .O(N__9965),
            .I(N__9950));
    CascadeMux I__1980 (
            .O(N__9964),
            .I(N__9947));
    InMux I__1979 (
            .O(N__9963),
            .I(N__9934));
    InMux I__1978 (
            .O(N__9962),
            .I(N__9934));
    InMux I__1977 (
            .O(N__9961),
            .I(N__9934));
    InMux I__1976 (
            .O(N__9960),
            .I(N__9934));
    InMux I__1975 (
            .O(N__9959),
            .I(N__9934));
    InMux I__1974 (
            .O(N__9958),
            .I(N__9927));
    InMux I__1973 (
            .O(N__9955),
            .I(N__9927));
    InMux I__1972 (
            .O(N__9954),
            .I(N__9927));
    InMux I__1971 (
            .O(N__9953),
            .I(N__9918));
    InMux I__1970 (
            .O(N__9950),
            .I(N__9918));
    InMux I__1969 (
            .O(N__9947),
            .I(N__9918));
    InMux I__1968 (
            .O(N__9946),
            .I(N__9918));
    CascadeMux I__1967 (
            .O(N__9945),
            .I(N__9914));
    LocalMux I__1966 (
            .O(N__9934),
            .I(N__9905));
    LocalMux I__1965 (
            .O(N__9927),
            .I(N__9900));
    LocalMux I__1964 (
            .O(N__9918),
            .I(N__9900));
    InMux I__1963 (
            .O(N__9917),
            .I(N__9895));
    InMux I__1962 (
            .O(N__9914),
            .I(N__9895));
    CascadeMux I__1961 (
            .O(N__9913),
            .I(N__9892));
    InMux I__1960 (
            .O(N__9912),
            .I(N__9887));
    InMux I__1959 (
            .O(N__9911),
            .I(N__9887));
    InMux I__1958 (
            .O(N__9910),
            .I(N__9884));
    InMux I__1957 (
            .O(N__9909),
            .I(N__9879));
    InMux I__1956 (
            .O(N__9908),
            .I(N__9879));
    Span4Mux_h I__1955 (
            .O(N__9905),
            .I(N__9872));
    Span4Mux_v I__1954 (
            .O(N__9900),
            .I(N__9872));
    LocalMux I__1953 (
            .O(N__9895),
            .I(N__9872));
    InMux I__1952 (
            .O(N__9892),
            .I(N__9869));
    LocalMux I__1951 (
            .O(N__9887),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__1950 (
            .O(N__9884),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__1949 (
            .O(N__9879),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    Odrv4 I__1948 (
            .O(N__9872),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__1947 (
            .O(N__9869),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    CascadeMux I__1946 (
            .O(N__9858),
            .I(N__9855));
    InMux I__1945 (
            .O(N__9855),
            .I(N__9852));
    LocalMux I__1944 (
            .O(N__9852),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2 ));
    CEMux I__1943 (
            .O(N__9849),
            .I(N__9846));
    LocalMux I__1942 (
            .O(N__9846),
            .I(N__9842));
    CEMux I__1941 (
            .O(N__9845),
            .I(N__9839));
    Span4Mux_h I__1940 (
            .O(N__9842),
            .I(N__9836));
    LocalMux I__1939 (
            .O(N__9839),
            .I(N__9833));
    Odrv4 I__1938 (
            .O(N__9836),
            .I(N_100_i_0));
    Odrv12 I__1937 (
            .O(N__9833),
            .I(N_100_i_0));
    SRMux I__1936 (
            .O(N__9828),
            .I(N__9824));
    SRMux I__1935 (
            .O(N__9827),
            .I(N__9821));
    LocalMux I__1934 (
            .O(N__9824),
            .I(N__9818));
    LocalMux I__1933 (
            .O(N__9821),
            .I(N__9815));
    Span4Mux_v I__1932 (
            .O(N__9818),
            .I(N__9811));
    Span4Mux_h I__1931 (
            .O(N__9815),
            .I(N__9808));
    InMux I__1930 (
            .O(N__9814),
            .I(N__9805));
    Odrv4 I__1929 (
            .O(N__9811),
            .I(rFifoDatarff_0_RNIHJV05));
    Odrv4 I__1928 (
            .O(N__9808),
            .I(rFifoDatarff_0_RNIHJV05));
    LocalMux I__1927 (
            .O(N__9805),
            .I(rFifoDatarff_0_RNIHJV05));
    InMux I__1926 (
            .O(N__9798),
            .I(N__9795));
    LocalMux I__1925 (
            .O(N__9795),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_1 ));
    InMux I__1924 (
            .O(N__9792),
            .I(N__9789));
    LocalMux I__1923 (
            .O(N__9789),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_0 ));
    InMux I__1922 (
            .O(N__9786),
            .I(N__9783));
    LocalMux I__1921 (
            .O(N__9783),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_2 ));
    InMux I__1920 (
            .O(N__9780),
            .I(N__9777));
    LocalMux I__1919 (
            .O(N__9777),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_4 ));
    InMux I__1918 (
            .O(N__9774),
            .I(N__9769));
    CEMux I__1917 (
            .O(N__9773),
            .I(N__9766));
    CEMux I__1916 (
            .O(N__9772),
            .I(N__9763));
    LocalMux I__1915 (
            .O(N__9769),
            .I(N__9760));
    LocalMux I__1914 (
            .O(N__9766),
            .I(N__9757));
    LocalMux I__1913 (
            .O(N__9763),
            .I(N__9754));
    Span4Mux_v I__1912 (
            .O(N__9760),
            .I(N__9751));
    Span4Mux_v I__1911 (
            .O(N__9757),
            .I(N__9748));
    Span12Mux_h I__1910 (
            .O(N__9754),
            .I(N__9745));
    Span4Mux_h I__1909 (
            .O(N__9751),
            .I(N__9742));
    Odrv4 I__1908 (
            .O(N__9748),
            .I(\DUT.fifo_rx_inst.rFifoData_awe3 ));
    Odrv12 I__1907 (
            .O(N__9745),
            .I(\DUT.fifo_rx_inst.rFifoData_awe3 ));
    Odrv4 I__1906 (
            .O(N__9742),
            .I(\DUT.fifo_rx_inst.rFifoData_awe3 ));
    InMux I__1905 (
            .O(N__9735),
            .I(N__9732));
    LocalMux I__1904 (
            .O(N__9732),
            .I(N__9729));
    Odrv12 I__1903 (
            .O(N__9729),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_0 ));
    InMux I__1902 (
            .O(N__9726),
            .I(N__9722));
    InMux I__1901 (
            .O(N__9725),
            .I(N__9719));
    LocalMux I__1900 (
            .O(N__9722),
            .I(N__9714));
    LocalMux I__1899 (
            .O(N__9719),
            .I(N__9711));
    InMux I__1898 (
            .O(N__9718),
            .I(N__9708));
    InMux I__1897 (
            .O(N__9717),
            .I(N__9705));
    Span4Mux_h I__1896 (
            .O(N__9714),
            .I(N__9701));
    Span4Mux_h I__1895 (
            .O(N__9711),
            .I(N__9698));
    LocalMux I__1894 (
            .O(N__9708),
            .I(N__9695));
    LocalMux I__1893 (
            .O(N__9705),
            .I(N__9692));
    InMux I__1892 (
            .O(N__9704),
            .I(N__9689));
    Odrv4 I__1891 (
            .O(N__9701),
            .I(\DUT.wRxByte_1 ));
    Odrv4 I__1890 (
            .O(N__9698),
            .I(\DUT.wRxByte_1 ));
    Odrv4 I__1889 (
            .O(N__9695),
            .I(\DUT.wRxByte_1 ));
    Odrv4 I__1888 (
            .O(N__9692),
            .I(\DUT.wRxByte_1 ));
    LocalMux I__1887 (
            .O(N__9689),
            .I(\DUT.wRxByte_1 ));
    CascadeMux I__1886 (
            .O(N__9678),
            .I(N__9675));
    InMux I__1885 (
            .O(N__9675),
            .I(N__9672));
    LocalMux I__1884 (
            .O(N__9672),
            .I(N__9669));
    Odrv4 I__1883 (
            .O(N__9669),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_1 ));
    InMux I__1882 (
            .O(N__9666),
            .I(N__9662));
    InMux I__1881 (
            .O(N__9665),
            .I(N__9659));
    LocalMux I__1880 (
            .O(N__9662),
            .I(N__9653));
    LocalMux I__1879 (
            .O(N__9659),
            .I(N__9653));
    InMux I__1878 (
            .O(N__9658),
            .I(N__9650));
    Span4Mux_v I__1877 (
            .O(N__9653),
            .I(N__9645));
    LocalMux I__1876 (
            .O(N__9650),
            .I(N__9642));
    InMux I__1875 (
            .O(N__9649),
            .I(N__9639));
    InMux I__1874 (
            .O(N__9648),
            .I(N__9636));
    Odrv4 I__1873 (
            .O(N__9645),
            .I(\DUT.wRxByte_2 ));
    Odrv4 I__1872 (
            .O(N__9642),
            .I(\DUT.wRxByte_2 ));
    LocalMux I__1871 (
            .O(N__9639),
            .I(\DUT.wRxByte_2 ));
    LocalMux I__1870 (
            .O(N__9636),
            .I(\DUT.wRxByte_2 ));
    InMux I__1869 (
            .O(N__9627),
            .I(N__9624));
    LocalMux I__1868 (
            .O(N__9624),
            .I(N__9621));
    Odrv4 I__1867 (
            .O(N__9621),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_2 ));
    InMux I__1866 (
            .O(N__9618),
            .I(N__9615));
    LocalMux I__1865 (
            .O(N__9615),
            .I(N__9611));
    InMux I__1864 (
            .O(N__9614),
            .I(N__9608));
    Span4Mux_h I__1863 (
            .O(N__9611),
            .I(N__9602));
    LocalMux I__1862 (
            .O(N__9608),
            .I(N__9599));
    InMux I__1861 (
            .O(N__9607),
            .I(N__9596));
    InMux I__1860 (
            .O(N__9606),
            .I(N__9593));
    InMux I__1859 (
            .O(N__9605),
            .I(N__9590));
    Odrv4 I__1858 (
            .O(N__9602),
            .I(\DUT.wRxByte_3 ));
    Odrv4 I__1857 (
            .O(N__9599),
            .I(\DUT.wRxByte_3 ));
    LocalMux I__1856 (
            .O(N__9596),
            .I(\DUT.wRxByte_3 ));
    LocalMux I__1855 (
            .O(N__9593),
            .I(\DUT.wRxByte_3 ));
    LocalMux I__1854 (
            .O(N__9590),
            .I(\DUT.wRxByte_3 ));
    InMux I__1853 (
            .O(N__9579),
            .I(N__9575));
    InMux I__1852 (
            .O(N__9578),
            .I(N__9572));
    LocalMux I__1851 (
            .O(N__9575),
            .I(\DUT.fifo_rx_inst.rFifoDataro_3 ));
    LocalMux I__1850 (
            .O(N__9572),
            .I(\DUT.fifo_rx_inst.rFifoDataro_3 ));
    InMux I__1849 (
            .O(N__9567),
            .I(N__9564));
    LocalMux I__1848 (
            .O(N__9564),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_1 ));
    InMux I__1847 (
            .O(N__9561),
            .I(N__9558));
    LocalMux I__1846 (
            .O(N__9558),
            .I(\fifo_inst.ft2232h_inst.N_103 ));
    InMux I__1845 (
            .O(N__9555),
            .I(N__9551));
    InMux I__1844 (
            .O(N__9554),
            .I(N__9548));
    LocalMux I__1843 (
            .O(N__9551),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_2 ));
    LocalMux I__1842 (
            .O(N__9548),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_2 ));
    InMux I__1841 (
            .O(N__9543),
            .I(N__9539));
    InMux I__1840 (
            .O(N__9542),
            .I(N__9536));
    LocalMux I__1839 (
            .O(N__9539),
            .I(\DUT.fifo_rx_inst.rFifoDataro_2 ));
    LocalMux I__1838 (
            .O(N__9536),
            .I(\DUT.fifo_rx_inst.rFifoDataro_2 ));
    CascadeMux I__1837 (
            .O(N__9531),
            .I(N__9528));
    InMux I__1836 (
            .O(N__9528),
            .I(N__9521));
    InMux I__1835 (
            .O(N__9527),
            .I(N__9516));
    InMux I__1834 (
            .O(N__9526),
            .I(N__9516));
    InMux I__1833 (
            .O(N__9525),
            .I(N__9511));
    InMux I__1832 (
            .O(N__9524),
            .I(N__9511));
    LocalMux I__1831 (
            .O(N__9521),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_0 ));
    LocalMux I__1830 (
            .O(N__9516),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_0 ));
    LocalMux I__1829 (
            .O(N__9511),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_0 ));
    InMux I__1828 (
            .O(N__9504),
            .I(N__9499));
    InMux I__1827 (
            .O(N__9503),
            .I(N__9494));
    InMux I__1826 (
            .O(N__9502),
            .I(N__9494));
    LocalMux I__1825 (
            .O(N__9499),
            .I(N__9491));
    LocalMux I__1824 (
            .O(N__9494),
            .I(N__9488));
    Span4Mux_h I__1823 (
            .O(N__9491),
            .I(N__9485));
    Span4Mux_h I__1822 (
            .O(N__9488),
            .I(N__9482));
    Span4Mux_v I__1821 (
            .O(N__9485),
            .I(N__9479));
    Sp12to4 I__1820 (
            .O(N__9482),
            .I(N__9476));
    Span4Mux_v I__1819 (
            .O(N__9479),
            .I(N__9473));
    Span12Mux_v I__1818 (
            .O(N__9476),
            .I(N__9470));
    Span4Mux_v I__1817 (
            .O(N__9473),
            .I(N__9467));
    Odrv12 I__1816 (
            .O(N__9470),
            .I(iTxE_n_c));
    Odrv4 I__1815 (
            .O(N__9467),
            .I(iTxE_n_c));
    InMux I__1814 (
            .O(N__9462),
            .I(N__9455));
    InMux I__1813 (
            .O(N__9461),
            .I(N__9455));
    InMux I__1812 (
            .O(N__9460),
            .I(N__9450));
    LocalMux I__1811 (
            .O(N__9455),
            .I(N__9447));
    InMux I__1810 (
            .O(N__9454),
            .I(N__9442));
    InMux I__1809 (
            .O(N__9453),
            .I(N__9442));
    LocalMux I__1808 (
            .O(N__9450),
            .I(N__9435));
    Span4Mux_h I__1807 (
            .O(N__9447),
            .I(N__9435));
    LocalMux I__1806 (
            .O(N__9442),
            .I(N__9435));
    Span4Mux_v I__1805 (
            .O(N__9435),
            .I(N__9432));
    Sp12to4 I__1804 (
            .O(N__9432),
            .I(N__9429));
    Span12Mux_h I__1803 (
            .O(N__9429),
            .I(N__9426));
    Odrv12 I__1802 (
            .O(N__9426),
            .I(iRxF_n_c));
    CascadeMux I__1801 (
            .O(N__9423),
            .I(N__9420));
    InMux I__1800 (
            .O(N__9420),
            .I(N__9417));
    LocalMux I__1799 (
            .O(N__9417),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_0 ));
    InMux I__1798 (
            .O(N__9414),
            .I(N__9408));
    InMux I__1797 (
            .O(N__9413),
            .I(N__9401));
    InMux I__1796 (
            .O(N__9412),
            .I(N__9401));
    InMux I__1795 (
            .O(N__9411),
            .I(N__9401));
    LocalMux I__1794 (
            .O(N__9408),
            .I(N__9390));
    LocalMux I__1793 (
            .O(N__9401),
            .I(N__9387));
    InMux I__1792 (
            .O(N__9400),
            .I(N__9382));
    InMux I__1791 (
            .O(N__9399),
            .I(N__9382));
    InMux I__1790 (
            .O(N__9398),
            .I(N__9374));
    InMux I__1789 (
            .O(N__9397),
            .I(N__9374));
    InMux I__1788 (
            .O(N__9396),
            .I(N__9374));
    InMux I__1787 (
            .O(N__9395),
            .I(N__9367));
    InMux I__1786 (
            .O(N__9394),
            .I(N__9367));
    InMux I__1785 (
            .O(N__9393),
            .I(N__9367));
    Span4Mux_h I__1784 (
            .O(N__9390),
            .I(N__9360));
    Span4Mux_v I__1783 (
            .O(N__9387),
            .I(N__9360));
    LocalMux I__1782 (
            .O(N__9382),
            .I(N__9360));
    InMux I__1781 (
            .O(N__9381),
            .I(N__9357));
    LocalMux I__1780 (
            .O(N__9374),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__1779 (
            .O(N__9367),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    Odrv4 I__1778 (
            .O(N__9360),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__1777 (
            .O(N__9357),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    CascadeMux I__1776 (
            .O(N__9348),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ));
    CascadeMux I__1775 (
            .O(N__9345),
            .I(N__9342));
    InMux I__1774 (
            .O(N__9342),
            .I(N__9339));
    LocalMux I__1773 (
            .O(N__9339),
            .I(N__9336));
    Span4Mux_h I__1772 (
            .O(N__9336),
            .I(N__9333));
    Odrv4 I__1771 (
            .O(N__9333),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7 ));
    InMux I__1770 (
            .O(N__9330),
            .I(N__9327));
    LocalMux I__1769 (
            .O(N__9327),
            .I(N__9324));
    Span4Mux_h I__1768 (
            .O(N__9324),
            .I(N__9321));
    Odrv4 I__1767 (
            .O(N__9321),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_7 ));
    InMux I__1766 (
            .O(N__9318),
            .I(N__9315));
    LocalMux I__1765 (
            .O(N__9315),
            .I(N__9312));
    Span4Mux_h I__1764 (
            .O(N__9312),
            .I(N__9309));
    Odrv4 I__1763 (
            .O(N__9309),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1 ));
    InMux I__1762 (
            .O(N__9306),
            .I(N__9303));
    LocalMux I__1761 (
            .O(N__9303),
            .I(N__9292));
    InMux I__1760 (
            .O(N__9302),
            .I(N__9287));
    InMux I__1759 (
            .O(N__9301),
            .I(N__9287));
    InMux I__1758 (
            .O(N__9300),
            .I(N__9282));
    InMux I__1757 (
            .O(N__9299),
            .I(N__9282));
    InMux I__1756 (
            .O(N__9298),
            .I(N__9279));
    InMux I__1755 (
            .O(N__9297),
            .I(N__9274));
    InMux I__1754 (
            .O(N__9296),
            .I(N__9274));
    InMux I__1753 (
            .O(N__9295),
            .I(N__9271));
    Span4Mux_h I__1752 (
            .O(N__9292),
            .I(N__9268));
    LocalMux I__1751 (
            .O(N__9287),
            .I(N__9263));
    LocalMux I__1750 (
            .O(N__9282),
            .I(N__9263));
    LocalMux I__1749 (
            .O(N__9279),
            .I(\DUT.uart_inst0.N_77 ));
    LocalMux I__1748 (
            .O(N__9274),
            .I(\DUT.uart_inst0.N_77 ));
    LocalMux I__1747 (
            .O(N__9271),
            .I(\DUT.uart_inst0.N_77 ));
    Odrv4 I__1746 (
            .O(N__9268),
            .I(\DUT.uart_inst0.N_77 ));
    Odrv4 I__1745 (
            .O(N__9263),
            .I(\DUT.uart_inst0.N_77 ));
    InMux I__1744 (
            .O(N__9252),
            .I(N__9249));
    LocalMux I__1743 (
            .O(N__9249),
            .I(\DUT.uart_inst0.tx_bits_remaining_RNO_0Z0Z_3 ));
    InMux I__1742 (
            .O(N__9246),
            .I(N__9243));
    LocalMux I__1741 (
            .O(N__9243),
            .I(\DUT.uart_inst0.tx_bits_remaining_RNIAIE4LZ0Z_1 ));
    CascadeMux I__1740 (
            .O(N__9240),
            .I(N__9236));
    InMux I__1739 (
            .O(N__9239),
            .I(N__9232));
    InMux I__1738 (
            .O(N__9236),
            .I(N__9229));
    InMux I__1737 (
            .O(N__9235),
            .I(N__9226));
    LocalMux I__1736 (
            .O(N__9232),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_1 ));
    LocalMux I__1735 (
            .O(N__9229),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_1 ));
    LocalMux I__1734 (
            .O(N__9226),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_1 ));
    CascadeMux I__1733 (
            .O(N__9219),
            .I(N__9216));
    InMux I__1732 (
            .O(N__9216),
            .I(N__9213));
    LocalMux I__1731 (
            .O(N__9213),
            .I(N__9207));
    InMux I__1730 (
            .O(N__9212),
            .I(N__9204));
    InMux I__1729 (
            .O(N__9211),
            .I(N__9201));
    InMux I__1728 (
            .O(N__9210),
            .I(N__9198));
    Span4Mux_h I__1727 (
            .O(N__9207),
            .I(N__9195));
    LocalMux I__1726 (
            .O(N__9204),
            .I(N__9192));
    LocalMux I__1725 (
            .O(N__9201),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_0 ));
    LocalMux I__1724 (
            .O(N__9198),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_0 ));
    Odrv4 I__1723 (
            .O(N__9195),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_0 ));
    Odrv4 I__1722 (
            .O(N__9192),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_0 ));
    CascadeMux I__1721 (
            .O(N__9183),
            .I(N__9179));
    InMux I__1720 (
            .O(N__9182),
            .I(N__9174));
    InMux I__1719 (
            .O(N__9179),
            .I(N__9168));
    InMux I__1718 (
            .O(N__9178),
            .I(N__9168));
    InMux I__1717 (
            .O(N__9177),
            .I(N__9165));
    LocalMux I__1716 (
            .O(N__9174),
            .I(N__9162));
    InMux I__1715 (
            .O(N__9173),
            .I(N__9159));
    LocalMux I__1714 (
            .O(N__9168),
            .I(N__9156));
    LocalMux I__1713 (
            .O(N__9165),
            .I(N__9149));
    Span4Mux_h I__1712 (
            .O(N__9162),
            .I(N__9149));
    LocalMux I__1711 (
            .O(N__9159),
            .I(N__9149));
    Odrv12 I__1710 (
            .O(N__9156),
            .I(\DUT.uart_inst0.N_124 ));
    Odrv4 I__1709 (
            .O(N__9149),
            .I(\DUT.uart_inst0.N_124 ));
    CascadeMux I__1708 (
            .O(N__9144),
            .I(N__9141));
    InMux I__1707 (
            .O(N__9141),
            .I(N__9136));
    InMux I__1706 (
            .O(N__9140),
            .I(N__9131));
    InMux I__1705 (
            .O(N__9139),
            .I(N__9131));
    LocalMux I__1704 (
            .O(N__9136),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_2 ));
    LocalMux I__1703 (
            .O(N__9131),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_2 ));
    InMux I__1702 (
            .O(N__9126),
            .I(N__9123));
    LocalMux I__1701 (
            .O(N__9123),
            .I(\DUT.uart_inst0.tx_bits_remaining_RNIBJE4LZ0Z_2 ));
    CascadeMux I__1700 (
            .O(N__9120),
            .I(N__9116));
    InMux I__1699 (
            .O(N__9119),
            .I(N__9111));
    InMux I__1698 (
            .O(N__9116),
            .I(N__9111));
    LocalMux I__1697 (
            .O(N__9111),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_3 ));
    InMux I__1696 (
            .O(N__9108),
            .I(N__9103));
    InMux I__1695 (
            .O(N__9107),
            .I(N__9096));
    InMux I__1694 (
            .O(N__9106),
            .I(N__9093));
    LocalMux I__1693 (
            .O(N__9103),
            .I(N__9090));
    InMux I__1692 (
            .O(N__9102),
            .I(N__9083));
    InMux I__1691 (
            .O(N__9101),
            .I(N__9083));
    InMux I__1690 (
            .O(N__9100),
            .I(N__9083));
    InMux I__1689 (
            .O(N__9099),
            .I(N__9080));
    LocalMux I__1688 (
            .O(N__9096),
            .I(\DUT.uart_inst0.N_96 ));
    LocalMux I__1687 (
            .O(N__9093),
            .I(\DUT.uart_inst0.N_96 ));
    Odrv4 I__1686 (
            .O(N__9090),
            .I(\DUT.uart_inst0.N_96 ));
    LocalMux I__1685 (
            .O(N__9083),
            .I(\DUT.uart_inst0.N_96 ));
    LocalMux I__1684 (
            .O(N__9080),
            .I(\DUT.uart_inst0.N_96 ));
    InMux I__1683 (
            .O(N__9069),
            .I(N__9064));
    InMux I__1682 (
            .O(N__9068),
            .I(N__9061));
    InMux I__1681 (
            .O(N__9067),
            .I(N__9055));
    LocalMux I__1680 (
            .O(N__9064),
            .I(N__9050));
    LocalMux I__1679 (
            .O(N__9061),
            .I(N__9050));
    InMux I__1678 (
            .O(N__9060),
            .I(N__9043));
    InMux I__1677 (
            .O(N__9059),
            .I(N__9043));
    InMux I__1676 (
            .O(N__9058),
            .I(N__9043));
    LocalMux I__1675 (
            .O(N__9055),
            .I(\DUT.uart_inst0.N_99 ));
    Odrv4 I__1674 (
            .O(N__9050),
            .I(\DUT.uart_inst0.N_99 ));
    LocalMux I__1673 (
            .O(N__9043),
            .I(\DUT.uart_inst0.N_99 ));
    InMux I__1672 (
            .O(N__9036),
            .I(N__9033));
    LocalMux I__1671 (
            .O(N__9033),
            .I(\DUT.uart_inst0.un1_tx_bits_remaining_axb_3 ));
    IoInMux I__1670 (
            .O(N__9030),
            .I(N__9026));
    IoInMux I__1669 (
            .O(N__9029),
            .I(N__9023));
    LocalMux I__1668 (
            .O(N__9026),
            .I(N__9020));
    LocalMux I__1667 (
            .O(N__9023),
            .I(N__9017));
    Span4Mux_s0_v I__1666 (
            .O(N__9020),
            .I(N__9014));
    Span4Mux_s2_v I__1665 (
            .O(N__9017),
            .I(N__9011));
    Sp12to4 I__1664 (
            .O(N__9014),
            .I(N__9008));
    Span4Mux_v I__1663 (
            .O(N__9011),
            .I(N__9005));
    Span12Mux_h I__1662 (
            .O(N__9008),
            .I(N__9002));
    Span4Mux_v I__1661 (
            .O(N__9005),
            .I(N__8999));
    Span12Mux_v I__1660 (
            .O(N__9002),
            .I(N__8995));
    Span4Mux_v I__1659 (
            .O(N__8999),
            .I(N__8992));
    InMux I__1658 (
            .O(N__8998),
            .I(N__8989));
    Odrv12 I__1657 (
            .O(N__8995),
            .I(P1A4_c));
    Odrv4 I__1656 (
            .O(N__8992),
            .I(P1A4_c));
    LocalMux I__1655 (
            .O(N__8989),
            .I(P1A4_c));
    CascadeMux I__1654 (
            .O(N__8982),
            .I(\DUT.uart_inst0.tx_countdown_7_i_a3_0_sx_3_cascade_ ));
    InMux I__1653 (
            .O(N__8979),
            .I(N__8976));
    LocalMux I__1652 (
            .O(N__8976),
            .I(\DUT.uart_inst0.N_116 ));
    SRMux I__1651 (
            .O(N__8973),
            .I(N__8969));
    SRMux I__1650 (
            .O(N__8972),
            .I(N__8966));
    LocalMux I__1649 (
            .O(N__8969),
            .I(N__8963));
    LocalMux I__1648 (
            .O(N__8966),
            .I(N__8960));
    Odrv4 I__1647 (
            .O(N__8963),
            .I(\DUT.uart_inst0.N_76_i ));
    Odrv4 I__1646 (
            .O(N__8960),
            .I(\DUT.uart_inst0.N_76_i ));
    CascadeMux I__1645 (
            .O(N__8955),
            .I(N__8947));
    InMux I__1644 (
            .O(N__8954),
            .I(N__8944));
    InMux I__1643 (
            .O(N__8953),
            .I(N__8939));
    InMux I__1642 (
            .O(N__8952),
            .I(N__8939));
    InMux I__1641 (
            .O(N__8951),
            .I(N__8936));
    InMux I__1640 (
            .O(N__8950),
            .I(N__8933));
    InMux I__1639 (
            .O(N__8947),
            .I(N__8930));
    LocalMux I__1638 (
            .O(N__8944),
            .I(N__8927));
    LocalMux I__1637 (
            .O(N__8939),
            .I(N__8924));
    LocalMux I__1636 (
            .O(N__8936),
            .I(N__8921));
    LocalMux I__1635 (
            .O(N__8933),
            .I(\DUT.uart_inst0.tx_countdown_3_2 ));
    LocalMux I__1634 (
            .O(N__8930),
            .I(\DUT.uart_inst0.tx_countdown_3_2 ));
    Odrv4 I__1633 (
            .O(N__8927),
            .I(\DUT.uart_inst0.tx_countdown_3_2 ));
    Odrv4 I__1632 (
            .O(N__8924),
            .I(\DUT.uart_inst0.tx_countdown_3_2 ));
    Odrv4 I__1631 (
            .O(N__8921),
            .I(\DUT.uart_inst0.tx_countdown_3_2 ));
    CascadeMux I__1630 (
            .O(N__8910),
            .I(N__8905));
    InMux I__1629 (
            .O(N__8909),
            .I(N__8900));
    InMux I__1628 (
            .O(N__8908),
            .I(N__8895));
    InMux I__1627 (
            .O(N__8905),
            .I(N__8895));
    InMux I__1626 (
            .O(N__8904),
            .I(N__8891));
    InMux I__1625 (
            .O(N__8903),
            .I(N__8888));
    LocalMux I__1624 (
            .O(N__8900),
            .I(N__8883));
    LocalMux I__1623 (
            .O(N__8895),
            .I(N__8883));
    InMux I__1622 (
            .O(N__8894),
            .I(N__8880));
    LocalMux I__1621 (
            .O(N__8891),
            .I(\DUT.uart_inst0.tx_countdown_3_4 ));
    LocalMux I__1620 (
            .O(N__8888),
            .I(\DUT.uart_inst0.tx_countdown_3_4 ));
    Odrv4 I__1619 (
            .O(N__8883),
            .I(\DUT.uart_inst0.tx_countdown_3_4 ));
    LocalMux I__1618 (
            .O(N__8880),
            .I(\DUT.uart_inst0.tx_countdown_3_4 ));
    InMux I__1617 (
            .O(N__8871),
            .I(N__8863));
    InMux I__1616 (
            .O(N__8870),
            .I(N__8858));
    InMux I__1615 (
            .O(N__8869),
            .I(N__8858));
    CascadeMux I__1614 (
            .O(N__8868),
            .I(N__8855));
    InMux I__1613 (
            .O(N__8867),
            .I(N__8852));
    InMux I__1612 (
            .O(N__8866),
            .I(N__8849));
    LocalMux I__1611 (
            .O(N__8863),
            .I(N__8844));
    LocalMux I__1610 (
            .O(N__8858),
            .I(N__8844));
    InMux I__1609 (
            .O(N__8855),
            .I(N__8841));
    LocalMux I__1608 (
            .O(N__8852),
            .I(\DUT.uart_inst0.tx_countdown_3_1 ));
    LocalMux I__1607 (
            .O(N__8849),
            .I(\DUT.uart_inst0.tx_countdown_3_1 ));
    Odrv4 I__1606 (
            .O(N__8844),
            .I(\DUT.uart_inst0.tx_countdown_3_1 ));
    LocalMux I__1605 (
            .O(N__8841),
            .I(\DUT.uart_inst0.tx_countdown_3_1 ));
    InMux I__1604 (
            .O(N__8832),
            .I(N__8826));
    InMux I__1603 (
            .O(N__8831),
            .I(N__8821));
    InMux I__1602 (
            .O(N__8830),
            .I(N__8821));
    InMux I__1601 (
            .O(N__8829),
            .I(N__8817));
    LocalMux I__1600 (
            .O(N__8826),
            .I(N__8814));
    LocalMux I__1599 (
            .O(N__8821),
            .I(N__8811));
    InMux I__1598 (
            .O(N__8820),
            .I(N__8808));
    LocalMux I__1597 (
            .O(N__8817),
            .I(\DUT.uart_inst0.tx_countdown_3_3 ));
    Odrv4 I__1596 (
            .O(N__8814),
            .I(\DUT.uart_inst0.tx_countdown_3_3 ));
    Odrv4 I__1595 (
            .O(N__8811),
            .I(\DUT.uart_inst0.tx_countdown_3_3 ));
    LocalMux I__1594 (
            .O(N__8808),
            .I(\DUT.uart_inst0.tx_countdown_3_3 ));
    InMux I__1593 (
            .O(N__8799),
            .I(N__8795));
    InMux I__1592 (
            .O(N__8798),
            .I(N__8790));
    LocalMux I__1591 (
            .O(N__8795),
            .I(N__8786));
    InMux I__1590 (
            .O(N__8794),
            .I(N__8781));
    InMux I__1589 (
            .O(N__8793),
            .I(N__8781));
    LocalMux I__1588 (
            .O(N__8790),
            .I(N__8778));
    InMux I__1587 (
            .O(N__8789),
            .I(N__8775));
    Span4Mux_h I__1586 (
            .O(N__8786),
            .I(N__8772));
    LocalMux I__1585 (
            .O(N__8781),
            .I(N__8769));
    Span4Mux_v I__1584 (
            .O(N__8778),
            .I(N__8764));
    LocalMux I__1583 (
            .O(N__8775),
            .I(N__8764));
    Odrv4 I__1582 (
            .O(N__8772),
            .I(\DUT.uart_inst0.tx_countdown_3_0 ));
    Odrv4 I__1581 (
            .O(N__8769),
            .I(\DUT.uart_inst0.tx_countdown_3_0 ));
    Odrv4 I__1580 (
            .O(N__8764),
            .I(\DUT.uart_inst0.tx_countdown_3_0 ));
    CascadeMux I__1579 (
            .O(N__8757),
            .I(\DUT.uart_inst0.N_77_cascade_ ));
    CascadeMux I__1578 (
            .O(N__8754),
            .I(N__8750));
    InMux I__1577 (
            .O(N__8753),
            .I(N__8744));
    InMux I__1576 (
            .O(N__8750),
            .I(N__8739));
    InMux I__1575 (
            .O(N__8749),
            .I(N__8739));
    InMux I__1574 (
            .O(N__8748),
            .I(N__8735));
    InMux I__1573 (
            .O(N__8747),
            .I(N__8732));
    LocalMux I__1572 (
            .O(N__8744),
            .I(N__8729));
    LocalMux I__1571 (
            .O(N__8739),
            .I(N__8726));
    InMux I__1570 (
            .O(N__8738),
            .I(N__8723));
    LocalMux I__1569 (
            .O(N__8735),
            .I(\DUT.uart_inst0.tx_countdown_3_5 ));
    LocalMux I__1568 (
            .O(N__8732),
            .I(\DUT.uart_inst0.tx_countdown_3_5 ));
    Odrv4 I__1567 (
            .O(N__8729),
            .I(\DUT.uart_inst0.tx_countdown_3_5 ));
    Odrv4 I__1566 (
            .O(N__8726),
            .I(\DUT.uart_inst0.tx_countdown_3_5 ));
    LocalMux I__1565 (
            .O(N__8723),
            .I(\DUT.uart_inst0.tx_countdown_3_5 ));
    CascadeMux I__1564 (
            .O(N__8712),
            .I(\DUT.uart_inst0.tx_state_RNI9DTT5Z0Z_0_cascade_ ));
    InMux I__1563 (
            .O(N__8709),
            .I(N__8706));
    LocalMux I__1562 (
            .O(N__8706),
            .I(\DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIMJ5ECZ0 ));
    CascadeMux I__1561 (
            .O(N__8703),
            .I(\DUT.uart_inst0.N_99_cascade_ ));
    InMux I__1560 (
            .O(N__8700),
            .I(N__8697));
    LocalMux I__1559 (
            .O(N__8697),
            .I(\DUT.uart_inst0.un1_tx_bits_remaining_cry_0_c_RNOZ0 ));
    InMux I__1558 (
            .O(N__8694),
            .I(N__8683));
    InMux I__1557 (
            .O(N__8693),
            .I(N__8683));
    InMux I__1556 (
            .O(N__8692),
            .I(N__8680));
    InMux I__1555 (
            .O(N__8691),
            .I(N__8675));
    InMux I__1554 (
            .O(N__8690),
            .I(N__8675));
    InMux I__1553 (
            .O(N__8689),
            .I(N__8670));
    InMux I__1552 (
            .O(N__8688),
            .I(N__8670));
    LocalMux I__1551 (
            .O(N__8683),
            .I(N__8667));
    LocalMux I__1550 (
            .O(N__8680),
            .I(\DUT.tx_state_1 ));
    LocalMux I__1549 (
            .O(N__8675),
            .I(\DUT.tx_state_1 ));
    LocalMux I__1548 (
            .O(N__8670),
            .I(\DUT.tx_state_1 ));
    Odrv4 I__1547 (
            .O(N__8667),
            .I(\DUT.tx_state_1 ));
    CascadeMux I__1546 (
            .O(N__8658),
            .I(N__8655));
    InMux I__1545 (
            .O(N__8655),
            .I(N__8652));
    LocalMux I__1544 (
            .O(N__8652),
            .I(N__8649));
    Span4Mux_v I__1543 (
            .O(N__8649),
            .I(N__8646));
    Odrv4 I__1542 (
            .O(N__8646),
            .I(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_3 ));
    CascadeMux I__1541 (
            .O(N__8643),
            .I(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_3_cascade_ ));
    IoInMux I__1540 (
            .O(N__8640),
            .I(N__8637));
    LocalMux I__1539 (
            .O(N__8637),
            .I(N__8634));
    Span4Mux_s2_v I__1538 (
            .O(N__8634),
            .I(N__8631));
    Span4Mux_v I__1537 (
            .O(N__8631),
            .I(N__8628));
    Span4Mux_v I__1536 (
            .O(N__8628),
            .I(N__8624));
    CascadeMux I__1535 (
            .O(N__8627),
            .I(N__8621));
    Span4Mux_h I__1534 (
            .O(N__8624),
            .I(N__8617));
    InMux I__1533 (
            .O(N__8621),
            .I(N__8614));
    InMux I__1532 (
            .O(N__8620),
            .I(N__8611));
    Odrv4 I__1531 (
            .O(N__8617),
            .I(P1A7_c));
    LocalMux I__1530 (
            .O(N__8614),
            .I(P1A7_c));
    LocalMux I__1529 (
            .O(N__8611),
            .I(P1A7_c));
    InMux I__1528 (
            .O(N__8604),
            .I(N__8601));
    LocalMux I__1527 (
            .O(N__8601),
            .I(\DUT.uart_inst0.N_112 ));
    CascadeMux I__1526 (
            .O(N__8598),
            .I(\DUT.uart_inst0.tx_out_6_iv_0_a3_1_1_cascade_ ));
    CascadeMux I__1525 (
            .O(N__8595),
            .I(\DUT.uart_inst0.tx_out_6_iv_0_a3_1_sx_cascade_ ));
    InMux I__1524 (
            .O(N__8592),
            .I(N__8589));
    LocalMux I__1523 (
            .O(N__8589),
            .I(\DUT.uart_inst0.N_113 ));
    CascadeMux I__1522 (
            .O(N__8586),
            .I(N__8583));
    InMux I__1521 (
            .O(N__8583),
            .I(N__8580));
    LocalMux I__1520 (
            .O(N__8580),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_3 ));
    InMux I__1519 (
            .O(N__8577),
            .I(N__8574));
    LocalMux I__1518 (
            .O(N__8574),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_3 ));
    CascadeMux I__1517 (
            .O(N__8571),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ));
    InMux I__1516 (
            .O(N__8568),
            .I(N__8565));
    LocalMux I__1515 (
            .O(N__8565),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6 ));
    InMux I__1514 (
            .O(N__8562),
            .I(N__8559));
    LocalMux I__1513 (
            .O(N__8559),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_6 ));
    InMux I__1512 (
            .O(N__8556),
            .I(N__8553));
    LocalMux I__1511 (
            .O(N__8553),
            .I(N__8550));
    Odrv12 I__1510 (
            .O(N__8550),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_3 ));
    InMux I__1509 (
            .O(N__8547),
            .I(N__8544));
    LocalMux I__1508 (
            .O(N__8544),
            .I(N__8541));
    Odrv4 I__1507 (
            .O(N__8541),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_5 ));
    CascadeMux I__1506 (
            .O(N__8538),
            .I(N__8528));
    CascadeMux I__1505 (
            .O(N__8537),
            .I(N__8525));
    CascadeMux I__1504 (
            .O(N__8536),
            .I(N__8521));
    CascadeMux I__1503 (
            .O(N__8535),
            .I(N__8517));
    CascadeMux I__1502 (
            .O(N__8534),
            .I(N__8513));
    CascadeMux I__1501 (
            .O(N__8533),
            .I(N__8509));
    CascadeMux I__1500 (
            .O(N__8532),
            .I(N__8505));
    InMux I__1499 (
            .O(N__8531),
            .I(N__8484));
    InMux I__1498 (
            .O(N__8528),
            .I(N__8484));
    InMux I__1497 (
            .O(N__8525),
            .I(N__8484));
    InMux I__1496 (
            .O(N__8524),
            .I(N__8484));
    InMux I__1495 (
            .O(N__8521),
            .I(N__8484));
    InMux I__1494 (
            .O(N__8520),
            .I(N__8484));
    InMux I__1493 (
            .O(N__8517),
            .I(N__8469));
    InMux I__1492 (
            .O(N__8516),
            .I(N__8469));
    InMux I__1491 (
            .O(N__8513),
            .I(N__8469));
    InMux I__1490 (
            .O(N__8512),
            .I(N__8469));
    InMux I__1489 (
            .O(N__8509),
            .I(N__8469));
    InMux I__1488 (
            .O(N__8508),
            .I(N__8469));
    InMux I__1487 (
            .O(N__8505),
            .I(N__8469));
    CascadeMux I__1486 (
            .O(N__8504),
            .I(N__8464));
    CascadeMux I__1485 (
            .O(N__8503),
            .I(N__8460));
    CascadeMux I__1484 (
            .O(N__8502),
            .I(N__8456));
    CascadeMux I__1483 (
            .O(N__8501),
            .I(N__8452));
    CascadeMux I__1482 (
            .O(N__8500),
            .I(N__8447));
    CascadeMux I__1481 (
            .O(N__8499),
            .I(N__8444));
    CascadeMux I__1480 (
            .O(N__8498),
            .I(N__8441));
    CascadeMux I__1479 (
            .O(N__8497),
            .I(N__8436));
    LocalMux I__1478 (
            .O(N__8484),
            .I(N__8430));
    LocalMux I__1477 (
            .O(N__8469),
            .I(N__8430));
    InMux I__1476 (
            .O(N__8468),
            .I(N__8427));
    InMux I__1475 (
            .O(N__8467),
            .I(N__8410));
    InMux I__1474 (
            .O(N__8464),
            .I(N__8410));
    InMux I__1473 (
            .O(N__8463),
            .I(N__8410));
    InMux I__1472 (
            .O(N__8460),
            .I(N__8410));
    InMux I__1471 (
            .O(N__8459),
            .I(N__8410));
    InMux I__1470 (
            .O(N__8456),
            .I(N__8410));
    InMux I__1469 (
            .O(N__8455),
            .I(N__8410));
    InMux I__1468 (
            .O(N__8452),
            .I(N__8410));
    InMux I__1467 (
            .O(N__8451),
            .I(N__8407));
    InMux I__1466 (
            .O(N__8450),
            .I(N__8392));
    InMux I__1465 (
            .O(N__8447),
            .I(N__8392));
    InMux I__1464 (
            .O(N__8444),
            .I(N__8392));
    InMux I__1463 (
            .O(N__8441),
            .I(N__8392));
    InMux I__1462 (
            .O(N__8440),
            .I(N__8392));
    InMux I__1461 (
            .O(N__8439),
            .I(N__8392));
    InMux I__1460 (
            .O(N__8436),
            .I(N__8392));
    InMux I__1459 (
            .O(N__8435),
            .I(N__8389));
    Span4Mux_v I__1458 (
            .O(N__8430),
            .I(N__8381));
    LocalMux I__1457 (
            .O(N__8427),
            .I(N__8381));
    LocalMux I__1456 (
            .O(N__8410),
            .I(N__8381));
    LocalMux I__1455 (
            .O(N__8407),
            .I(N__8376));
    LocalMux I__1454 (
            .O(N__8392),
            .I(N__8376));
    LocalMux I__1453 (
            .O(N__8389),
            .I(N__8373));
    InMux I__1452 (
            .O(N__8388),
            .I(N__8370));
    Span4Mux_v I__1451 (
            .O(N__8381),
            .I(N__8365));
    Span4Mux_v I__1450 (
            .O(N__8376),
            .I(N__8365));
    Span4Mux_v I__1449 (
            .O(N__8373),
            .I(N__8362));
    LocalMux I__1448 (
            .O(N__8370),
            .I(N__8359));
    Odrv4 I__1447 (
            .O(N__8365),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1446 (
            .O(N__8362),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__1445 (
            .O(N__8359),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__1444 (
            .O(N__8352),
            .I(N__8345));
    CascadeMux I__1443 (
            .O(N__8351),
            .I(N__8342));
    InMux I__1442 (
            .O(N__8350),
            .I(N__8337));
    CascadeMux I__1441 (
            .O(N__8349),
            .I(N__8330));
    InMux I__1440 (
            .O(N__8348),
            .I(N__8322));
    InMux I__1439 (
            .O(N__8345),
            .I(N__8322));
    InMux I__1438 (
            .O(N__8342),
            .I(N__8322));
    CascadeMux I__1437 (
            .O(N__8341),
            .I(N__8312));
    InMux I__1436 (
            .O(N__8340),
            .I(N__8309));
    LocalMux I__1435 (
            .O(N__8337),
            .I(N__8306));
    InMux I__1434 (
            .O(N__8336),
            .I(N__8303));
    InMux I__1433 (
            .O(N__8335),
            .I(N__8298));
    InMux I__1432 (
            .O(N__8334),
            .I(N__8293));
    InMux I__1431 (
            .O(N__8333),
            .I(N__8293));
    InMux I__1430 (
            .O(N__8330),
            .I(N__8288));
    InMux I__1429 (
            .O(N__8329),
            .I(N__8288));
    LocalMux I__1428 (
            .O(N__8322),
            .I(N__8275));
    InMux I__1427 (
            .O(N__8321),
            .I(N__8270));
    InMux I__1426 (
            .O(N__8320),
            .I(N__8270));
    InMux I__1425 (
            .O(N__8319),
            .I(N__8265));
    InMux I__1424 (
            .O(N__8318),
            .I(N__8265));
    InMux I__1423 (
            .O(N__8317),
            .I(N__8256));
    InMux I__1422 (
            .O(N__8316),
            .I(N__8256));
    InMux I__1421 (
            .O(N__8315),
            .I(N__8256));
    InMux I__1420 (
            .O(N__8312),
            .I(N__8256));
    LocalMux I__1419 (
            .O(N__8309),
            .I(N__8253));
    Span4Mux_v I__1418 (
            .O(N__8306),
            .I(N__8248));
    LocalMux I__1417 (
            .O(N__8303),
            .I(N__8248));
    InMux I__1416 (
            .O(N__8302),
            .I(N__8245));
    InMux I__1415 (
            .O(N__8301),
            .I(N__8242));
    LocalMux I__1414 (
            .O(N__8298),
            .I(N__8235));
    LocalMux I__1413 (
            .O(N__8293),
            .I(N__8235));
    LocalMux I__1412 (
            .O(N__8288),
            .I(N__8235));
    InMux I__1411 (
            .O(N__8287),
            .I(N__8220));
    InMux I__1410 (
            .O(N__8286),
            .I(N__8220));
    InMux I__1409 (
            .O(N__8285),
            .I(N__8220));
    InMux I__1408 (
            .O(N__8284),
            .I(N__8220));
    InMux I__1407 (
            .O(N__8283),
            .I(N__8220));
    InMux I__1406 (
            .O(N__8282),
            .I(N__8220));
    InMux I__1405 (
            .O(N__8281),
            .I(N__8220));
    InMux I__1404 (
            .O(N__8280),
            .I(N__8217));
    InMux I__1403 (
            .O(N__8279),
            .I(N__8212));
    InMux I__1402 (
            .O(N__8278),
            .I(N__8212));
    Span4Mux_v I__1401 (
            .O(N__8275),
            .I(N__8207));
    LocalMux I__1400 (
            .O(N__8270),
            .I(N__8207));
    LocalMux I__1399 (
            .O(N__8265),
            .I(N__8202));
    LocalMux I__1398 (
            .O(N__8256),
            .I(N__8202));
    Span4Mux_v I__1397 (
            .O(N__8253),
            .I(N__8199));
    Span4Mux_v I__1396 (
            .O(N__8248),
            .I(N__8194));
    LocalMux I__1395 (
            .O(N__8245),
            .I(N__8194));
    LocalMux I__1394 (
            .O(N__8242),
            .I(N__8183));
    Span4Mux_v I__1393 (
            .O(N__8235),
            .I(N__8183));
    LocalMux I__1392 (
            .O(N__8220),
            .I(N__8183));
    LocalMux I__1391 (
            .O(N__8217),
            .I(N__8183));
    LocalMux I__1390 (
            .O(N__8212),
            .I(N__8183));
    Span4Mux_v I__1389 (
            .O(N__8207),
            .I(N__8178));
    Span4Mux_v I__1388 (
            .O(N__8202),
            .I(N__8178));
    Span4Mux_h I__1387 (
            .O(N__8199),
            .I(N__8171));
    Span4Mux_v I__1386 (
            .O(N__8194),
            .I(N__8171));
    Span4Mux_v I__1385 (
            .O(N__8183),
            .I(N__8171));
    Sp12to4 I__1384 (
            .O(N__8178),
            .I(N__8166));
    Sp12to4 I__1383 (
            .O(N__8171),
            .I(N__8166));
    Span12Mux_h I__1382 (
            .O(N__8166),
            .I(N__8163));
    Odrv12 I__1381 (
            .O(N__8163),
            .I(P1A1_c));
    InMux I__1380 (
            .O(N__8160),
            .I(N__8157));
    LocalMux I__1379 (
            .O(N__8157),
            .I(N__8154));
    Span4Mux_h I__1378 (
            .O(N__8154),
            .I(N__8151));
    Odrv4 I__1377 (
            .O(N__8151),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO ));
    CascadeMux I__1376 (
            .O(N__8148),
            .I(N__8141));
    CascadeMux I__1375 (
            .O(N__8147),
            .I(N__8134));
    CascadeMux I__1374 (
            .O(N__8146),
            .I(N__8131));
    CascadeMux I__1373 (
            .O(N__8145),
            .I(N__8128));
    CascadeMux I__1372 (
            .O(N__8144),
            .I(N__8125));
    InMux I__1371 (
            .O(N__8141),
            .I(N__8116));
    CascadeMux I__1370 (
            .O(N__8140),
            .I(N__8111));
    InMux I__1369 (
            .O(N__8139),
            .I(N__8096));
    InMux I__1368 (
            .O(N__8138),
            .I(N__8096));
    InMux I__1367 (
            .O(N__8137),
            .I(N__8096));
    InMux I__1366 (
            .O(N__8134),
            .I(N__8096));
    InMux I__1365 (
            .O(N__8131),
            .I(N__8096));
    InMux I__1364 (
            .O(N__8128),
            .I(N__8096));
    InMux I__1363 (
            .O(N__8125),
            .I(N__8096));
    InMux I__1362 (
            .O(N__8124),
            .I(N__8091));
    InMux I__1361 (
            .O(N__8123),
            .I(N__8091));
    CascadeMux I__1360 (
            .O(N__8122),
            .I(N__8088));
    CascadeMux I__1359 (
            .O(N__8121),
            .I(N__8085));
    CascadeMux I__1358 (
            .O(N__8120),
            .I(N__8082));
    CascadeMux I__1357 (
            .O(N__8119),
            .I(N__8079));
    LocalMux I__1356 (
            .O(N__8116),
            .I(N__8074));
    InMux I__1355 (
            .O(N__8115),
            .I(N__8071));
    InMux I__1354 (
            .O(N__8114),
            .I(N__8065));
    InMux I__1353 (
            .O(N__8111),
            .I(N__8065));
    LocalMux I__1352 (
            .O(N__8096),
            .I(N__8060));
    LocalMux I__1351 (
            .O(N__8091),
            .I(N__8060));
    InMux I__1350 (
            .O(N__8088),
            .I(N__8047));
    InMux I__1349 (
            .O(N__8085),
            .I(N__8047));
    InMux I__1348 (
            .O(N__8082),
            .I(N__8047));
    InMux I__1347 (
            .O(N__8079),
            .I(N__8047));
    InMux I__1346 (
            .O(N__8078),
            .I(N__8047));
    InMux I__1345 (
            .O(N__8077),
            .I(N__8047));
    Span4Mux_v I__1344 (
            .O(N__8074),
            .I(N__8042));
    LocalMux I__1343 (
            .O(N__8071),
            .I(N__8042));
    InMux I__1342 (
            .O(N__8070),
            .I(N__8037));
    LocalMux I__1341 (
            .O(N__8065),
            .I(N__8034));
    Span4Mux_v I__1340 (
            .O(N__8060),
            .I(N__8031));
    LocalMux I__1339 (
            .O(N__8047),
            .I(N__8026));
    Span4Mux_h I__1338 (
            .O(N__8042),
            .I(N__8026));
    InMux I__1337 (
            .O(N__8041),
            .I(N__8021));
    InMux I__1336 (
            .O(N__8040),
            .I(N__8021));
    LocalMux I__1335 (
            .O(N__8037),
            .I(\DUT.uart_inst0.recv_stateZ0Z_0 ));
    Odrv12 I__1334 (
            .O(N__8034),
            .I(\DUT.uart_inst0.recv_stateZ0Z_0 ));
    Odrv4 I__1333 (
            .O(N__8031),
            .I(\DUT.uart_inst0.recv_stateZ0Z_0 ));
    Odrv4 I__1332 (
            .O(N__8026),
            .I(\DUT.uart_inst0.recv_stateZ0Z_0 ));
    LocalMux I__1331 (
            .O(N__8021),
            .I(\DUT.uart_inst0.recv_stateZ0Z_0 ));
    CascadeMux I__1330 (
            .O(N__8010),
            .I(N__8006));
    CascadeMux I__1329 (
            .O(N__8009),
            .I(N__8003));
    InMux I__1328 (
            .O(N__8006),
            .I(N__7999));
    InMux I__1327 (
            .O(N__8003),
            .I(N__7996));
    InMux I__1326 (
            .O(N__8002),
            .I(N__7993));
    LocalMux I__1325 (
            .O(N__7999),
            .I(N__7988));
    LocalMux I__1324 (
            .O(N__7996),
            .I(N__7988));
    LocalMux I__1323 (
            .O(N__7993),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_4 ));
    Odrv12 I__1322 (
            .O(N__7988),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_4 ));
    CascadeMux I__1321 (
            .O(N__7983),
            .I(N__7980));
    InMux I__1320 (
            .O(N__7980),
            .I(N__7977));
    LocalMux I__1319 (
            .O(N__7977),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_6 ));
    CascadeMux I__1318 (
            .O(N__7974),
            .I(N__7971));
    InMux I__1317 (
            .O(N__7971),
            .I(N__7968));
    LocalMux I__1316 (
            .O(N__7968),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_7 ));
    CEMux I__1315 (
            .O(N__7965),
            .I(N__7962));
    LocalMux I__1314 (
            .O(N__7962),
            .I(N__7959));
    Span4Mux_h I__1313 (
            .O(N__7959),
            .I(N__7955));
    InMux I__1312 (
            .O(N__7958),
            .I(N__7952));
    Odrv4 I__1311 (
            .O(N__7955),
            .I(\DUT.fifo_rx_inst.rFifoData_awe1 ));
    LocalMux I__1310 (
            .O(N__7952),
            .I(\DUT.fifo_rx_inst.rFifoData_awe1 ));
    InMux I__1309 (
            .O(N__7947),
            .I(N__7944));
    LocalMux I__1308 (
            .O(N__7944),
            .I(N__7941));
    Odrv4 I__1307 (
            .O(N__7941),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_4 ));
    InMux I__1306 (
            .O(N__7938),
            .I(N__7935));
    LocalMux I__1305 (
            .O(N__7935),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_4 ));
    CascadeMux I__1304 (
            .O(N__7932),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4_cascade_ ));
    InMux I__1303 (
            .O(N__7929),
            .I(N__7926));
    LocalMux I__1302 (
            .O(N__7926),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_5 ));
    CascadeMux I__1301 (
            .O(N__7923),
            .I(N__7920));
    InMux I__1300 (
            .O(N__7920),
            .I(N__7917));
    LocalMux I__1299 (
            .O(N__7917),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_5 ));
    InMux I__1298 (
            .O(N__7914),
            .I(N__7911));
    LocalMux I__1297 (
            .O(N__7911),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5 ));
    InMux I__1296 (
            .O(N__7908),
            .I(N__7905));
    LocalMux I__1295 (
            .O(N__7905),
            .I(N_100_i));
    InMux I__1294 (
            .O(N__7902),
            .I(N__7899));
    LocalMux I__1293 (
            .O(N__7899),
            .I(\DUT.fifo_rx_inst.rTxByte_52_1 ));
    CascadeMux I__1292 (
            .O(N__7896),
            .I(\DUT.fifo_rx_inst.rTxByte_52_0_cascade_ ));
    InMux I__1291 (
            .O(N__7893),
            .I(N__7886));
    InMux I__1290 (
            .O(N__7892),
            .I(N__7886));
    InMux I__1289 (
            .O(N__7891),
            .I(N__7883));
    LocalMux I__1288 (
            .O(N__7886),
            .I(N__7880));
    LocalMux I__1287 (
            .O(N__7883),
            .I(N__7875));
    Span4Mux_v I__1286 (
            .O(N__7880),
            .I(N__7875));
    Odrv4 I__1285 (
            .O(N__7875),
            .I(\DUT.fifo_rx_inst.rFifoCount_RNIHH0D1Z0Z_0 ));
    CascadeMux I__1284 (
            .O(N__7872),
            .I(N__7869));
    InMux I__1283 (
            .O(N__7869),
            .I(N__7866));
    LocalMux I__1282 (
            .O(N__7866),
            .I(N__7863));
    Odrv4 I__1281 (
            .O(N__7863),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_2 ));
    CascadeMux I__1280 (
            .O(N__7860),
            .I(N__7857));
    InMux I__1279 (
            .O(N__7857),
            .I(N__7854));
    LocalMux I__1278 (
            .O(N__7854),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_1 ));
    InMux I__1277 (
            .O(N__7851),
            .I(N__7848));
    LocalMux I__1276 (
            .O(N__7848),
            .I(N__7845));
    Odrv4 I__1275 (
            .O(N__7845),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_2 ));
    InMux I__1274 (
            .O(N__7842),
            .I(N__7839));
    LocalMux I__1273 (
            .O(N__7839),
            .I(\DUT.uart_inst0.tx_countdown_3_axb_5 ));
    InMux I__1272 (
            .O(N__7836),
            .I(\DUT.uart_inst0.tx_countdown_3_cry_4 ));
    CascadeMux I__1271 (
            .O(N__7833),
            .I(N__7829));
    CascadeMux I__1270 (
            .O(N__7832),
            .I(N__7826));
    InMux I__1269 (
            .O(N__7829),
            .I(N__7823));
    InMux I__1268 (
            .O(N__7826),
            .I(N__7820));
    LocalMux I__1267 (
            .O(N__7823),
            .I(N__7817));
    LocalMux I__1266 (
            .O(N__7820),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_1 ));
    Odrv4 I__1265 (
            .O(N__7817),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_1 ));
    InMux I__1264 (
            .O(N__7812),
            .I(N__7809));
    LocalMux I__1263 (
            .O(N__7809),
            .I(\DUT.uart_inst0.tx_countdown_RNI4K692Z0Z_1 ));
    InMux I__1262 (
            .O(N__7806),
            .I(N__7795));
    InMux I__1261 (
            .O(N__7805),
            .I(N__7795));
    InMux I__1260 (
            .O(N__7804),
            .I(N__7790));
    InMux I__1259 (
            .O(N__7803),
            .I(N__7790));
    InMux I__1258 (
            .O(N__7802),
            .I(N__7783));
    InMux I__1257 (
            .O(N__7801),
            .I(N__7783));
    InMux I__1256 (
            .O(N__7800),
            .I(N__7783));
    LocalMux I__1255 (
            .O(N__7795),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_10 ));
    LocalMux I__1254 (
            .O(N__7790),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_10 ));
    LocalMux I__1253 (
            .O(N__7783),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_10 ));
    CascadeMux I__1252 (
            .O(N__7776),
            .I(N__7772));
    InMux I__1251 (
            .O(N__7775),
            .I(N__7769));
    InMux I__1250 (
            .O(N__7772),
            .I(N__7766));
    LocalMux I__1249 (
            .O(N__7769),
            .I(\DUT.uart_inst0.tx_countdownZ1Z_3 ));
    LocalMux I__1248 (
            .O(N__7766),
            .I(\DUT.uart_inst0.tx_countdownZ1Z_3 ));
    InMux I__1247 (
            .O(N__7761),
            .I(N__7756));
    CascadeMux I__1246 (
            .O(N__7760),
            .I(N__7752));
    CascadeMux I__1245 (
            .O(N__7759),
            .I(N__7748));
    LocalMux I__1244 (
            .O(N__7756),
            .I(N__7743));
    InMux I__1243 (
            .O(N__7755),
            .I(N__7740));
    InMux I__1242 (
            .O(N__7752),
            .I(N__7735));
    InMux I__1241 (
            .O(N__7751),
            .I(N__7735));
    InMux I__1240 (
            .O(N__7748),
            .I(N__7728));
    InMux I__1239 (
            .O(N__7747),
            .I(N__7728));
    InMux I__1238 (
            .O(N__7746),
            .I(N__7728));
    Odrv12 I__1237 (
            .O(N__7743),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_8 ));
    LocalMux I__1236 (
            .O(N__7740),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_8 ));
    LocalMux I__1235 (
            .O(N__7735),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_8 ));
    LocalMux I__1234 (
            .O(N__7728),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_8 ));
    InMux I__1233 (
            .O(N__7719),
            .I(N__7710));
    InMux I__1232 (
            .O(N__7718),
            .I(N__7705));
    InMux I__1231 (
            .O(N__7717),
            .I(N__7705));
    InMux I__1230 (
            .O(N__7716),
            .I(N__7696));
    InMux I__1229 (
            .O(N__7715),
            .I(N__7696));
    InMux I__1228 (
            .O(N__7714),
            .I(N__7696));
    InMux I__1227 (
            .O(N__7713),
            .I(N__7696));
    LocalMux I__1226 (
            .O(N__7710),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_9 ));
    LocalMux I__1225 (
            .O(N__7705),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_9 ));
    LocalMux I__1224 (
            .O(N__7696),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_9 ));
    InMux I__1223 (
            .O(N__7689),
            .I(N__7686));
    LocalMux I__1222 (
            .O(N__7686),
            .I(\DUT.uart_inst0.tx_countdown_RNI6M692Z0Z_3 ));
    InMux I__1221 (
            .O(N__7683),
            .I(\DUT.uart_inst0.un1_tx_bits_remaining_cry_0 ));
    InMux I__1220 (
            .O(N__7680),
            .I(\DUT.uart_inst0.un1_tx_bits_remaining_cry_1 ));
    InMux I__1219 (
            .O(N__7677),
            .I(\DUT.uart_inst0.un1_tx_bits_remaining_cry_2 ));
    IoInMux I__1218 (
            .O(N__7674),
            .I(N__7671));
    LocalMux I__1217 (
            .O(N__7671),
            .I(N__7668));
    IoSpan4Mux I__1216 (
            .O(N__7668),
            .I(N__7664));
    IoInMux I__1215 (
            .O(N__7667),
            .I(N__7661));
    Span4Mux_s3_v I__1214 (
            .O(N__7664),
            .I(N__7658));
    LocalMux I__1213 (
            .O(N__7661),
            .I(N__7655));
    Span4Mux_h I__1212 (
            .O(N__7658),
            .I(N__7650));
    Span4Mux_s3_v I__1211 (
            .O(N__7655),
            .I(N__7650));
    Sp12to4 I__1210 (
            .O(N__7650),
            .I(N__7647));
    Span12Mux_s11_h I__1209 (
            .O(N__7647),
            .I(N__7643));
    InMux I__1208 (
            .O(N__7646),
            .I(N__7640));
    Odrv12 I__1207 (
            .O(N__7643),
            .I(P1A3_c));
    LocalMux I__1206 (
            .O(N__7640),
            .I(P1A3_c));
    InMux I__1205 (
            .O(N__7635),
            .I(N__7631));
    InMux I__1204 (
            .O(N__7634),
            .I(N__7628));
    LocalMux I__1203 (
            .O(N__7631),
            .I(\DUT.uart_inst0.N_82 ));
    LocalMux I__1202 (
            .O(N__7628),
            .I(\DUT.uart_inst0.N_82 ));
    InMux I__1201 (
            .O(N__7623),
            .I(N__7620));
    LocalMux I__1200 (
            .O(N__7620),
            .I(\DUT.uart_inst0.tx_countdown_3_cry_0_c_RNOZ0 ));
    CascadeMux I__1199 (
            .O(N__7617),
            .I(N__7613));
    CascadeMux I__1198 (
            .O(N__7616),
            .I(N__7609));
    InMux I__1197 (
            .O(N__7613),
            .I(N__7606));
    InMux I__1196 (
            .O(N__7612),
            .I(N__7603));
    InMux I__1195 (
            .O(N__7609),
            .I(N__7600));
    LocalMux I__1194 (
            .O(N__7606),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_3 ));
    LocalMux I__1193 (
            .O(N__7603),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_3 ));
    LocalMux I__1192 (
            .O(N__7600),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_3 ));
    InMux I__1191 (
            .O(N__7593),
            .I(\DUT.uart_inst0.tx_countdown_3_cry_0 ));
    InMux I__1190 (
            .O(N__7590),
            .I(N__7587));
    LocalMux I__1189 (
            .O(N__7587),
            .I(\DUT.uart_inst0.tx_countdown_RNI5L692Z0Z_2 ));
    InMux I__1188 (
            .O(N__7584),
            .I(N__7580));
    CascadeMux I__1187 (
            .O(N__7583),
            .I(N__7577));
    LocalMux I__1186 (
            .O(N__7580),
            .I(N__7574));
    InMux I__1185 (
            .O(N__7577),
            .I(N__7571));
    Span12Mux_v I__1184 (
            .O(N__7574),
            .I(N__7568));
    LocalMux I__1183 (
            .O(N__7571),
            .I(N__7565));
    Odrv12 I__1182 (
            .O(N__7568),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_2 ));
    Odrv4 I__1181 (
            .O(N__7565),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_2 ));
    InMux I__1180 (
            .O(N__7560),
            .I(\DUT.uart_inst0.tx_countdown_3_cry_1 ));
    InMux I__1179 (
            .O(N__7557),
            .I(\DUT.uart_inst0.tx_countdown_3_cry_2 ));
    InMux I__1178 (
            .O(N__7554),
            .I(N__7551));
    LocalMux I__1177 (
            .O(N__7551),
            .I(\DUT.uart_inst0.tx_countdown_RNI7N692Z0Z_4 ));
    InMux I__1176 (
            .O(N__7548),
            .I(N__7544));
    CascadeMux I__1175 (
            .O(N__7547),
            .I(N__7541));
    LocalMux I__1174 (
            .O(N__7544),
            .I(N__7538));
    InMux I__1173 (
            .O(N__7541),
            .I(N__7535));
    Odrv4 I__1172 (
            .O(N__7538),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_4 ));
    LocalMux I__1171 (
            .O(N__7535),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_4 ));
    InMux I__1170 (
            .O(N__7530),
            .I(\DUT.uart_inst0.tx_countdown_3_cry_3 ));
    CascadeMux I__1169 (
            .O(N__7527),
            .I(\DUT.uart_inst0.tx_bits_remaining_RNI5UON8Z0Z_3_cascade_ ));
    CascadeMux I__1168 (
            .O(N__7524),
            .I(\DUT.uart_inst0.N_109_cascade_ ));
    CascadeMux I__1167 (
            .O(N__7521),
            .I(\DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIKK41CZ0_cascade_ ));
    InMux I__1166 (
            .O(N__7518),
            .I(N__7515));
    LocalMux I__1165 (
            .O(N__7515),
            .I(\DUT.uart_inst0.N_109 ));
    InMux I__1164 (
            .O(N__7512),
            .I(N__7509));
    LocalMux I__1163 (
            .O(N__7509),
            .I(\DUT.uart_inst0.tx_state_ns_i_i_a3_1_0 ));
    InMux I__1162 (
            .O(N__7506),
            .I(N__7503));
    LocalMux I__1161 (
            .O(N__7503),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_6 ));
    CEMux I__1160 (
            .O(N__7500),
            .I(N__7496));
    CEMux I__1159 (
            .O(N__7499),
            .I(N__7492));
    LocalMux I__1158 (
            .O(N__7496),
            .I(N__7489));
    CEMux I__1157 (
            .O(N__7495),
            .I(N__7486));
    LocalMux I__1156 (
            .O(N__7492),
            .I(N__7483));
    Span4Mux_h I__1155 (
            .O(N__7489),
            .I(N__7478));
    LocalMux I__1154 (
            .O(N__7486),
            .I(N__7478));
    Span4Mux_h I__1153 (
            .O(N__7483),
            .I(N__7475));
    Span4Mux_h I__1152 (
            .O(N__7478),
            .I(N__7472));
    Span4Mux_v I__1151 (
            .O(N__7475),
            .I(N__7469));
    Span4Mux_v I__1150 (
            .O(N__7472),
            .I(N__7466));
    Odrv4 I__1149 (
            .O(N__7469),
            .I(\DUT.uart_inst0.rx_bits_remaining_2_sqmuxa ));
    Odrv4 I__1148 (
            .O(N__7466),
            .I(\DUT.uart_inst0.rx_bits_remaining_2_sqmuxa ));
    CascadeMux I__1147 (
            .O(N__7461),
            .I(\DUT.uart_inst0.g0_0_1_cascade_ ));
    InMux I__1146 (
            .O(N__7458),
            .I(N__7450));
    InMux I__1145 (
            .O(N__7457),
            .I(N__7447));
    InMux I__1144 (
            .O(N__7456),
            .I(N__7440));
    InMux I__1143 (
            .O(N__7455),
            .I(N__7440));
    InMux I__1142 (
            .O(N__7454),
            .I(N__7440));
    InMux I__1141 (
            .O(N__7453),
            .I(N__7437));
    LocalMux I__1140 (
            .O(N__7450),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_0 ));
    LocalMux I__1139 (
            .O(N__7447),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_0 ));
    LocalMux I__1138 (
            .O(N__7440),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_0 ));
    LocalMux I__1137 (
            .O(N__7437),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_0 ));
    InMux I__1136 (
            .O(N__7428),
            .I(N__7424));
    InMux I__1135 (
            .O(N__7427),
            .I(N__7421));
    LocalMux I__1134 (
            .O(N__7424),
            .I(\DUT.uart_inst0.N_62_4 ));
    LocalMux I__1133 (
            .O(N__7421),
            .I(\DUT.uart_inst0.N_62_4 ));
    InMux I__1132 (
            .O(N__7416),
            .I(N__7407));
    InMux I__1131 (
            .O(N__7415),
            .I(N__7407));
    InMux I__1130 (
            .O(N__7414),
            .I(N__7403));
    InMux I__1129 (
            .O(N__7413),
            .I(N__7398));
    InMux I__1128 (
            .O(N__7412),
            .I(N__7398));
    LocalMux I__1127 (
            .O(N__7407),
            .I(N__7395));
    InMux I__1126 (
            .O(N__7406),
            .I(N__7392));
    LocalMux I__1125 (
            .O(N__7403),
            .I(N__7387));
    LocalMux I__1124 (
            .O(N__7398),
            .I(N__7380));
    Span4Mux_h I__1123 (
            .O(N__7395),
            .I(N__7380));
    LocalMux I__1122 (
            .O(N__7392),
            .I(N__7380));
    InMux I__1121 (
            .O(N__7391),
            .I(N__7375));
    InMux I__1120 (
            .O(N__7390),
            .I(N__7375));
    Odrv12 I__1119 (
            .O(N__7387),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    Odrv4 I__1118 (
            .O(N__7380),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    LocalMux I__1117 (
            .O(N__7375),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    CascadeMux I__1116 (
            .O(N__7368),
            .I(\DUT.uart_inst0.recv_state_srsts_1_2_cascade_ ));
    InMux I__1115 (
            .O(N__7365),
            .I(N__7355));
    InMux I__1114 (
            .O(N__7364),
            .I(N__7350));
    InMux I__1113 (
            .O(N__7363),
            .I(N__7350));
    InMux I__1112 (
            .O(N__7362),
            .I(N__7341));
    InMux I__1111 (
            .O(N__7361),
            .I(N__7341));
    InMux I__1110 (
            .O(N__7360),
            .I(N__7341));
    InMux I__1109 (
            .O(N__7359),
            .I(N__7336));
    InMux I__1108 (
            .O(N__7358),
            .I(N__7336));
    LocalMux I__1107 (
            .O(N__7355),
            .I(N__7333));
    LocalMux I__1106 (
            .O(N__7350),
            .I(N__7330));
    InMux I__1105 (
            .O(N__7349),
            .I(N__7325));
    InMux I__1104 (
            .O(N__7348),
            .I(N__7325));
    LocalMux I__1103 (
            .O(N__7341),
            .I(N__7320));
    LocalMux I__1102 (
            .O(N__7336),
            .I(N__7320));
    Span4Mux_h I__1101 (
            .O(N__7333),
            .I(N__7317));
    Odrv4 I__1100 (
            .O(N__7330),
            .I(\DUT.uart_inst0.N_42 ));
    LocalMux I__1099 (
            .O(N__7325),
            .I(\DUT.uart_inst0.N_42 ));
    Odrv4 I__1098 (
            .O(N__7320),
            .I(\DUT.uart_inst0.N_42 ));
    Odrv4 I__1097 (
            .O(N__7317),
            .I(\DUT.uart_inst0.N_42 ));
    InMux I__1096 (
            .O(N__7308),
            .I(N__7303));
    InMux I__1095 (
            .O(N__7307),
            .I(N__7300));
    InMux I__1094 (
            .O(N__7306),
            .I(N__7297));
    LocalMux I__1093 (
            .O(N__7303),
            .I(N__7294));
    LocalMux I__1092 (
            .O(N__7300),
            .I(N__7289));
    LocalMux I__1091 (
            .O(N__7297),
            .I(N__7289));
    Span4Mux_h I__1090 (
            .O(N__7294),
            .I(N__7277));
    Span4Mux_v I__1089 (
            .O(N__7289),
            .I(N__7274));
    InMux I__1088 (
            .O(N__7288),
            .I(N__7267));
    InMux I__1087 (
            .O(N__7287),
            .I(N__7267));
    InMux I__1086 (
            .O(N__7286),
            .I(N__7267));
    InMux I__1085 (
            .O(N__7285),
            .I(N__7262));
    InMux I__1084 (
            .O(N__7284),
            .I(N__7262));
    InMux I__1083 (
            .O(N__7283),
            .I(N__7253));
    InMux I__1082 (
            .O(N__7282),
            .I(N__7253));
    InMux I__1081 (
            .O(N__7281),
            .I(N__7253));
    InMux I__1080 (
            .O(N__7280),
            .I(N__7253));
    Odrv4 I__1079 (
            .O(N__7277),
            .I(\DUT.uart_inst0.recv_stateZ0Z_2 ));
    Odrv4 I__1078 (
            .O(N__7274),
            .I(\DUT.uart_inst0.recv_stateZ0Z_2 ));
    LocalMux I__1077 (
            .O(N__7267),
            .I(\DUT.uart_inst0.recv_stateZ0Z_2 ));
    LocalMux I__1076 (
            .O(N__7262),
            .I(\DUT.uart_inst0.recv_stateZ0Z_2 ));
    LocalMux I__1075 (
            .O(N__7253),
            .I(\DUT.uart_inst0.recv_stateZ0Z_2 ));
    InMux I__1074 (
            .O(N__7242),
            .I(N__7239));
    LocalMux I__1073 (
            .O(N__7239),
            .I(\DUT.uart_inst0.m5_0_0 ));
    InMux I__1072 (
            .O(N__7236),
            .I(N__7230));
    InMux I__1071 (
            .O(N__7235),
            .I(N__7230));
    LocalMux I__1070 (
            .O(N__7230),
            .I(\DUT.fifo_rx_inst.rFifoDataro_0 ));
    InMux I__1069 (
            .O(N__7227),
            .I(N__7221));
    InMux I__1068 (
            .O(N__7226),
            .I(N__7221));
    LocalMux I__1067 (
            .O(N__7221),
            .I(\DUT.fifo_rx_inst.rFifoDataro_1 ));
    InMux I__1066 (
            .O(N__7218),
            .I(N__7215));
    LocalMux I__1065 (
            .O(N__7215),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_1 ));
    InMux I__1064 (
            .O(N__7212),
            .I(N__7209));
    LocalMux I__1063 (
            .O(N__7209),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_7 ));
    CascadeMux I__1062 (
            .O(N__7206),
            .I(\DUT.uart_inst0.tx_countdown_3_0_cascade_ ));
    CascadeMux I__1061 (
            .O(N__7203),
            .I(N__7200));
    InMux I__1060 (
            .O(N__7200),
            .I(N__7196));
    InMux I__1059 (
            .O(N__7199),
            .I(N__7193));
    LocalMux I__1058 (
            .O(N__7196),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_11 ));
    LocalMux I__1057 (
            .O(N__7193),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_11 ));
    InMux I__1056 (
            .O(N__7188),
            .I(N__7184));
    InMux I__1055 (
            .O(N__7187),
            .I(N__7181));
    LocalMux I__1054 (
            .O(N__7184),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_10 ));
    LocalMux I__1053 (
            .O(N__7181),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_10 ));
    CascadeMux I__1052 (
            .O(N__7176),
            .I(N__7173));
    InMux I__1051 (
            .O(N__7173),
            .I(N__7169));
    InMux I__1050 (
            .O(N__7172),
            .I(N__7166));
    LocalMux I__1049 (
            .O(N__7169),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_9 ));
    LocalMux I__1048 (
            .O(N__7166),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_9 ));
    InMux I__1047 (
            .O(N__7161),
            .I(N__7157));
    InMux I__1046 (
            .O(N__7160),
            .I(N__7154));
    LocalMux I__1045 (
            .O(N__7157),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_8 ));
    LocalMux I__1044 (
            .O(N__7154),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_8 ));
    InMux I__1043 (
            .O(N__7149),
            .I(N__7145));
    InMux I__1042 (
            .O(N__7148),
            .I(N__7142));
    LocalMux I__1041 (
            .O(N__7145),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_1 ));
    LocalMux I__1040 (
            .O(N__7142),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_1 ));
    CascadeMux I__1039 (
            .O(N__7137),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_7_cascade_ ));
    CascadeMux I__1038 (
            .O(N__7134),
            .I(N__7130));
    InMux I__1037 (
            .O(N__7133),
            .I(N__7126));
    InMux I__1036 (
            .O(N__7130),
            .I(N__7123));
    InMux I__1035 (
            .O(N__7129),
            .I(N__7120));
    LocalMux I__1034 (
            .O(N__7126),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_0 ));
    LocalMux I__1033 (
            .O(N__7123),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_0 ));
    LocalMux I__1032 (
            .O(N__7120),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_0 ));
    CascadeMux I__1031 (
            .O(N__7113),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_10_cascade_ ));
    CascadeMux I__1030 (
            .O(N__7110),
            .I(\DUT.uart_inst0.tx_clk_divider_1_sqmuxa_1_0_cascade_ ));
    SRMux I__1029 (
            .O(N__7107),
            .I(N__7103));
    SRMux I__1028 (
            .O(N__7106),
            .I(N__7100));
    LocalMux I__1027 (
            .O(N__7103),
            .I(\DUT.uart_inst0.tx_clk_divider_1_sqmuxa_1_i ));
    LocalMux I__1026 (
            .O(N__7100),
            .I(\DUT.uart_inst0.tx_clk_divider_1_sqmuxa_1_i ));
    InMux I__1025 (
            .O(N__7095),
            .I(N__7092));
    LocalMux I__1024 (
            .O(N__7092),
            .I(N__7089));
    Odrv12 I__1023 (
            .O(N__7089),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_5 ));
    CascadeMux I__1022 (
            .O(N__7086),
            .I(N__7082));
    InMux I__1021 (
            .O(N__7085),
            .I(N__7075));
    InMux I__1020 (
            .O(N__7082),
            .I(N__7075));
    InMux I__1019 (
            .O(N__7081),
            .I(N__7072));
    CascadeMux I__1018 (
            .O(N__7080),
            .I(N__7069));
    LocalMux I__1017 (
            .O(N__7075),
            .I(N__7064));
    LocalMux I__1016 (
            .O(N__7072),
            .I(N__7064));
    InMux I__1015 (
            .O(N__7069),
            .I(N__7061));
    Span4Mux_v I__1014 (
            .O(N__7064),
            .I(N__7058));
    LocalMux I__1013 (
            .O(N__7061),
            .I(N__7054));
    Span4Mux_h I__1012 (
            .O(N__7058),
            .I(N__7051));
    InMux I__1011 (
            .O(N__7057),
            .I(N__7048));
    Odrv12 I__1010 (
            .O(N__7054),
            .I(\DUT.uart_inst0.N_47 ));
    Odrv4 I__1009 (
            .O(N__7051),
            .I(\DUT.uart_inst0.N_47 ));
    LocalMux I__1008 (
            .O(N__7048),
            .I(\DUT.uart_inst0.N_47 ));
    InMux I__1007 (
            .O(N__7041),
            .I(N__7038));
    LocalMux I__1006 (
            .O(N__7038),
            .I(\DUT.uart_inst0.N_68 ));
    CascadeMux I__1005 (
            .O(N__7035),
            .I(N__7031));
    CascadeMux I__1004 (
            .O(N__7034),
            .I(N__7028));
    InMux I__1003 (
            .O(N__7031),
            .I(N__7024));
    InMux I__1002 (
            .O(N__7028),
            .I(N__7019));
    InMux I__1001 (
            .O(N__7027),
            .I(N__7019));
    LocalMux I__1000 (
            .O(N__7024),
            .I(N__7012));
    LocalMux I__999 (
            .O(N__7019),
            .I(N__7009));
    InMux I__998 (
            .O(N__7018),
            .I(N__7002));
    InMux I__997 (
            .O(N__7017),
            .I(N__7002));
    InMux I__996 (
            .O(N__7016),
            .I(N__7002));
    CascadeMux I__995 (
            .O(N__7015),
            .I(N__6999));
    Span4Mux_v I__994 (
            .O(N__7012),
            .I(N__6992));
    Span4Mux_v I__993 (
            .O(N__7009),
            .I(N__6992));
    LocalMux I__992 (
            .O(N__7002),
            .I(N__6992));
    InMux I__991 (
            .O(N__6999),
            .I(N__6989));
    Span4Mux_h I__990 (
            .O(N__6992),
            .I(N__6986));
    LocalMux I__989 (
            .O(N__6989),
            .I(\DUT.uart_inst0.recv_stateZ0Z_5 ));
    Odrv4 I__988 (
            .O(N__6986),
            .I(\DUT.uart_inst0.recv_stateZ0Z_5 ));
    CascadeMux I__987 (
            .O(N__6981),
            .I(N__6977));
    InMux I__986 (
            .O(N__6980),
            .I(N__6974));
    InMux I__985 (
            .O(N__6977),
            .I(N__6971));
    LocalMux I__984 (
            .O(N__6974),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_2 ));
    LocalMux I__983 (
            .O(N__6971),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_2 ));
    InMux I__982 (
            .O(N__6966),
            .I(N__6961));
    InMux I__981 (
            .O(N__6965),
            .I(N__6956));
    InMux I__980 (
            .O(N__6964),
            .I(N__6956));
    LocalMux I__979 (
            .O(N__6961),
            .I(\DUT.uart_inst0.rx_countdown_3_2 ));
    LocalMux I__978 (
            .O(N__6956),
            .I(\DUT.uart_inst0.rx_countdown_3_2 ));
    CascadeMux I__977 (
            .O(N__6951),
            .I(N__6948));
    InMux I__976 (
            .O(N__6948),
            .I(N__6945));
    LocalMux I__975 (
            .O(N__6945),
            .I(N__6939));
    InMux I__974 (
            .O(N__6944),
            .I(N__6934));
    InMux I__973 (
            .O(N__6943),
            .I(N__6934));
    InMux I__972 (
            .O(N__6942),
            .I(N__6931));
    Odrv12 I__971 (
            .O(N__6939),
            .I(\DUT.uart_inst0.rx_countdown_3_3 ));
    LocalMux I__970 (
            .O(N__6934),
            .I(\DUT.uart_inst0.rx_countdown_3_3 ));
    LocalMux I__969 (
            .O(N__6931),
            .I(\DUT.uart_inst0.rx_countdown_3_3 ));
    InMux I__968 (
            .O(N__6924),
            .I(N__6918));
    InMux I__967 (
            .O(N__6923),
            .I(N__6913));
    InMux I__966 (
            .O(N__6922),
            .I(N__6913));
    InMux I__965 (
            .O(N__6921),
            .I(N__6910));
    LocalMux I__964 (
            .O(N__6918),
            .I(\DUT.uart_inst0.rx_countdown_3_4 ));
    LocalMux I__963 (
            .O(N__6913),
            .I(\DUT.uart_inst0.rx_countdown_3_4 ));
    LocalMux I__962 (
            .O(N__6910),
            .I(\DUT.uart_inst0.rx_countdown_3_4 ));
    CascadeMux I__961 (
            .O(N__6903),
            .I(\DUT.uart_inst0.rx_bits_remaining_2_sqmuxa_0_a2_0_a2_1_cascade_ ));
    InMux I__960 (
            .O(N__6900),
            .I(N__6896));
    InMux I__959 (
            .O(N__6899),
            .I(N__6893));
    LocalMux I__958 (
            .O(N__6896),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_2_2 ));
    LocalMux I__957 (
            .O(N__6893),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_2_2 ));
    InMux I__956 (
            .O(N__6888),
            .I(N__6884));
    InMux I__955 (
            .O(N__6887),
            .I(N__6881));
    LocalMux I__954 (
            .O(N__6884),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_12 ));
    LocalMux I__953 (
            .O(N__6881),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_12 ));
    InMux I__952 (
            .O(N__6876),
            .I(N__6872));
    InMux I__951 (
            .O(N__6875),
            .I(N__6869));
    LocalMux I__950 (
            .O(N__6872),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_7 ));
    LocalMux I__949 (
            .O(N__6869),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_7 ));
    CascadeMux I__948 (
            .O(N__6864),
            .I(N__6861));
    InMux I__947 (
            .O(N__6861),
            .I(N__6857));
    InMux I__946 (
            .O(N__6860),
            .I(N__6854));
    LocalMux I__945 (
            .O(N__6857),
            .I(N__6851));
    LocalMux I__944 (
            .O(N__6854),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_13 ));
    Odrv4 I__943 (
            .O(N__6851),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_13 ));
    CascadeMux I__942 (
            .O(N__6846),
            .I(N__6843));
    InMux I__941 (
            .O(N__6843),
            .I(N__6839));
    InMux I__940 (
            .O(N__6842),
            .I(N__6836));
    LocalMux I__939 (
            .O(N__6839),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_6 ));
    LocalMux I__938 (
            .O(N__6836),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_6 ));
    CascadeMux I__937 (
            .O(N__6831),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_8_cascade_ ));
    CascadeMux I__936 (
            .O(N__6828),
            .I(N__6825));
    InMux I__935 (
            .O(N__6825),
            .I(N__6821));
    InMux I__934 (
            .O(N__6824),
            .I(N__6818));
    LocalMux I__933 (
            .O(N__6821),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_4 ));
    LocalMux I__932 (
            .O(N__6818),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_4 ));
    InMux I__931 (
            .O(N__6813),
            .I(N__6809));
    InMux I__930 (
            .O(N__6812),
            .I(N__6806));
    LocalMux I__929 (
            .O(N__6809),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_3 ));
    LocalMux I__928 (
            .O(N__6806),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_3 ));
    CascadeMux I__927 (
            .O(N__6801),
            .I(N__6798));
    InMux I__926 (
            .O(N__6798),
            .I(N__6794));
    InMux I__925 (
            .O(N__6797),
            .I(N__6791));
    LocalMux I__924 (
            .O(N__6794),
            .I(N__6788));
    LocalMux I__923 (
            .O(N__6791),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_5 ));
    Odrv4 I__922 (
            .O(N__6788),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_5 ));
    CascadeMux I__921 (
            .O(N__6783),
            .I(N__6780));
    InMux I__920 (
            .O(N__6780),
            .I(N__6776));
    InMux I__919 (
            .O(N__6779),
            .I(N__6773));
    LocalMux I__918 (
            .O(N__6776),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_2 ));
    LocalMux I__917 (
            .O(N__6773),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_2 ));
    CascadeMux I__916 (
            .O(N__6768),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_9_cascade_ ));
    CascadeMux I__915 (
            .O(N__6765),
            .I(N__6760));
    CascadeMux I__914 (
            .O(N__6764),
            .I(N__6757));
    InMux I__913 (
            .O(N__6763),
            .I(N__6753));
    InMux I__912 (
            .O(N__6760),
            .I(N__6748));
    InMux I__911 (
            .O(N__6757),
            .I(N__6748));
    InMux I__910 (
            .O(N__6756),
            .I(N__6745));
    LocalMux I__909 (
            .O(N__6753),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    LocalMux I__908 (
            .O(N__6748),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    LocalMux I__907 (
            .O(N__6745),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    CascadeMux I__906 (
            .O(N__6738),
            .I(N__6735));
    InMux I__905 (
            .O(N__6735),
            .I(N__6732));
    LocalMux I__904 (
            .O(N__6732),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_0_c_RNOZ0 ));
    InMux I__903 (
            .O(N__6729),
            .I(N__6725));
    InMux I__902 (
            .O(N__6728),
            .I(N__6722));
    LocalMux I__901 (
            .O(N__6725),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_1 ));
    LocalMux I__900 (
            .O(N__6722),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_1 ));
    CascadeMux I__899 (
            .O(N__6717),
            .I(N__6714));
    InMux I__898 (
            .O(N__6714),
            .I(N__6711));
    LocalMux I__897 (
            .O(N__6711),
            .I(\DUT.uart_inst0.rx_countdown_RNICSMA4Z0Z_1 ));
    InMux I__896 (
            .O(N__6708),
            .I(N__6704));
    InMux I__895 (
            .O(N__6707),
            .I(N__6701));
    LocalMux I__894 (
            .O(N__6704),
            .I(\DUT.uart_inst0.rx_countdown_3_1 ));
    LocalMux I__893 (
            .O(N__6701),
            .I(\DUT.uart_inst0.rx_countdown_3_1 ));
    InMux I__892 (
            .O(N__6696),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_0 ));
    InMux I__891 (
            .O(N__6693),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_1 ));
    InMux I__890 (
            .O(N__6690),
            .I(N__6686));
    InMux I__889 (
            .O(N__6689),
            .I(N__6683));
    LocalMux I__888 (
            .O(N__6686),
            .I(\DUT.uart_inst0.rx_countdownZ1Z_3 ));
    LocalMux I__887 (
            .O(N__6683),
            .I(\DUT.uart_inst0.rx_countdownZ1Z_3 ));
    CascadeMux I__886 (
            .O(N__6678),
            .I(N__6675));
    InMux I__885 (
            .O(N__6675),
            .I(N__6672));
    LocalMux I__884 (
            .O(N__6672),
            .I(N__6669));
    Odrv4 I__883 (
            .O(N__6669),
            .I(\DUT.uart_inst0.rx_countdown_RNIEUMA4Z0Z_3 ));
    InMux I__882 (
            .O(N__6666),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_2 ));
    InMux I__881 (
            .O(N__6663),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_3 ));
    InMux I__880 (
            .O(N__6660),
            .I(N__6657));
    LocalMux I__879 (
            .O(N__6657),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_5 ));
    InMux I__878 (
            .O(N__6654),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_4 ));
    CascadeMux I__877 (
            .O(N__6651),
            .I(N__6648));
    InMux I__876 (
            .O(N__6648),
            .I(N__6645));
    LocalMux I__875 (
            .O(N__6645),
            .I(N__6641));
    InMux I__874 (
            .O(N__6644),
            .I(N__6638));
    Odrv4 I__873 (
            .O(N__6641),
            .I(\DUT.uart_inst0.rx_countdown_3_5 ));
    LocalMux I__872 (
            .O(N__6638),
            .I(\DUT.uart_inst0.rx_countdown_3_5 ));
    CascadeMux I__871 (
            .O(N__6633),
            .I(N__6629));
    InMux I__870 (
            .O(N__6632),
            .I(N__6624));
    InMux I__869 (
            .O(N__6629),
            .I(N__6624));
    LocalMux I__868 (
            .O(N__6624),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_4 ));
    InMux I__867 (
            .O(N__6621),
            .I(N__6618));
    LocalMux I__866 (
            .O(N__6618),
            .I(\DUT.uart_inst0.rx_countdown_RNIFVMA4Z0Z_4 ));
    InMux I__865 (
            .O(N__6615),
            .I(N__6604));
    InMux I__864 (
            .O(N__6614),
            .I(N__6604));
    CascadeMux I__863 (
            .O(N__6613),
            .I(N__6601));
    CascadeMux I__862 (
            .O(N__6612),
            .I(N__6597));
    CascadeMux I__861 (
            .O(N__6611),
            .I(N__6592));
    InMux I__860 (
            .O(N__6610),
            .I(N__6589));
    InMux I__859 (
            .O(N__6609),
            .I(N__6586));
    LocalMux I__858 (
            .O(N__6604),
            .I(N__6583));
    InMux I__857 (
            .O(N__6601),
            .I(N__6578));
    InMux I__856 (
            .O(N__6600),
            .I(N__6578));
    InMux I__855 (
            .O(N__6597),
            .I(N__6571));
    InMux I__854 (
            .O(N__6596),
            .I(N__6571));
    InMux I__853 (
            .O(N__6595),
            .I(N__6571));
    InMux I__852 (
            .O(N__6592),
            .I(N__6568));
    LocalMux I__851 (
            .O(N__6589),
            .I(N__6565));
    LocalMux I__850 (
            .O(N__6586),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_15 ));
    Odrv4 I__849 (
            .O(N__6583),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_15 ));
    LocalMux I__848 (
            .O(N__6578),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_15 ));
    LocalMux I__847 (
            .O(N__6571),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_15 ));
    LocalMux I__846 (
            .O(N__6568),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_15 ));
    Odrv4 I__845 (
            .O(N__6565),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_15 ));
    InMux I__844 (
            .O(N__6552),
            .I(N__6538));
    InMux I__843 (
            .O(N__6551),
            .I(N__6538));
    InMux I__842 (
            .O(N__6550),
            .I(N__6538));
    InMux I__841 (
            .O(N__6549),
            .I(N__6533));
    InMux I__840 (
            .O(N__6548),
            .I(N__6533));
    InMux I__839 (
            .O(N__6547),
            .I(N__6528));
    InMux I__838 (
            .O(N__6546),
            .I(N__6528));
    InMux I__837 (
            .O(N__6545),
            .I(N__6525));
    LocalMux I__836 (
            .O(N__6538),
            .I(N__6519));
    LocalMux I__835 (
            .O(N__6533),
            .I(N__6512));
    LocalMux I__834 (
            .O(N__6528),
            .I(N__6512));
    LocalMux I__833 (
            .O(N__6525),
            .I(N__6512));
    InMux I__832 (
            .O(N__6524),
            .I(N__6507));
    InMux I__831 (
            .O(N__6523),
            .I(N__6507));
    InMux I__830 (
            .O(N__6522),
            .I(N__6504));
    Span4Mux_h I__829 (
            .O(N__6519),
            .I(N__6497));
    Span4Mux_v I__828 (
            .O(N__6512),
            .I(N__6497));
    LocalMux I__827 (
            .O(N__6507),
            .I(N__6497));
    LocalMux I__826 (
            .O(N__6504),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_14 ));
    Odrv4 I__825 (
            .O(N__6497),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_14 ));
    InMux I__824 (
            .O(N__6492),
            .I(N__6489));
    LocalMux I__823 (
            .O(N__6489),
            .I(\DUT.uart_inst0.rx_countdown_RNIDTMA4Z0Z_2 ));
    IoInMux I__822 (
            .O(N__6486),
            .I(N__6483));
    LocalMux I__821 (
            .O(N__6483),
            .I(wPllLocked_i));
    InMux I__820 (
            .O(N__6480),
            .I(N__6477));
    LocalMux I__819 (
            .O(N__6477),
            .I(N__6474));
    Odrv4 I__818 (
            .O(N__6474),
            .I(\DUT.uart_inst0.rx_clk_divider_1_5 ));
    InMux I__817 (
            .O(N__6471),
            .I(N__6467));
    InMux I__816 (
            .O(N__6470),
            .I(N__6464));
    LocalMux I__815 (
            .O(N__6467),
            .I(N__6459));
    LocalMux I__814 (
            .O(N__6464),
            .I(N__6459));
    Odrv12 I__813 (
            .O(N__6459),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_5 ));
    InMux I__812 (
            .O(N__6456),
            .I(N__6453));
    LocalMux I__811 (
            .O(N__6453),
            .I(N__6450));
    Odrv4 I__810 (
            .O(N__6450),
            .I(\DUT.uart_inst0.rx_clk_divider_1_6 ));
    CascadeMux I__809 (
            .O(N__6447),
            .I(N__6444));
    InMux I__808 (
            .O(N__6444),
            .I(N__6440));
    InMux I__807 (
            .O(N__6443),
            .I(N__6437));
    LocalMux I__806 (
            .O(N__6440),
            .I(N__6432));
    LocalMux I__805 (
            .O(N__6437),
            .I(N__6432));
    Span4Mux_h I__804 (
            .O(N__6432),
            .I(N__6429));
    Odrv4 I__803 (
            .O(N__6429),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_6 ));
    InMux I__802 (
            .O(N__6426),
            .I(N__6423));
    LocalMux I__801 (
            .O(N__6423),
            .I(\DUT.fifo_rx_inst.un1_i11_2_i ));
    CascadeMux I__800 (
            .O(N__6420),
            .I(\DUT.fifo_rx_inst.un1_i11_2_i_cascade_ ));
    CascadeMux I__799 (
            .O(N__6417),
            .I(N__6413));
    InMux I__798 (
            .O(N__6416),
            .I(N__6408));
    InMux I__797 (
            .O(N__6413),
            .I(N__6401));
    InMux I__796 (
            .O(N__6412),
            .I(N__6401));
    InMux I__795 (
            .O(N__6411),
            .I(N__6401));
    LocalMux I__794 (
            .O(N__6408),
            .I(\DUT.fifo_rx_inst.N_88 ));
    LocalMux I__793 (
            .O(N__6401),
            .I(\DUT.fifo_rx_inst.N_88 ));
    InMux I__792 (
            .O(N__6396),
            .I(N__6386));
    InMux I__791 (
            .O(N__6395),
            .I(N__6386));
    InMux I__790 (
            .O(N__6394),
            .I(N__6386));
    CascadeMux I__789 (
            .O(N__6393),
            .I(N__6381));
    LocalMux I__788 (
            .O(N__6386),
            .I(N__6378));
    InMux I__787 (
            .O(N__6385),
            .I(N__6371));
    InMux I__786 (
            .O(N__6384),
            .I(N__6371));
    InMux I__785 (
            .O(N__6381),
            .I(N__6371));
    Odrv4 I__784 (
            .O(N__6378),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_0 ));
    LocalMux I__783 (
            .O(N__6371),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_0 ));
    InMux I__782 (
            .O(N__6366),
            .I(N__6360));
    InMux I__781 (
            .O(N__6365),
            .I(N__6355));
    InMux I__780 (
            .O(N__6364),
            .I(N__6355));
    CascadeMux I__779 (
            .O(N__6363),
            .I(N__6352));
    LocalMux I__778 (
            .O(N__6360),
            .I(N__6346));
    LocalMux I__777 (
            .O(N__6355),
            .I(N__6346));
    InMux I__776 (
            .O(N__6352),
            .I(N__6341));
    InMux I__775 (
            .O(N__6351),
            .I(N__6341));
    Odrv4 I__774 (
            .O(N__6346),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_1 ));
    LocalMux I__773 (
            .O(N__6341),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_1 ));
    InMux I__772 (
            .O(N__6336),
            .I(N__6327));
    InMux I__771 (
            .O(N__6335),
            .I(N__6327));
    InMux I__770 (
            .O(N__6334),
            .I(N__6320));
    InMux I__769 (
            .O(N__6333),
            .I(N__6320));
    InMux I__768 (
            .O(N__6332),
            .I(N__6320));
    LocalMux I__767 (
            .O(N__6327),
            .I(\DUT.fifo_rx_inst.N_85 ));
    LocalMux I__766 (
            .O(N__6320),
            .I(\DUT.fifo_rx_inst.N_85 ));
    CascadeMux I__765 (
            .O(N__6315),
            .I(N__6309));
    CascadeMux I__764 (
            .O(N__6314),
            .I(N__6306));
    InMux I__763 (
            .O(N__6313),
            .I(N__6302));
    InMux I__762 (
            .O(N__6312),
            .I(N__6293));
    InMux I__761 (
            .O(N__6309),
            .I(N__6293));
    InMux I__760 (
            .O(N__6306),
            .I(N__6293));
    InMux I__759 (
            .O(N__6305),
            .I(N__6293));
    LocalMux I__758 (
            .O(N__6302),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_1 ));
    LocalMux I__757 (
            .O(N__6293),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_1 ));
    CascadeMux I__756 (
            .O(N__6288),
            .I(\DUT.uart_inst0.m5_1_cascade_ ));
    CascadeMux I__755 (
            .O(N__6285),
            .I(N__6282));
    InMux I__754 (
            .O(N__6282),
            .I(N__6279));
    LocalMux I__753 (
            .O(N__6279),
            .I(N__6276));
    Odrv4 I__752 (
            .O(N__6276),
            .I(\DUT.uart_inst0.N_6_0 ));
    CascadeMux I__751 (
            .O(N__6273),
            .I(\DUT.uart_inst0.N_12_cascade_ ));
    CascadeMux I__750 (
            .O(N__6270),
            .I(\DUT.uart_inst0.N_7_0_cascade_ ));
    CascadeMux I__749 (
            .O(N__6267),
            .I(N__6262));
    InMux I__748 (
            .O(N__6266),
            .I(N__6255));
    InMux I__747 (
            .O(N__6265),
            .I(N__6255));
    InMux I__746 (
            .O(N__6262),
            .I(N__6255));
    LocalMux I__745 (
            .O(N__6255),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_3 ));
    CascadeMux I__744 (
            .O(N__6252),
            .I(\DUT.uart_inst0.m5_0_1_cascade_ ));
    CascadeMux I__743 (
            .O(N__6249),
            .I(\DUT.uart_inst0.N_6_cascade_ ));
    InMux I__742 (
            .O(N__6246),
            .I(N__6234));
    InMux I__741 (
            .O(N__6245),
            .I(N__6234));
    InMux I__740 (
            .O(N__6244),
            .I(N__6234));
    InMux I__739 (
            .O(N__6243),
            .I(N__6234));
    LocalMux I__738 (
            .O(N__6234),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_2 ));
    InMux I__737 (
            .O(N__6231),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_4 ));
    InMux I__736 (
            .O(N__6228),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_5 ));
    InMux I__735 (
            .O(N__6225),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_6 ));
    InMux I__734 (
            .O(N__6222),
            .I(bfn_12_15_0_));
    InMux I__733 (
            .O(N__6219),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_8 ));
    InMux I__732 (
            .O(N__6216),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_9 ));
    InMux I__731 (
            .O(N__6213),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_10 ));
    InMux I__730 (
            .O(N__6210),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_11 ));
    InMux I__729 (
            .O(N__6207),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_12 ));
    CascadeMux I__728 (
            .O(N__6204),
            .I(\DUT.uart_inst0.rx_countdown_RNI8KQG9Z0Z_0_cascade_ ));
    CascadeMux I__727 (
            .O(N__6201),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_2_2_cascade_ ));
    CascadeMux I__726 (
            .O(N__6198),
            .I(\DUT.uart_inst0.N_42_cascade_ ));
    InMux I__725 (
            .O(N__6195),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_0 ));
    InMux I__724 (
            .O(N__6192),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_1 ));
    InMux I__723 (
            .O(N__6189),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_2 ));
    InMux I__722 (
            .O(N__6186),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_3 ));
    InMux I__721 (
            .O(N__6183),
            .I(N__6180));
    LocalMux I__720 (
            .O(N__6180),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO ));
    CascadeMux I__719 (
            .O(N__6177),
            .I(N__6172));
    InMux I__718 (
            .O(N__6176),
            .I(N__6169));
    InMux I__717 (
            .O(N__6175),
            .I(N__6166));
    InMux I__716 (
            .O(N__6172),
            .I(N__6163));
    LocalMux I__715 (
            .O(N__6169),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_13 ));
    LocalMux I__714 (
            .O(N__6166),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_13 ));
    LocalMux I__713 (
            .O(N__6163),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_13 ));
    CascadeMux I__712 (
            .O(N__6156),
            .I(N__6153));
    InMux I__711 (
            .O(N__6153),
            .I(N__6150));
    LocalMux I__710 (
            .O(N__6150),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO ));
    CascadeMux I__709 (
            .O(N__6147),
            .I(N__6143));
    InMux I__708 (
            .O(N__6146),
            .I(N__6139));
    InMux I__707 (
            .O(N__6143),
            .I(N__6136));
    InMux I__706 (
            .O(N__6142),
            .I(N__6133));
    LocalMux I__705 (
            .O(N__6139),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_14 ));
    LocalMux I__704 (
            .O(N__6136),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_14 ));
    LocalMux I__703 (
            .O(N__6133),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_14 ));
    InMux I__702 (
            .O(N__6126),
            .I(N__6123));
    LocalMux I__701 (
            .O(N__6123),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO ));
    InMux I__700 (
            .O(N__6120),
            .I(N__6115));
    InMux I__699 (
            .O(N__6119),
            .I(N__6112));
    InMux I__698 (
            .O(N__6118),
            .I(N__6109));
    LocalMux I__697 (
            .O(N__6115),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_15 ));
    LocalMux I__696 (
            .O(N__6112),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_15 ));
    LocalMux I__695 (
            .O(N__6109),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_15 ));
    CascadeMux I__694 (
            .O(N__6102),
            .I(N__6099));
    InMux I__693 (
            .O(N__6099),
            .I(N__6096));
    LocalMux I__692 (
            .O(N__6096),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO ));
    CascadeMux I__691 (
            .O(N__6093),
            .I(N__6089));
    InMux I__690 (
            .O(N__6092),
            .I(N__6085));
    InMux I__689 (
            .O(N__6089),
            .I(N__6082));
    InMux I__688 (
            .O(N__6088),
            .I(N__6079));
    LocalMux I__687 (
            .O(N__6085),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_16 ));
    LocalMux I__686 (
            .O(N__6082),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_16 ));
    LocalMux I__685 (
            .O(N__6079),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_16 ));
    CascadeMux I__684 (
            .O(N__6072),
            .I(\DUT.uart_inst0.N_46_cascade_ ));
    InMux I__683 (
            .O(N__6069),
            .I(N__6066));
    LocalMux I__682 (
            .O(N__6066),
            .I(\DUT.uart_inst0.rx_countdown_3_0 ));
    InMux I__681 (
            .O(N__6063),
            .I(N__6060));
    LocalMux I__680 (
            .O(N__6060),
            .I(\DUT.fifo_rx_inst.N_97 ));
    CascadeMux I__679 (
            .O(N__6057),
            .I(N__6054));
    InMux I__678 (
            .O(N__6054),
            .I(N__6047));
    InMux I__677 (
            .O(N__6053),
            .I(N__6044));
    InMux I__676 (
            .O(N__6052),
            .I(N__6037));
    InMux I__675 (
            .O(N__6051),
            .I(N__6037));
    InMux I__674 (
            .O(N__6050),
            .I(N__6037));
    LocalMux I__673 (
            .O(N__6047),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_0 ));
    LocalMux I__672 (
            .O(N__6044),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_0 ));
    LocalMux I__671 (
            .O(N__6037),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_0 ));
    InMux I__670 (
            .O(N__6030),
            .I(N__6020));
    InMux I__669 (
            .O(N__6029),
            .I(N__6015));
    InMux I__668 (
            .O(N__6028),
            .I(N__6015));
    InMux I__667 (
            .O(N__6027),
            .I(N__6012));
    InMux I__666 (
            .O(N__6026),
            .I(N__6009));
    InMux I__665 (
            .O(N__6025),
            .I(N__6004));
    InMux I__664 (
            .O(N__6024),
            .I(N__6004));
    InMux I__663 (
            .O(N__6023),
            .I(N__6001));
    LocalMux I__662 (
            .O(N__6020),
            .I(N__5996));
    LocalMux I__661 (
            .O(N__6015),
            .I(N__5996));
    LocalMux I__660 (
            .O(N__6012),
            .I(\DUT.wRcvd ));
    LocalMux I__659 (
            .O(N__6009),
            .I(\DUT.wRcvd ));
    LocalMux I__658 (
            .O(N__6004),
            .I(\DUT.wRcvd ));
    LocalMux I__657 (
            .O(N__6001),
            .I(\DUT.wRcvd ));
    Odrv4 I__656 (
            .O(N__5996),
            .I(\DUT.wRcvd ));
    CascadeMux I__655 (
            .O(N__5985),
            .I(N__5982));
    InMux I__654 (
            .O(N__5982),
            .I(N__5973));
    InMux I__653 (
            .O(N__5981),
            .I(N__5970));
    InMux I__652 (
            .O(N__5980),
            .I(N__5965));
    InMux I__651 (
            .O(N__5979),
            .I(N__5965));
    InMux I__650 (
            .O(N__5978),
            .I(N__5958));
    InMux I__649 (
            .O(N__5977),
            .I(N__5958));
    InMux I__648 (
            .O(N__5976),
            .I(N__5958));
    LocalMux I__647 (
            .O(N__5973),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ));
    LocalMux I__646 (
            .O(N__5970),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ));
    LocalMux I__645 (
            .O(N__5965),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ));
    LocalMux I__644 (
            .O(N__5958),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ));
    InMux I__643 (
            .O(N__5949),
            .I(N__5944));
    InMux I__642 (
            .O(N__5948),
            .I(N__5941));
    InMux I__641 (
            .O(N__5947),
            .I(N__5938));
    LocalMux I__640 (
            .O(N__5944),
            .I(\DUT.uart_inst0.rx_clk_dividerZ1Z_1 ));
    LocalMux I__639 (
            .O(N__5941),
            .I(\DUT.uart_inst0.rx_clk_dividerZ1Z_1 ));
    LocalMux I__638 (
            .O(N__5938),
            .I(\DUT.uart_inst0.rx_clk_dividerZ1Z_1 ));
    InMux I__637 (
            .O(N__5931),
            .I(N__5927));
    InMux I__636 (
            .O(N__5930),
            .I(N__5924));
    LocalMux I__635 (
            .O(N__5927),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_3 ));
    LocalMux I__634 (
            .O(N__5924),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_3 ));
    CascadeMux I__633 (
            .O(N__5919),
            .I(N__5916));
    InMux I__632 (
            .O(N__5916),
            .I(N__5912));
    InMux I__631 (
            .O(N__5915),
            .I(N__5908));
    LocalMux I__630 (
            .O(N__5912),
            .I(N__5905));
    InMux I__629 (
            .O(N__5911),
            .I(N__5902));
    LocalMux I__628 (
            .O(N__5908),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_2 ));
    Odrv4 I__627 (
            .O(N__5905),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_2 ));
    LocalMux I__626 (
            .O(N__5902),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_2 ));
    CascadeMux I__625 (
            .O(N__5895),
            .I(N__5891));
    InMux I__624 (
            .O(N__5894),
            .I(N__5887));
    InMux I__623 (
            .O(N__5891),
            .I(N__5884));
    InMux I__622 (
            .O(N__5890),
            .I(N__5881));
    LocalMux I__621 (
            .O(N__5887),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_1 ));
    LocalMux I__620 (
            .O(N__5884),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_1 ));
    LocalMux I__619 (
            .O(N__5881),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_1 ));
    CascadeMux I__618 (
            .O(N__5874),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_9_cascade_ ));
    CascadeMux I__617 (
            .O(N__5871),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_15_cascade_ ));
    CascadeMux I__616 (
            .O(N__5868),
            .I(N__5864));
    InMux I__615 (
            .O(N__5867),
            .I(N__5861));
    InMux I__614 (
            .O(N__5864),
            .I(N__5858));
    LocalMux I__613 (
            .O(N__5861),
            .I(N__5855));
    LocalMux I__612 (
            .O(N__5858),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_17 ));
    Odrv4 I__611 (
            .O(N__5855),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_17 ));
    InMux I__610 (
            .O(N__5850),
            .I(N__5847));
    LocalMux I__609 (
            .O(N__5847),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_12 ));
    InMux I__608 (
            .O(N__5844),
            .I(N__5841));
    LocalMux I__607 (
            .O(N__5841),
            .I(\DUT.uart_inst0.N_50 ));
    CascadeMux I__606 (
            .O(N__5838),
            .I(\DUT.uart_inst0.recv_state_srsts_1_3_cascade_ ));
    InMux I__605 (
            .O(N__5835),
            .I(N__5826));
    InMux I__604 (
            .O(N__5834),
            .I(N__5826));
    InMux I__603 (
            .O(N__5833),
            .I(N__5826));
    LocalMux I__602 (
            .O(N__5826),
            .I(\DUT.uart_inst0.recv_stateZ0Z_3 ));
    CascadeMux I__601 (
            .O(N__5823),
            .I(\DUT.fifo_rx_inst.N_88_cascade_ ));
    CascadeMux I__600 (
            .O(N__5820),
            .I(N__5817));
    InMux I__599 (
            .O(N__5817),
            .I(N__5814));
    LocalMux I__598 (
            .O(N__5814),
            .I(\DUT.fifo_rx_inst.rFifoCount_RNIK3G92Z0Z_1 ));
    CascadeMux I__597 (
            .O(N__5811),
            .I(N__5806));
    InMux I__596 (
            .O(N__5810),
            .I(N__5802));
    InMux I__595 (
            .O(N__5809),
            .I(N__5795));
    InMux I__594 (
            .O(N__5806),
            .I(N__5795));
    InMux I__593 (
            .O(N__5805),
            .I(N__5795));
    LocalMux I__592 (
            .O(N__5802),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_1 ));
    LocalMux I__591 (
            .O(N__5795),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_1 ));
    CascadeMux I__590 (
            .O(N__5790),
            .I(\DUT.fifo_rx_inst.rFifoCount_RNIHH0D1Z0Z_0_cascade_ ));
    CascadeMux I__589 (
            .O(N__5787),
            .I(\DUT.fifo_rx_inst.N_97_cascade_ ));
    CascadeMux I__588 (
            .O(N__5784),
            .I(N__5781));
    InMux I__587 (
            .O(N__5781),
            .I(N__5778));
    LocalMux I__586 (
            .O(N__5778),
            .I(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0 ));
    InMux I__585 (
            .O(N__5775),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_12 ));
    InMux I__584 (
            .O(N__5772),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_13 ));
    InMux I__583 (
            .O(N__5769),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_14 ));
    InMux I__582 (
            .O(N__5766),
            .I(bfn_11_13_0_));
    InMux I__581 (
            .O(N__5763),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_16 ));
    InMux I__580 (
            .O(N__5760),
            .I(N__5754));
    InMux I__579 (
            .O(N__5759),
            .I(N__5754));
    LocalMux I__578 (
            .O(N__5754),
            .I(\DUT.uart_inst0.recv_stateZ0Z_4 ));
    CascadeMux I__577 (
            .O(N__5751),
            .I(\DUT.uart_inst0.recv_state_ns_0_0_0_cascade_ ));
    InMux I__576 (
            .O(N__5748),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_4 ));
    InMux I__575 (
            .O(N__5745),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_5 ));
    InMux I__574 (
            .O(N__5742),
            .I(N__5737));
    InMux I__573 (
            .O(N__5741),
            .I(N__5734));
    InMux I__572 (
            .O(N__5740),
            .I(N__5731));
    LocalMux I__571 (
            .O(N__5737),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_7 ));
    LocalMux I__570 (
            .O(N__5734),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_7 ));
    LocalMux I__569 (
            .O(N__5731),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_7 ));
    InMux I__568 (
            .O(N__5724),
            .I(N__5721));
    LocalMux I__567 (
            .O(N__5721),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO ));
    InMux I__566 (
            .O(N__5718),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_6 ));
    CascadeMux I__565 (
            .O(N__5715),
            .I(N__5711));
    InMux I__564 (
            .O(N__5714),
            .I(N__5707));
    InMux I__563 (
            .O(N__5711),
            .I(N__5704));
    InMux I__562 (
            .O(N__5710),
            .I(N__5701));
    LocalMux I__561 (
            .O(N__5707),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_8 ));
    LocalMux I__560 (
            .O(N__5704),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_8 ));
    LocalMux I__559 (
            .O(N__5701),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_8 ));
    InMux I__558 (
            .O(N__5694),
            .I(N__5691));
    LocalMux I__557 (
            .O(N__5691),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO ));
    InMux I__556 (
            .O(N__5688),
            .I(bfn_11_12_0_));
    InMux I__555 (
            .O(N__5685),
            .I(N__5680));
    InMux I__554 (
            .O(N__5684),
            .I(N__5677));
    InMux I__553 (
            .O(N__5683),
            .I(N__5674));
    LocalMux I__552 (
            .O(N__5680),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_9 ));
    LocalMux I__551 (
            .O(N__5677),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_9 ));
    LocalMux I__550 (
            .O(N__5674),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_9 ));
    InMux I__549 (
            .O(N__5667),
            .I(N__5664));
    LocalMux I__548 (
            .O(N__5664),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO ));
    InMux I__547 (
            .O(N__5661),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_8 ));
    CascadeMux I__546 (
            .O(N__5658),
            .I(N__5654));
    InMux I__545 (
            .O(N__5657),
            .I(N__5650));
    InMux I__544 (
            .O(N__5654),
            .I(N__5647));
    InMux I__543 (
            .O(N__5653),
            .I(N__5644));
    LocalMux I__542 (
            .O(N__5650),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_10 ));
    LocalMux I__541 (
            .O(N__5647),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_10 ));
    LocalMux I__540 (
            .O(N__5644),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_10 ));
    InMux I__539 (
            .O(N__5637),
            .I(N__5634));
    LocalMux I__538 (
            .O(N__5634),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO ));
    InMux I__537 (
            .O(N__5631),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_9 ));
    InMux I__536 (
            .O(N__5628),
            .I(N__5623));
    InMux I__535 (
            .O(N__5627),
            .I(N__5620));
    InMux I__534 (
            .O(N__5626),
            .I(N__5617));
    LocalMux I__533 (
            .O(N__5623),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_11 ));
    LocalMux I__532 (
            .O(N__5620),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_11 ));
    LocalMux I__531 (
            .O(N__5617),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_11 ));
    InMux I__530 (
            .O(N__5610),
            .I(N__5607));
    LocalMux I__529 (
            .O(N__5607),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO ));
    InMux I__528 (
            .O(N__5604),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_10 ));
    CascadeMux I__527 (
            .O(N__5601),
            .I(N__5596));
    CascadeMux I__526 (
            .O(N__5600),
            .I(N__5593));
    InMux I__525 (
            .O(N__5599),
            .I(N__5590));
    InMux I__524 (
            .O(N__5596),
            .I(N__5587));
    InMux I__523 (
            .O(N__5593),
            .I(N__5584));
    LocalMux I__522 (
            .O(N__5590),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_12 ));
    LocalMux I__521 (
            .O(N__5587),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_12 ));
    LocalMux I__520 (
            .O(N__5584),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_12 ));
    CascadeMux I__519 (
            .O(N__5577),
            .I(N__5574));
    InMux I__518 (
            .O(N__5574),
            .I(N__5571));
    LocalMux I__517 (
            .O(N__5571),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO ));
    InMux I__516 (
            .O(N__5568),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_11 ));
    CascadeMux I__515 (
            .O(N__5565),
            .I(\DUT.fifo_rx_inst.un1_i11_i_cascade_ ));
    InMux I__514 (
            .O(N__5562),
            .I(N__5559));
    LocalMux I__513 (
            .O(N__5559),
            .I(\DUT.fifo_rx_inst.un1_i11_i ));
    InMux I__512 (
            .O(N__5556),
            .I(N__5553));
    LocalMux I__511 (
            .O(N__5553),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO ));
    InMux I__510 (
            .O(N__5550),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_0 ));
    CascadeMux I__509 (
            .O(N__5547),
            .I(N__5544));
    InMux I__508 (
            .O(N__5544),
            .I(N__5541));
    LocalMux I__507 (
            .O(N__5541),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO ));
    InMux I__506 (
            .O(N__5538),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_1 ));
    InMux I__505 (
            .O(N__5535),
            .I(N__5532));
    LocalMux I__504 (
            .O(N__5532),
            .I(\DUT.uart_inst0.rx_clk_divider_1_3 ));
    InMux I__503 (
            .O(N__5529),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_2 ));
    InMux I__502 (
            .O(N__5526),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_3 ));
    InMux I__501 (
            .O(N__5523),
            .I(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0 ));
    InMux I__500 (
            .O(N__5520),
            .I(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1 ));
    CascadeMux I__499 (
            .O(N__5517),
            .I(\DUT.fifo_rx_inst.rFifoData_awe3_cascade_ ));
    IoInMux I__498 (
            .O(N__5514),
            .I(N__5511));
    LocalMux I__497 (
            .O(N__5511),
            .I(N__5508));
    Span12Mux_s3_v I__496 (
            .O(N__5508),
            .I(N__5505));
    Odrv12 I__495 (
            .O(N__5505),
            .I(wTxRdData_4));
    IoInMux I__494 (
            .O(N__5502),
            .I(N__5499));
    LocalMux I__493 (
            .O(N__5499),
            .I(N__5496));
    Span4Mux_s3_v I__492 (
            .O(N__5496),
            .I(N__5493));
    Span4Mux_v I__491 (
            .O(N__5493),
            .I(N__5490));
    Span4Mux_h I__490 (
            .O(N__5490),
            .I(N__5487));
    Odrv4 I__489 (
            .O(N__5487),
            .I(wTxRdData_1));
    InMux I__488 (
            .O(N__5484),
            .I(N__5481));
    LocalMux I__487 (
            .O(N__5481),
            .I(\PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO ));
    CascadeMux I__486 (
            .O(N__5478),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_3_cascade_ ));
    InMux I__485 (
            .O(N__5475),
            .I(N__5472));
    LocalMux I__484 (
            .O(N__5472),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_11 ));
    IoInMux I__483 (
            .O(N__5469),
            .I(N__5466));
    LocalMux I__482 (
            .O(N__5466),
            .I(N__5463));
    Sp12to4 I__481 (
            .O(N__5463),
            .I(N__5460));
    Span12Mux_v I__480 (
            .O(N__5460),
            .I(N__5457));
    Odrv12 I__479 (
            .O(N__5457),
            .I(wTxRdData_7));
    IoInMux I__478 (
            .O(N__5454),
            .I(N__5451));
    LocalMux I__477 (
            .O(N__5451),
            .I(N__5448));
    Span4Mux_s1_v I__476 (
            .O(N__5448),
            .I(N__5445));
    Span4Mux_v I__475 (
            .O(N__5445),
            .I(N__5442));
    Span4Mux_v I__474 (
            .O(N__5442),
            .I(N__5439));
    Span4Mux_h I__473 (
            .O(N__5439),
            .I(N__5436));
    Odrv4 I__472 (
            .O(N__5436),
            .I(wTxRdData_0));
    IoInMux I__471 (
            .O(N__5433),
            .I(N__5430));
    LocalMux I__470 (
            .O(N__5430),
            .I(N__5427));
    Span12Mux_s9_v I__469 (
            .O(N__5427),
            .I(N__5424));
    Span12Mux_v I__468 (
            .O(N__5424),
            .I(N__5421));
    Odrv12 I__467 (
            .O(N__5421),
            .I(BTN_N_c));
    IoInMux I__466 (
            .O(N__5418),
            .I(N__5415));
    LocalMux I__465 (
            .O(N__5415),
            .I(N__5412));
    Span4Mux_s1_v I__464 (
            .O(N__5412),
            .I(N__5409));
    Span4Mux_v I__463 (
            .O(N__5409),
            .I(N__5406));
    Span4Mux_v I__462 (
            .O(N__5406),
            .I(N__5403));
    Odrv4 I__461 (
            .O(N__5403),
            .I(wTxRdData_3));
    IoInMux I__460 (
            .O(N__5400),
            .I(N__5397));
    LocalMux I__459 (
            .O(N__5397),
            .I(N__5394));
    Span12Mux_s8_v I__458 (
            .O(N__5394),
            .I(N__5391));
    Odrv12 I__457 (
            .O(N__5391),
            .I(wTxRdData_5));
    IoInMux I__456 (
            .O(N__5388),
            .I(N__5385));
    LocalMux I__455 (
            .O(N__5385),
            .I(N__5382));
    Span4Mux_s1_v I__454 (
            .O(N__5382),
            .I(N__5379));
    Span4Mux_v I__453 (
            .O(N__5379),
            .I(N__5376));
    Span4Mux_v I__452 (
            .O(N__5376),
            .I(N__5373));
    Odrv4 I__451 (
            .O(N__5373),
            .I(wTxRdData_2));
    IoInMux I__450 (
            .O(N__5370),
            .I(N__5367));
    LocalMux I__449 (
            .O(N__5367),
            .I(N__5364));
    Span12Mux_s10_v I__448 (
            .O(N__5364),
            .I(N__5361));
    Odrv12 I__447 (
            .O(N__5361),
            .I(wTxRdData_6));
    defparam IN_MUX_bfv_17_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_12_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_12_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_14_0_));
    defparam IN_MUX_bfv_12_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_15_0_ (
            .carryinitin(\DUT.uart_inst0.tx_clk_divider_cry_7 ),
            .carryinitout(bfn_12_15_0_));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_11_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_12_0_ (
            .carryinitin(\DUT.uart_inst0.rx_clk_divider_1_cry_7 ),
            .carryinitout(bfn_11_12_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(\DUT.uart_inst0.rx_clk_divider_1_cry_15 ),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_20_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_17_0_));
    defparam IN_MUX_bfv_10_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_16_0_));
    ICE_GB wPllLocked_i_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__6486),
            .GLOBALBUFFEROUTPUT(wPllLocked_i_g));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB \top_pll_inst.top_pll_inst_RNISDA2  (
            .USERSIGNALTOGLOBALBUFFER(N__12454),
            .GLOBALBUFFEROUTPUT(wPllLocked_g));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0 .C_ON=1'b0;
    defparam \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0 .SEQ_MODE=4'b0000;
    defparam \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5484),
            .lcout(wPllLocked),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIL7JJ_7_LC_10_11_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIL7JJ_7_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIL7JJ_7_LC_10_11_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIL7JJ_7_LC_10_11_2  (
            .in0(_gnd_net_),
            .in1(N__5710),
            .in2(_gnd_net_),
            .in3(N__5740),
            .lcout(),
            .ltout(\DUT.uart_inst0.un2_rx_clk_divider_a_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIHKFQ1_5_LC_10_11_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIHKFQ1_5_LC_10_11_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIHKFQ1_5_LC_10_11_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIHKFQ1_5_LC_10_11_3  (
            .in0(N__6443),
            .in1(N__6470),
            .in2(N__5478),
            .in3(N__5475),
            .lcout(\DUT.uart_inst0.un2_rx_clk_divider_a_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIB99J_10_LC_10_11_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIB99J_10_LC_10_11_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIB99J_10_LC_10_11_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIB99J_10_LC_10_11_5  (
            .in0(N__5683),
            .in1(N__5626),
            .in2(N__5600),
            .in3(N__5653),
            .lcout(\DUT.uart_inst0.un2_rx_clk_divider_a_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_8_LC_10_12_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_8_LC_10_12_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_8_LC_10_12_1 .LUT_INIT=16'b1000110000100011;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_8_LC_10_12_1  (
            .in0(N__8319),
            .in1(N__5694),
            .in2(N__8120),
            .in3(N__5714),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13474),
            .ce(N__12011),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_12_LC_10_12_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_12_LC_10_12_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_12_LC_10_12_2 .LUT_INIT=16'b1011000000001011;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_12_LC_10_12_2  (
            .in0(N__8315),
            .in1(N__8078),
            .in2(N__5577),
            .in3(N__5599),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13474),
            .ce(N__12011),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_7_LC_10_12_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_7_LC_10_12_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_7_LC_10_12_3 .LUT_INIT=16'b1000101001000101;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_7_LC_10_12_3  (
            .in0(N__5724),
            .in1(N__8316),
            .in2(N__8121),
            .in3(N__5742),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13474),
            .ce(N__12011),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_9_LC_10_12_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_9_LC_10_12_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_9_LC_10_12_5 .LUT_INIT=16'b1000101001000101;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_9_LC_10_12_5  (
            .in0(N__5667),
            .in1(N__8317),
            .in2(N__8122),
            .in3(N__5685),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13474),
            .ce(N__12011),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_10_LC_10_12_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_10_LC_10_12_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_10_LC_10_12_6 .LUT_INIT=16'b1010001001010001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_10_LC_10_12_6  (
            .in0(N__5637),
            .in1(N__8077),
            .in2(N__8341),
            .in3(N__5657),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13474),
            .ce(N__12011),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_11_LC_10_12_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_11_LC_10_12_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_11_LC_10_12_7 .LUT_INIT=16'b1000110000100011;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_11_LC_10_12_7  (
            .in0(N__8318),
            .in1(N__5610),
            .in2(N__8119),
            .in3(N__5628),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13474),
            .ce(N__12011),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_5_LC_10_14_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_5_LC_10_14_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_5_LC_10_14_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \DUT.uart_inst0.recv_state_5_LC_10_14_7  (
            .in0(N__12296),
            .in1(N__5844),
            .in2(_gnd_net_),
            .in3(N__7365),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13463),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_LC_10_16_0 .C_ON=1'b1;
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_LC_10_16_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_LC_10_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_LC_10_16_0  (
            .in0(_gnd_net_),
            .in1(N__6053),
            .in2(N__5784),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_16_0_),
            .carryout(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_1_LC_10_16_1 .C_ON=1'b1;
    defparam \DUT.fifo_rx_inst.rFifoCount_1_LC_10_16_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoCount_1_LC_10_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_1_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(N__5810),
            .in2(N__5820),
            .in3(N__5523),
            .lcout(\DUT.fifo_rx_inst.rFifoCountZ0Z_1 ),
            .ltout(),
            .carryin(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0 ),
            .carryout(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1 ),
            .clk(N__13452),
            .ce(),
            .sr(N__13280));
    defparam \DUT.fifo_rx_inst.rFifoCount_2_LC_10_16_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_2_LC_10_16_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoCount_2_LC_10_16_2 .LUT_INIT=16'b0001111011100001;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_2_LC_10_16_2  (
            .in0(N__6027),
            .in1(N__6416),
            .in2(N__5985),
            .in3(N__5520),
            .lcout(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13452),
            .ce(),
            .sr(N__13280));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_2_1_LC_10_17_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_2_1_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_2_1_LC_10_17_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI96D91_2_1_LC_10_17_1  (
            .in0(N__6030),
            .in1(N__6351),
            .in2(N__6393),
            .in3(N__5981),
            .lcout(\DUT.fifo_rx_inst.rFifoData_awe3 ),
            .ltout(\DUT.fifo_rx_inst.rFifoData_awe3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1_1_LC_10_17_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1_1_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1_1_LC_10_17_2 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1_1_LC_10_17_2  (
            .in0(N__12188),
            .in1(_gnd_net_),
            .in2(N__5517),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.un1_i11_i ),
            .ltout(\DUT.fifo_rx_inst.un1_i11_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_0_LC_10_17_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_0_LC_10_17_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rWritePtr_0_LC_10_17_3 .LUT_INIT=16'b0000101000000101;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_0_LC_10_17_3  (
            .in0(N__6384),
            .in1(_gnd_net_),
            .in2(N__5565),
            .in3(N__6335),
            .lcout(\DUT.fifo_rx_inst.rWritePtrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13448),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_1_LC_10_17_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_1_LC_10_17_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rWritePtr_1_LC_10_17_6 .LUT_INIT=16'b0000000010110100;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_1_LC_10_17_6  (
            .in0(N__6336),
            .in1(N__6385),
            .in2(N__6363),
            .in3(N__5562),
            .lcout(\DUT.fifo_rx_inst.rWritePtrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13448),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_3_LC_11_10_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_3_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_3_LC_11_10_3 .LUT_INIT=16'b1110111111001111;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_3_LC_11_10_3  (
            .in0(N__6609),
            .in1(N__5535),
            .in2(N__7080),
            .in3(N__6522),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13481),
            .ce(N__12008),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_LC_11_10_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_1_LC_11_10_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_LC_11_10_6 .LUT_INIT=16'b1000110000100011;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_LC_11_10_6  (
            .in0(N__8278),
            .in1(N__5556),
            .in2(N__8140),
            .in3(N__5949),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13481),
            .ce(N__12008),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_2_LC_11_10_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_2_LC_11_10_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_2_LC_11_10_7 .LUT_INIT=16'b1000010010100101;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_2_LC_11_10_7  (
            .in0(N__5915),
            .in1(N__8279),
            .in2(N__5547),
            .in3(N__8114),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13481),
            .ce(N__12008),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_11_11_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_11_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5895),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_11_11_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_11_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(N__5948),
            .in2(N__8497),
            .in3(N__5550),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_0 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_11_11_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_11_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__8439),
            .in2(N__5919),
            .in3(N__5538),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_1 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_3_LC_11_11_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_3_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_3_LC_11_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNO_0_3_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(N__5931),
            .in2(N__8499),
            .in3(N__5529),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_3 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_2 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_11_11_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_11_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(N__8440),
            .in2(N__8010),
            .in3(N__5526),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_3 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_5_LC_11_11_5 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_5_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_5_LC_11_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNO_0_5_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(N__6471),
            .in2(N__8500),
            .in3(N__5748),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_5 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_4 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_6_LC_11_11_6 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_6_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_6_LC_11_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNO_0_6_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(N__8450),
            .in2(N__6447),
            .in3(N__5745),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_6 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_5 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_11_11_7 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_11_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(N__5741),
            .in2(N__8498),
            .in3(N__5718),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_6 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_11_12_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_11_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(N__8463),
            .in2(N__5715),
            .in3(N__5688),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_11_12_0_),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_11_12_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_11_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(N__5684),
            .in2(N__8504),
            .in3(N__5661),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_8 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_LUT4_0_LC_11_12_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_LUT4_0_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_LUT4_0_LC_11_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_LUT4_0_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(N__8467),
            .in2(N__5658),
            .in3(N__5631),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_9 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_LUT4_0_LC_11_12_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_LUT4_0_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_LUT4_0_LC_11_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_LUT4_0_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(N__5627),
            .in2(N__8501),
            .in3(N__5604),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_10 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_LUT4_0_LC_11_12_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_LUT4_0_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_LUT4_0_LC_11_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_LUT4_0_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(N__8455),
            .in2(N__5601),
            .in3(N__5568),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_11 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_LUT4_0_LC_11_12_5 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_LUT4_0_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_LUT4_0_LC_11_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_LUT4_0_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(N__6175),
            .in2(N__8502),
            .in3(N__5775),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_12 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_LUT4_0_LC_11_12_6 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_LUT4_0_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_LUT4_0_LC_11_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_LUT4_0_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(N__8459),
            .in2(N__6147),
            .in3(N__5772),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_13 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_LUT4_0_LC_11_12_7 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_LUT4_0_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_LUT4_0_LC_11_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_LUT4_0_LC_11_12_7  (
            .in0(_gnd_net_),
            .in1(N__6119),
            .in2(N__8503),
            .in3(N__5769),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_14 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_LUT4_0_LC_11_13_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_LUT4_0_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_LUT4_0_LC_11_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_LUT4_0_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__8468),
            .in2(N__6093),
            .in3(N__5766),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_17_LC_11_13_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_17_LC_11_13_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_17_LC_11_13_1 .LUT_INIT=16'b1011000000001011;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_17_LC_11_13_1  (
            .in0(N__8302),
            .in1(N__8070),
            .in2(N__5868),
            .in3(N__5763),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13464),
            .ce(N__12012),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNI237O_0_LC_11_14_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNI237O_0_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNI237O_0_LC_11_14_0 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \DUT.uart_inst0.recv_state_RNI237O_0_LC_11_14_0  (
            .in0(N__8329),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8040),
            .lcout(\DUT.uart_inst0.N_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_4_LC_11_14_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_4_LC_11_14_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_4_LC_11_14_1 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \DUT.uart_inst0.recv_state_4_LC_11_14_1  (
            .in0(N__12298),
            .in1(N__5760),
            .in2(N__7015),
            .in3(N__7349),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13457),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_0_LC_11_14_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_0_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_0_LC_11_14_4 .LUT_INIT=16'b0001010100010101;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_0_LC_11_14_4  (
            .in0(N__6026),
            .in1(N__8041),
            .in2(N__8349),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\DUT.uart_inst0.recv_state_ns_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_0_LC_11_14_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_0_LC_11_14_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_0_LC_11_14_5 .LUT_INIT=16'b0101111111011111;
    LogicCell40 \DUT.uart_inst0.recv_state_0_LC_11_14_5  (
            .in0(N__12297),
            .in1(N__5759),
            .in2(N__5751),
            .in3(N__7348),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13457),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_5_LC_11_15_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_5_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_5_LC_11_15_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_5_LC_11_15_2  (
            .in0(N__8334),
            .in1(N__5833),
            .in2(_gnd_net_),
            .in3(N__7406),
            .lcout(\DUT.uart_inst0.N_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_6_LC_11_15_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_6_LC_11_15_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_6_LC_11_15_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \DUT.uart_inst0.recv_state_6_LC_11_15_4  (
            .in0(N__8333),
            .in1(N__5835),
            .in2(N__12368),
            .in3(N__7358),
            .lcout(\DUT.wRcvd ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13453),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_3_LC_11_15_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_3_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_3_LC_11_15_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_3_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(N__7308),
            .in2(_gnd_net_),
            .in3(N__7427),
            .lcout(),
            .ltout(\DUT.uart_inst0.recv_state_srsts_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_3_LC_11_15_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_3_LC_11_15_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_3_LC_11_15_6 .LUT_INIT=16'b1000100000001010;
    LogicCell40 \DUT.uart_inst0.recv_state_3_LC_11_15_6  (
            .in0(N__12320),
            .in1(N__5834),
            .in2(N__5838),
            .in3(N__7359),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13453),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI9EGD1_0_LC_11_16_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI9EGD1_0_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI9EGD1_0_LC_11_16_0 .LUT_INIT=16'b0011001100110111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNI9EGD1_0_LC_11_16_0  (
            .in0(N__6051),
            .in1(N__13015),
            .in2(N__5811),
            .in3(N__5977),
            .lcout(\DUT.fifo_rx_inst.N_88 ),
            .ltout(\DUT.fifo_rx_inst.N_88_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIK3G92_1_LC_11_16_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIK3G92_1_LC_11_16_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIK3G92_1_LC_11_16_1 .LUT_INIT=16'b0000001100000011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNIK3G92_1_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(N__6025),
            .in2(N__5823),
            .in3(N__5809),
            .lcout(\DUT.fifo_rx_inst.rFifoCount_RNIK3G92Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_LC_11_16_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_LC_11_16_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_LC_11_16_5  (
            .in0(N__5976),
            .in1(N__5805),
            .in2(_gnd_net_),
            .in3(N__6050),
            .lcout(\DUT.fifo_rx_inst.rFifoCount_RNIHH0D1Z0Z_0 ),
            .ltout(\DUT.fifo_rx_inst.rFifoCount_RNIHH0D1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIPTFQ1_0_LC_11_16_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIPTFQ1_0_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIPTFQ1_0_LC_11_16_6 .LUT_INIT=16'b1111110000110011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNIPTFQ1_0_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__6023),
            .in2(N__5790),
            .in3(N__13016),
            .lcout(\DUT.fifo_rx_inst.N_97 ),
            .ltout(\DUT.fifo_rx_inst.N_97_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_11_16_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_11_16_7 .LUT_INIT=16'b0000011100000111;
    LogicCell40 \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_11_16_7  (
            .in0(N__5978),
            .in1(N__6024),
            .in2(N__5787),
            .in3(N__6052),
            .lcout(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_0_LC_11_17_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_0_LC_11_17_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoCount_0_LC_11_17_3 .LUT_INIT=16'b1110000110100101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_0_LC_11_17_3  (
            .in0(N__6063),
            .in1(N__6029),
            .in2(N__6057),
            .in3(N__5980),
            .lcout(\DUT.fifo_rx_inst.rFifoCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13443),
            .ce(),
            .sr(N__13278));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_11_17_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_11_17_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(N__6028),
            .in2(_gnd_net_),
            .in3(N__5979),
            .lcout(\DUT.fifo_rx_inst.N_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_0_LC_12_10_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_0_LC_12_10_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_0_LC_12_10_7 .LUT_INIT=16'b0000000010111011;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_0_LC_12_10_7  (
            .in0(N__8280),
            .in1(N__8115),
            .in2(_gnd_net_),
            .in3(N__5894),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13473),
            .ce(N__12007),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIMQ571_1_LC_12_11_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIMQ571_1_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIMQ571_1_LC_12_11_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIMQ571_1_LC_12_11_2  (
            .in0(N__5947),
            .in1(N__5930),
            .in2(N__8009),
            .in3(N__5911),
            .lcout(),
            .ltout(\DUT.uart_inst0.un2_rx_clk_divider_a_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIMSP02_16_LC_12_11_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIMSP02_16_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIMSP02_16_LC_12_11_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIMSP02_16_LC_12_11_3  (
            .in0(N__6088),
            .in1(N__5890),
            .in2(N__5874),
            .in3(N__5850),
            .lcout(\DUT.uart_inst0.un2_rx_clk_divider_a_15 ),
            .ltout(\DUT.uart_inst0.un2_rx_clk_divider_a_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_c_RNO_LC_12_11_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_c_RNO_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_c_RNO_LC_12_11_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_0_c_RNO_LC_12_11_4  (
            .in0(N__6763),
            .in1(_gnd_net_),
            .in2(N__5871),
            .in3(N__6523),
            .lcout(\DUT.uart_inst0.rx_countdown_3_cry_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNI3ALC_17_LC_12_11_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI3ALC_17_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI3ALC_17_LC_12_11_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNI3ALC_17_LC_12_11_5  (
            .in0(N__6142),
            .in1(N__6118),
            .in2(N__6177),
            .in3(N__5867),
            .lcout(\DUT.uart_inst0.un2_rx_clk_divider_a_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNICSMA4_1_LC_12_11_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNICSMA4_1_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNICSMA4_1_LC_12_11_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNICSMA4_1_LC_12_11_7  (
            .in0(N__6524),
            .in1(N__6729),
            .in2(N__6611),
            .in3(_gnd_net_),
            .lcout(\DUT.uart_inst0.rx_countdown_RNICSMA4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_1_LC_12_12_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_1_LC_12_12_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_1_LC_12_12_0 .LUT_INIT=16'b0111001101010000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_1_LC_12_12_0  (
            .in0(N__8286),
            .in1(N__7018),
            .in2(N__8147),
            .in3(N__6708),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13462),
            .ce(N__12009),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_5_LC_12_12_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_5_LC_12_12_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_5_LC_12_12_1 .LUT_INIT=16'b0100000001010000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_5_LC_12_12_1  (
            .in0(N__7016),
            .in1(N__8287),
            .in2(N__6651),
            .in3(N__8137),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13462),
            .ce(N__12009),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_0_LC_12_12_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_0_LC_12_12_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_0_LC_12_12_2 .LUT_INIT=16'b0010001100000000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_0_LC_12_12_2  (
            .in0(N__8285),
            .in1(N__7017),
            .in2(N__8146),
            .in3(N__6069),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13462),
            .ce(N__12009),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_13_LC_12_12_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_13_LC_12_12_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_13_LC_12_12_4 .LUT_INIT=16'b1000110000100011;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_13_LC_12_12_4  (
            .in0(N__8281),
            .in1(N__6183),
            .in2(N__8144),
            .in3(N__6176),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13462),
            .ce(N__12009),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_14_LC_12_12_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_14_LC_12_12_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_14_LC_12_12_5 .LUT_INIT=16'b1000010010100101;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_14_LC_12_12_5  (
            .in0(N__6146),
            .in1(N__8282),
            .in2(N__6156),
            .in3(N__8138),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13462),
            .ce(N__12009),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_15_LC_12_12_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_15_LC_12_12_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_15_LC_12_12_6 .LUT_INIT=16'b1000110000100011;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_15_LC_12_12_6  (
            .in0(N__8283),
            .in1(N__6126),
            .in2(N__8145),
            .in3(N__6120),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13462),
            .ce(N__12009),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_16_LC_12_12_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_16_LC_12_12_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_16_LC_12_12_7 .LUT_INIT=16'b1000010010100101;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_16_LC_12_12_7  (
            .in0(N__6092),
            .in1(N__8284),
            .in2(N__6102),
            .in3(N__8139),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13462),
            .ce(N__12009),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_12_13_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_12_13_0 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_12_13_0  (
            .in0(N__8301),
            .in1(N__7390),
            .in2(_gnd_net_),
            .in3(N__7306),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_46_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_12_13_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_12_13_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_12_13_1  (
            .in0(N__6944),
            .in1(N__6923),
            .in2(N__6072),
            .in3(N__6899),
            .lcout(\DUT.uart_inst0.N_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_0_LC_12_13_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_0_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_0_LC_12_13_2 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_0_0_LC_12_13_2  (
            .in0(N__6615),
            .in1(_gnd_net_),
            .in2(N__6765),
            .in3(N__6549),
            .lcout(\DUT.uart_inst0.rx_countdown_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNI8KQG9_0_LC_12_13_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNI8KQG9_0_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNI8KQG9_0_LC_12_13_4 .LUT_INIT=16'b1101111011111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNI8KQG9_0_LC_12_13_4  (
            .in0(N__6614),
            .in1(N__6707),
            .in2(N__6764),
            .in3(N__6548),
            .lcout(),
            .ltout(\DUT.uart_inst0.rx_countdown_RNI8KQG9Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNI8EL7E_0_LC_12_13_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNI8EL7E_0_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNI8EL7E_0_LC_12_13_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNI8EL7E_0_LC_12_13_5  (
            .in0(N__6644),
            .in1(_gnd_net_),
            .in2(N__6204),
            .in3(N__8451),
            .lcout(\DUT.uart_inst0.rx_countdown_8_i_o2_2_2 ),
            .ltout(\DUT.uart_inst0.rx_countdown_8_i_o2_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_c_RNIHH7QT_LC_12_13_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_c_RNIHH7QT_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_c_RNIHH7QT_LC_12_13_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_1_c_RNIHH7QT_LC_12_13_6  (
            .in0(N__6922),
            .in1(N__6966),
            .in2(N__6201),
            .in3(N__6943),
            .lcout(\DUT.uart_inst0.N_42 ),
            .ltout(\DUT.uart_inst0.N_42_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_1_LC_12_13_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_1_LC_12_13_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_1_LC_12_13_7 .LUT_INIT=16'b1000000011001100;
    LogicCell40 \DUT.uart_inst0.recv_state_1_LC_12_13_7  (
            .in0(N__7391),
            .in1(N__12366),
            .in2(N__6198),
            .in3(N__7057),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13456),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_12_14_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_12_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7134),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_14_0_),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_1_LC_12_14_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_1_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_1_LC_12_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_1_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__7149),
            .in2(N__8532),
            .in3(N__6195),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_1 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_0 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_1 ),
            .clk(N__13451),
            .ce(),
            .sr(N__7107));
    defparam \DUT.uart_inst0.tx_clk_divider_2_LC_12_14_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_2_LC_12_14_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_2_LC_12_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_2_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(N__8508),
            .in2(N__6783),
            .in3(N__6192),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_2 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_1 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_2 ),
            .clk(N__13451),
            .ce(),
            .sr(N__7107));
    defparam \DUT.uart_inst0.tx_clk_divider_3_LC_12_14_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_3_LC_12_14_3 .SEQ_MODE=4'b1001;
    defparam \DUT.uart_inst0.tx_clk_divider_3_LC_12_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_3_LC_12_14_3  (
            .in0(_gnd_net_),
            .in1(N__6813),
            .in2(N__8533),
            .in3(N__6189),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_3 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_2 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_3 ),
            .clk(N__13451),
            .ce(),
            .sr(N__7107));
    defparam \DUT.uart_inst0.tx_clk_divider_4_LC_12_14_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_4_LC_12_14_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_4_LC_12_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_4_LC_12_14_4  (
            .in0(_gnd_net_),
            .in1(N__8512),
            .in2(N__6828),
            .in3(N__6186),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_4 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_3 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_4 ),
            .clk(N__13451),
            .ce(),
            .sr(N__7107));
    defparam \DUT.uart_inst0.tx_clk_divider_5_LC_12_14_5 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_5_LC_12_14_5 .SEQ_MODE=4'b1001;
    defparam \DUT.uart_inst0.tx_clk_divider_5_LC_12_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_5_LC_12_14_5  (
            .in0(_gnd_net_),
            .in1(N__6797),
            .in2(N__8534),
            .in3(N__6231),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_5 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_4 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_5 ),
            .clk(N__13451),
            .ce(),
            .sr(N__7107));
    defparam \DUT.uart_inst0.tx_clk_divider_6_LC_12_14_6 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_6_LC_12_14_6 .SEQ_MODE=4'b1001;
    defparam \DUT.uart_inst0.tx_clk_divider_6_LC_12_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_6_LC_12_14_6  (
            .in0(_gnd_net_),
            .in1(N__8516),
            .in2(N__6846),
            .in3(N__6228),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_6 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_5 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_6 ),
            .clk(N__13451),
            .ce(),
            .sr(N__7107));
    defparam \DUT.uart_inst0.tx_clk_divider_7_LC_12_14_7 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_7_LC_12_14_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_7_LC_12_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_7_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(N__6876),
            .in2(N__8535),
            .in3(N__6225),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_7 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_6 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_7 ),
            .clk(N__13451),
            .ce(),
            .sr(N__7107));
    defparam \DUT.uart_inst0.tx_clk_divider_8_LC_12_15_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_8_LC_12_15_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_8_LC_12_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_8_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(N__7161),
            .in2(N__8538),
            .in3(N__6222),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_8 ),
            .ltout(),
            .carryin(bfn_12_15_0_),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_8 ),
            .clk(N__13447),
            .ce(),
            .sr(N__7106));
    defparam \DUT.uart_inst0.tx_clk_divider_9_LC_12_15_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_9_LC_12_15_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_9_LC_12_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_9_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(N__8531),
            .in2(N__7176),
            .in3(N__6219),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_9 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_8 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_9 ),
            .clk(N__13447),
            .ce(),
            .sr(N__7106));
    defparam \DUT.uart_inst0.tx_clk_divider_10_LC_12_15_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_10_LC_12_15_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_10_LC_12_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_10_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(N__7188),
            .in2(N__8536),
            .in3(N__6216),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_10 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_9 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_10 ),
            .clk(N__13447),
            .ce(),
            .sr(N__7106));
    defparam \DUT.uart_inst0.tx_clk_divider_11_LC_12_15_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_11_LC_12_15_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_11_LC_12_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_11_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(N__8524),
            .in2(N__7203),
            .in3(N__6213),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_11 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_10 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_11 ),
            .clk(N__13447),
            .ce(),
            .sr(N__7106));
    defparam \DUT.uart_inst0.tx_clk_divider_12_LC_12_15_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_12_LC_12_15_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_12_LC_12_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_12_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(N__6888),
            .in2(N__8537),
            .in3(N__6210),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_12 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_11 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_12 ),
            .clk(N__13447),
            .ce(),
            .sr(N__7106));
    defparam \DUT.uart_inst0.tx_clk_divider_13_LC_12_15_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_13_LC_12_15_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_13_LC_12_15_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_13_LC_12_15_5  (
            .in0(_gnd_net_),
            .in1(N__6860),
            .in2(_gnd_net_),
            .in3(N__6207),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13447),
            .ce(),
            .sr(N__7106));
    defparam \DUT.uart_inst0.tx_clk_divider_0_LC_12_15_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_0_LC_12_15_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_0_LC_12_15_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_0_LC_12_15_6  (
            .in0(N__8520),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7133),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13447),
            .ce(),
            .sr(N__7106));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIUJI11_3_LC_12_16_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIUJI11_3_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIUJI11_3_LC_12_16_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNIUJI11_3_LC_12_16_0  (
            .in0(N__6243),
            .in1(N__6305),
            .in2(N__6267),
            .in3(N__7454),
            .lcout(\DUT.uart_inst0.N_62_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_3_LC_12_16_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_3_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_3_LC_12_16_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_1_3_LC_12_16_1  (
            .in0(N__7455),
            .in1(N__7286),
            .in2(N__6314),
            .in3(N__6244),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_3_LC_12_16_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_3_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_3_LC_12_16_2 .LUT_INIT=16'b0110010100100001;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_0_3_LC_12_16_2  (
            .in0(N__6265),
            .in1(N__7413),
            .in2(N__6273),
            .in3(N__7242),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_3_LC_12_16_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_3_LC_12_16_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_bits_remaining_3_LC_12_16_3 .LUT_INIT=16'b1011111100000100;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_3_LC_12_16_3  (
            .in0(N__7362),
            .in1(N__12326),
            .in2(N__6270),
            .in3(N__6266),
            .lcout(\DUT.uart_inst0.rx_bits_remainingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13442),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_1_LC_12_16_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_1_LC_12_16_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_bits_remaining_1_LC_12_16_4 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_1_LC_12_16_4  (
            .in0(N__12324),
            .in1(N__7360),
            .in2(N__6285),
            .in3(N__6312),
            .lcout(\DUT.uart_inst0.rx_bits_remainingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13442),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_2_LC_12_16_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_2_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_2_LC_12_16_5 .LUT_INIT=16'b0000010011111011;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_1_2_LC_12_16_5  (
            .in0(N__7456),
            .in1(N__7287),
            .in2(N__6315),
            .in3(N__6245),
            .lcout(),
            .ltout(\DUT.uart_inst0.m5_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_2_LC_12_16_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_2_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_2_LC_12_16_6 .LUT_INIT=16'b0000010000001111;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_0_2_LC_12_16_6  (
            .in0(N__7288),
            .in1(N__8336),
            .in2(N__6252),
            .in3(N__7412),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_2_LC_12_16_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_2_LC_12_16_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_bits_remaining_2_LC_12_16_7 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_2_LC_12_16_7  (
            .in0(N__7361),
            .in1(N__12325),
            .in2(N__6249),
            .in3(N__6246),
            .lcout(\DUT.uart_inst0.rx_bits_remainingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13442),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rReadPtr_1_LC_12_17_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rReadPtr_1_LC_12_17_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rReadPtr_1_LC_12_17_0 .LUT_INIT=16'b0100000101000100;
    LogicCell40 \DUT.fifo_rx_inst.rReadPtr_1_LC_12_17_0  (
            .in0(N__6426),
            .in1(N__9912),
            .in2(N__6417),
            .in3(N__9398),
            .lcout(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13439),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_12_17_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_12_17_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_12_17_1  (
            .in0(N__6394),
            .in1(N__6364),
            .in2(_gnd_net_),
            .in3(N__6332),
            .lcout(\DUT.fifo_rx_inst.rFifoData_awe1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rReadPtr_RNI4NC92_0_LC_12_17_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rReadPtr_RNI4NC92_0_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rReadPtr_RNI4NC92_0_LC_12_17_2 .LUT_INIT=16'b0100111100001111;
    LogicCell40 \DUT.fifo_rx_inst.rReadPtr_RNI4NC92_0_LC_12_17_2  (
            .in0(N__6411),
            .in1(N__9911),
            .in2(N__12192),
            .in3(N__9396),
            .lcout(\DUT.fifo_rx_inst.un1_i11_2_i ),
            .ltout(\DUT.fifo_rx_inst.un1_i11_2_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rReadPtr_0_LC_12_17_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rReadPtr_0_LC_12_17_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rReadPtr_0_LC_12_17_3 .LUT_INIT=16'b0000101000000101;
    LogicCell40 \DUT.fifo_rx_inst.rReadPtr_0_LC_12_17_3  (
            .in0(N__9397),
            .in1(_gnd_net_),
            .in2(N__6420),
            .in3(N__6412),
            .lcout(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13439),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_12_17_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_12_17_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_12_17_4  (
            .in0(N__6333),
            .in1(N__6395),
            .in2(_gnd_net_),
            .in3(N__6366),
            .lcout(\DUT.fifo_rx_inst.rFifoData_awe0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_12_17_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_12_17_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_12_17_5  (
            .in0(N__6396),
            .in1(N__6365),
            .in2(_gnd_net_),
            .in3(N__6334),
            .lcout(\DUT.fifo_rx_inst.rFifoData_awe2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_1_LC_12_17_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_1_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_1_LC_12_17_6 .LUT_INIT=16'b0011001110011001;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_1_1_LC_12_17_6  (
            .in0(N__7284),
            .in1(N__6313),
            .in2(_gnd_net_),
            .in3(N__7453),
            .lcout(),
            .ltout(\DUT.uart_inst0.m5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_1_LC_12_17_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_1_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_1_LC_12_17_7 .LUT_INIT=16'b0000001100001011;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_0_1_LC_12_17_7  (
            .in0(N__8335),
            .in1(N__7414),
            .in2(N__6288),
            .in3(N__7285),
            .lcout(\DUT.uart_inst0.N_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_12_18_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_12_18_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_12_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_12_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10187),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13436),
            .ce(N__10013),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_12_18_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_12_18_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_12_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_12_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9717),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13436),
            .ce(N__10013),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_12_18_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_12_18_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_12_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_12_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10118),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13436),
            .ce(N__10013),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_4_LC_12_19_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_4_LC_12_19_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_4_LC_12_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_4_LC_12_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10222),
            .lcout(\DUT.wRxByte_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13434),
            .ce(N__7499),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_7_LC_12_19_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_7_LC_12_19_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_7_LC_12_19_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.uart_inst0.rx_data_7_LC_12_19_5  (
            .in0(N__8350),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.wRxByte_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13434),
            .ce(N__7499),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_0_LC_12_20_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_0_LC_12_20_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_0_LC_12_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_0_LC_12_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9704),
            .lcout(\DUT.wRxByte_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13433),
            .ce(N__7500),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.wPllLocked_i_LC_12_30_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.wPllLocked_i_LC_12_30_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.wPllLocked_i_LC_12_30_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \DUT.uart_inst0.wPllLocked_i_LC_12_30_4  (
            .in0(N__12191),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(wPllLocked_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_5_LC_13_11_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_5_LC_13_11_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_5_LC_13_11_0 .LUT_INIT=16'b1110111110101111;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_5_LC_13_11_0  (
            .in0(N__6480),
            .in1(N__6596),
            .in2(N__7086),
            .in3(N__6551),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13475),
            .ce(N__12010),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_6_LC_13_11_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_6_LC_13_11_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_6_LC_13_11_1 .LUT_INIT=16'b1110110011111111;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_6_LC_13_11_1  (
            .in0(N__6552),
            .in1(N__6456),
            .in2(N__6612),
            .in3(N__7085),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13475),
            .ce(N__12010),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNIEUMA4_3_LC_13_11_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNIEUMA4_3_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNIEUMA4_3_LC_13_11_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNIEUMA4_3_LC_13_11_2  (
            .in0(N__6690),
            .in1(N__6595),
            .in2(_gnd_net_),
            .in3(N__6550),
            .lcout(\DUT.uart_inst0.rx_countdown_RNIEUMA4Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_LC_13_11_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_LC_13_11_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_3_LC_13_11_6 .LUT_INIT=16'b1010100011111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_LC_13_11_6  (
            .in0(N__8320),
            .in1(N__7027),
            .in2(N__6951),
            .in3(N__8124),
            .lcout(\DUT.uart_inst0.rx_countdownZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13475),
            .ce(N__12010),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_4_LC_13_11_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_4_LC_13_11_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_4_LC_13_11_7 .LUT_INIT=16'b0000110100000000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_4_LC_13_11_7  (
            .in0(N__8123),
            .in1(N__8321),
            .in2(N__7034),
            .in3(N__6924),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13475),
            .ce(N__12010),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_c_LC_13_12_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_c_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_c_LC_13_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_0_c_LC_13_12_0  (
            .in0(_gnd_net_),
            .in1(N__6756),
            .in2(N__6738),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_c_RNITO365_LC_13_12_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_c_RNITO365_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_c_RNITO365_LC_13_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_0_c_RNITO365_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__6728),
            .in2(N__6717),
            .in3(N__6696),
            .lcout(\DUT.uart_inst0.rx_countdown_3_1 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_countdown_3_cry_0 ),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_c_RNI0T465_LC_13_12_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_c_RNI0T465_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_c_RNI0T465_LC_13_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_1_c_RNI0T465_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(N__6492),
            .in2(N__6981),
            .in3(N__6693),
            .lcout(\DUT.uart_inst0.rx_countdown_3_2 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_countdown_3_cry_1 ),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_2_c_RNI31665_LC_13_12_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_2_c_RNI31665_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_2_c_RNI31665_LC_13_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_2_c_RNI31665_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(N__6689),
            .in2(N__6678),
            .in3(N__6666),
            .lcout(\DUT.uart_inst0.rx_countdown_3_3 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_countdown_3_cry_2 ),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_c_RNI65765_LC_13_12_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_c_RNI65765_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_c_RNI65765_LC_13_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_3_c_RNI65765_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(N__6621),
            .in2(N__6633),
            .in3(N__6663),
            .lcout(\DUT.uart_inst0.rx_countdown_3_4 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_countdown_3_cry_3 ),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_4_c_RNI0QQM4_LC_13_12_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_4_c_RNI0QQM4_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_4_c_RNI0QQM4_LC_13_12_5 .LUT_INIT=16'b1001001101101100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_4_c_RNI0QQM4_LC_13_12_5  (
            .in0(N__6547),
            .in1(N__6660),
            .in2(N__6613),
            .in3(N__6654),
            .lcout(\DUT.uart_inst0.rx_countdown_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNIFVMA4_4_LC_13_12_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNIFVMA4_4_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNIFVMA4_4_LC_13_12_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNIFVMA4_4_LC_13_12_6  (
            .in0(N__6632),
            .in1(N__6600),
            .in2(_gnd_net_),
            .in3(N__6546),
            .lcout(\DUT.uart_inst0.rx_countdown_RNIFVMA4Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNIDTMA4_2_LC_13_13_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNIDTMA4_2_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNIDTMA4_2_LC_13_13_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNIDTMA4_2_LC_13_13_0  (
            .in0(N__6980),
            .in1(N__6610),
            .in2(_gnd_net_),
            .in3(N__6545),
            .lcout(\DUT.uart_inst0.rx_countdown_RNIDTMA4Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_2_LC_13_13_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_2_LC_13_13_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_2_LC_13_13_4 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_2_LC_13_13_4  (
            .in0(N__7081),
            .in1(N__7041),
            .in2(N__7035),
            .in3(N__6965),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13465),
            .ce(N__12013),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_c_RNI93IIF_LC_13_13_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_c_RNI93IIF_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_c_RNI93IIF_LC_13_13_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_1_c_RNI93IIF_LC_13_13_5  (
            .in0(N__6964),
            .in1(N__6942),
            .in2(_gnd_net_),
            .in3(N__6921),
            .lcout(),
            .ltout(\DUT.uart_inst0.rx_bits_remaining_2_sqmuxa_0_a2_0_a2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNIPAH9U_2_LC_13_13_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNIPAH9U_2_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNIPAH9U_2_LC_13_13_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNIPAH9U_2_LC_13_13_6  (
            .in0(N__7307),
            .in1(N__12367),
            .in2(N__6903),
            .in3(N__6900),
            .lcout(\DUT.uart_inst0.rx_bits_remaining_2_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_5_LC_13_14_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_5_LC_13_14_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_5_LC_13_14_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_5_LC_13_14_0  (
            .in0(N__10536),
            .in1(N__8748),
            .in2(_gnd_net_),
            .in3(N__9302),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13458),
            .ce(N__12021),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_13_LC_13_14_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_13_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_13_LC_13_14_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_13_LC_13_14_1  (
            .in0(N__6887),
            .in1(N__6875),
            .in2(N__6864),
            .in3(N__6842),
            .lcout(\DUT.uart_inst0.un1_tx_clk_divider_8 ),
            .ltout(\DUT.uart_inst0.un1_tx_clk_divider_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNI7N692_4_LC_13_14_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNI7N692_4_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNI7N692_4_LC_13_14_2 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNI7N692_4_LC_13_14_2  (
            .in0(N__7548),
            .in1(N__7719),
            .in2(N__6831),
            .in3(N__7805),
            .lcout(\DUT.uart_inst0.tx_countdown_RNI7N692Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_RNI2V95_2_LC_13_14_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI2V95_2_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI2V95_2_LC_13_14_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNI2V95_2_LC_13_14_5  (
            .in0(N__6824),
            .in1(N__6812),
            .in2(N__6801),
            .in3(N__6779),
            .lcout(\DUT.uart_inst0.un1_tx_clk_divider_9 ),
            .ltout(\DUT.uart_inst0.un1_tx_clk_divider_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNI3J692_0_LC_13_14_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNI3J692_0_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNI3J692_0_LC_13_14_6 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNI3J692_0_LC_13_14_6  (
            .in0(N__7612),
            .in1(N__7755),
            .in2(N__6768),
            .in3(N__7806),
            .lcout(\DUT.uart_inst0.tx_countdown_3_0 ),
            .ltout(\DUT.uart_inst0.tx_countdown_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_0_LC_13_14_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_0_LC_13_14_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_0_LC_13_14_7 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_0_LC_13_14_7  (
            .in0(N__9301),
            .in1(_gnd_net_),
            .in2(N__7206),
            .in3(N__10537),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13458),
            .ce(N__12021),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_RNIR5NO_9_LC_13_15_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNIR5NO_9_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNIR5NO_9_LC_13_15_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNIR5NO_9_LC_13_15_1  (
            .in0(N__7199),
            .in1(N__7187),
            .in2(_gnd_net_),
            .in3(N__7172),
            .lcout(),
            .ltout(\DUT.uart_inst0.un1_tx_clk_divider_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_RNIJJMS_0_LC_13_15_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNIJJMS_0_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNIJJMS_0_LC_13_15_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNIJJMS_0_LC_13_15_2  (
            .in0(N__7160),
            .in1(N__7148),
            .in2(N__7137),
            .in3(N__7129),
            .lcout(\DUT.uart_inst0.un1_tx_clk_divider_10 ),
            .ltout(\DUT.uart_inst0.un1_tx_clk_divider_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNI5L692_2_LC_13_15_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNI5L692_2_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNI5L692_2_LC_13_15_3 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNI5L692_2_LC_13_15_3  (
            .in0(N__7747),
            .in1(N__7584),
            .in2(N__7113),
            .in3(N__7714),
            .lcout(\DUT.uart_inst0.tx_countdown_RNI5L692Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNI8CH01_0_LC_13_15_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNI8CH01_0_LC_13_15_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNI8CH01_0_LC_13_15_4 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \DUT.uart_inst0.tx_state_RNI8CH01_0_LC_13_15_4  (
            .in0(N__12166),
            .in1(N__10538),
            .in2(_gnd_net_),
            .in3(N__9306),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_clk_divider_1_sqmuxa_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNI5PJS2_0_LC_13_15_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNI5PJS2_0_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNI5PJS2_0_LC_13_15_5 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \DUT.uart_inst0.tx_state_RNI5PJS2_0_LC_13_15_5  (
            .in0(N__7802),
            .in1(N__7761),
            .in2(N__7110),
            .in3(N__7716),
            .lcout(\DUT.uart_inst0.tx_clk_divider_1_sqmuxa_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_3_cry_0_c_RNO_LC_13_15_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_3_cry_0_c_RNO_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_3_cry_0_c_RNO_LC_13_15_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_3_cry_0_c_RNO_LC_13_15_6  (
            .in0(N__7713),
            .in1(N__7746),
            .in2(N__7617),
            .in3(N__7800),
            .lcout(\DUT.uart_inst0.tx_countdown_3_cry_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNI8O692_5_LC_13_15_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNI8O692_5_LC_13_15_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNI8O692_5_LC_13_15_7 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNI8O692_5_LC_13_15_7  (
            .in0(N__7801),
            .in1(N__7095),
            .in2(N__7759),
            .in3(N__7715),
            .lcout(\DUT.uart_inst0.tx_countdown_3_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_0_LC_13_16_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_0_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_0_LC_13_16_1 .LUT_INIT=16'b0101000100100010;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_0_0_LC_13_16_1  (
            .in0(N__7281),
            .in1(N__7415),
            .in2(N__8352),
            .in3(N__7457),
            .lcout(),
            .ltout(\DUT.uart_inst0.g0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_0_LC_13_16_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_0_LC_13_16_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_bits_remaining_0_LC_13_16_2 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_0_LC_13_16_2  (
            .in0(N__12313),
            .in1(N__7458),
            .in2(N__7461),
            .in3(N__7364),
            .lcout(\DUT.uart_inst0.rx_bits_remainingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13449),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_2_LC_13_16_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_2_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_2_LC_13_16_3 .LUT_INIT=16'b0010111100100010;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_2_LC_13_16_3  (
            .in0(N__7282),
            .in1(N__7428),
            .in2(N__8351),
            .in3(N__7416),
            .lcout(),
            .ltout(\DUT.uart_inst0.recv_state_srsts_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_2_LC_13_16_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_2_LC_13_16_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_2_LC_13_16_4 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \DUT.uart_inst0.recv_state_2_LC_13_16_4  (
            .in0(N__12312),
            .in1(N__7283),
            .in2(N__7368),
            .in3(N__7363),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13449),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_2_3_LC_13_16_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_2_3_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_2_3_LC_13_16_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_2_3_LC_13_16_6  (
            .in0(_gnd_net_),
            .in1(N__8348),
            .in2(_gnd_net_),
            .in3(N__7280),
            .lcout(\DUT.uart_inst0.m5_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNI0AQO1_LC_13_17_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNI0AQO1_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNI0AQO1_LC_13_17_0 .LUT_INIT=16'b1111001011110111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_0_RNI0AQO1_LC_13_17_0  (
            .in0(N__9381),
            .in1(N__7226),
            .in2(N__9913),
            .in3(N__7235),
            .lcout(\DUT.fifo_rx_inst.rTxByte_52_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_LC_13_17_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_LC_13_17_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_LC_13_17_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_0_LC_13_17_1  (
            .in0(N__7236),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9988),
            .lcout(\DUT.fifo_rx_inst.rFifoDataro_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13444),
            .ce(),
            .sr(N__13279));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_1_LC_13_17_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_1_LC_13_17_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_1_LC_13_17_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_1_LC_13_17_2  (
            .in0(_gnd_net_),
            .in1(N__7958),
            .in2(_gnd_net_),
            .in3(N__7227),
            .lcout(\DUT.fifo_rx_inst.rFifoDataro_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13444),
            .ce(),
            .sr(N__13279));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_13_18_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_13_18_2 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_13_18_2  (
            .in0(N__7218),
            .in1(N__9908),
            .in2(N__7860),
            .in3(N__9394),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_13_18_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_13_18_3 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_13_18_3  (
            .in0(N__9393),
            .in1(N__7212),
            .in2(N__7974),
            .in3(N__9910),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_13_18_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_13_18_4 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_13_18_4  (
            .in0(N__7506),
            .in1(N__9909),
            .in2(N__7983),
            .in3(N__9395),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_13_19_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_13_19_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_13_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_13_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10220),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13437),
            .ce(N__10012),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_13_19_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_13_19_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_13_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_13_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9606),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13437),
            .ce(N__10012),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_13_19_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_13_19_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_13_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_13_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10263),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13437),
            .ce(N__10012),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_13_19_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_13_19_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_13_19_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_13_19_7  (
            .in0(_gnd_net_),
            .in1(N__9649),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13437),
            .ce(N__10012),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_2_LC_13_20_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_2_LC_13_20_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_2_LC_13_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_2_LC_13_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9605),
            .lcout(\DUT.wRxByte_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13435),
            .ce(N__7495),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_3_LC_13_20_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_3_LC_13_20_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_3_LC_13_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_3_LC_13_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10264),
            .lcout(\DUT.wRxByte_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13435),
            .ce(N__7495),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_1_LC_13_20_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_1_LC_13_20_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_1_LC_13_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_1_LC_13_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9648),
            .lcout(\DUT.wRxByte_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13435),
            .ce(N__7495),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_5_LC_13_20_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_5_LC_13_20_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_5_LC_13_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_5_LC_13_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10169),
            .lcout(\DUT.wRxByte_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13435),
            .ce(N__7495),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_6_LC_13_20_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_6_LC_13_20_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_6_LC_13_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_6_LC_13_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10119),
            .lcout(\DUT.wRxByte_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13435),
            .ce(N__7495),
            .sr(_gnd_net_));
    defparam \DUT.rTransmit_LC_14_11_5 .C_ON=1'b0;
    defparam \DUT.rTransmit_LC_14_11_5 .SEQ_MODE=4'b1000;
    defparam \DUT.rTransmit_LC_14_11_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \DUT.rTransmit_LC_14_11_5  (
            .in0(N__13119),
            .in1(N__10499),
            .in2(_gnd_net_),
            .in3(N__8692),
            .lcout(\DUT.rTransmitZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13482),
            .ce(),
            .sr(N__13286));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI5UON8_3_LC_14_12_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI5UON8_3_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI5UON8_3_LC_14_12_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNI5UON8_3_LC_14_12_0  (
            .in0(N__9182),
            .in1(N__8908),
            .in2(N__8754),
            .in3(N__8793),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_bits_remaining_RNI5UON8Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNIVQ9CI_0_LC_14_12_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNIVQ9CI_0_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNIVQ9CI_0_LC_14_12_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \DUT.uart_inst0.tx_state_RNIVQ9CI_0_LC_14_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7527),
            .in3(N__7512),
            .lcout(\DUT.uart_inst0.N_109 ),
            .ltout(\DUT.uart_inst0.N_109_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_1_LC_14_12_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_1_LC_14_12_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_state_1_LC_14_12_2 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \DUT.uart_inst0.tx_state_1_LC_14_12_2  (
            .in0(N__8690),
            .in1(N__7634),
            .in2(N__7524),
            .in3(N__8953),
            .lcout(\DUT.tx_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13476),
            .ce(),
            .sr(N__13285));
    defparam \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIKK41C_LC_14_12_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIKK41C_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIKK41C_LC_14_12_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIKK41C_LC_14_12_3  (
            .in0(N__8831),
            .in1(N__8749),
            .in2(N__8910),
            .in3(N__8870),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIKK41CZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNIN7BAE_0_LC_14_12_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNIN7BAE_0_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNIN7BAE_0_LC_14_12_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNIN7BAE_0_LC_14_12_4  (
            .in0(_gnd_net_),
            .in1(N__8435),
            .in2(N__7521),
            .in3(N__8794),
            .lcout(\DUT.uart_inst0.N_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_0_LC_14_12_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_0_LC_14_12_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_state_0_LC_14_12_5 .LUT_INIT=16'b0000000000110010;
    LogicCell40 \DUT.uart_inst0.tx_state_0_LC_14_12_5  (
            .in0(N__10490),
            .in1(N__8691),
            .in2(N__13078),
            .in3(N__7518),
            .lcout(\DUT.tx_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13476),
            .ce(),
            .sr(N__13285));
    defparam \DUT.uart_inst0.tx_state_RNIQSGK9_0_LC_14_12_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNIQSGK9_0_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNIQSGK9_0_LC_14_12_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \DUT.uart_inst0.tx_state_RNIQSGK9_0_LC_14_12_6  (
            .in0(N__8869),
            .in1(N__8952),
            .in2(N__10509),
            .in3(N__8830),
            .lcout(\DUT.uart_inst0.tx_state_ns_i_i_a3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_1_LC_14_13_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_1_LC_14_13_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_1_LC_14_13_1 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_1_LC_14_13_1  (
            .in0(N__10491),
            .in1(N__9298),
            .in2(_gnd_net_),
            .in3(N__8867),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13470),
            .ce(N__12022),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_4_LC_14_13_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_4_LC_14_13_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_4_LC_14_13_2 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_4_LC_14_13_2  (
            .in0(N__10498),
            .in1(N__9297),
            .in2(_gnd_net_),
            .in3(N__8904),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13470),
            .ce(N__12022),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_3_LC_14_13_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_3_LC_14_13_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_3_LC_14_13_3 .LUT_INIT=16'b1111111011001100;
    LogicCell40 \DUT.uart_inst0.tx_countdown_3_LC_14_13_3  (
            .in0(N__9296),
            .in1(N__8979),
            .in2(N__10535),
            .in3(N__8829),
            .lcout(\DUT.uart_inst0.tx_countdownZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13470),
            .ce(N__12022),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_2_LC_14_13_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_2_LC_14_13_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_2_LC_14_13_5 .LUT_INIT=16'b1111111100010101;
    LogicCell40 \DUT.uart_inst0.tx_countdown_2_LC_14_13_5  (
            .in0(N__9107),
            .in1(N__7635),
            .in2(N__10534),
            .in3(N__8950),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13470),
            .ce(N__12022),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNISDA2_0_LC_14_13_6 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNISDA2_0_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNISDA2_0_LC_14_13_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNISDA2_0_LC_14_13_6  (
            .in0(N__11889),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12165),
            .lcout(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_3_cry_0_c_LC_14_14_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_countdown_3_cry_0_c_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_3_cry_0_c_LC_14_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_3_cry_0_c_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(N__7623),
            .in2(N__7616),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(\DUT.uart_inst0.tx_countdown_3_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_3_cry_0_c_RNIPMF33_LC_14_14_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_countdown_3_cry_0_c_RNIPMF33_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_3_cry_0_c_RNIPMF33_LC_14_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_countdown_3_cry_0_c_RNIPMF33_LC_14_14_1  (
            .in0(_gnd_net_),
            .in1(N__7812),
            .in2(N__7833),
            .in3(N__7593),
            .lcout(\DUT.uart_inst0.tx_countdown_3_1 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_countdown_3_cry_0 ),
            .carryout(\DUT.uart_inst0.tx_countdown_3_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_3_cry_1_c_RNISQG33_LC_14_14_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_countdown_3_cry_1_c_RNISQG33_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_3_cry_1_c_RNISQG33_LC_14_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_countdown_3_cry_1_c_RNISQG33_LC_14_14_2  (
            .in0(_gnd_net_),
            .in1(N__7590),
            .in2(N__7583),
            .in3(N__7560),
            .lcout(\DUT.uart_inst0.tx_countdown_3_2 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_countdown_3_cry_1 ),
            .carryout(\DUT.uart_inst0.tx_countdown_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIVUH33_LC_14_14_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIVUH33_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIVUH33_LC_14_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIVUH33_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__7689),
            .in2(N__7776),
            .in3(N__7557),
            .lcout(\DUT.uart_inst0.tx_countdown_3_3 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_countdown_3_cry_2 ),
            .carryout(\DUT.uart_inst0.tx_countdown_3_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_3_cry_3_c_RNI23J33_LC_14_14_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_countdown_3_cry_3_c_RNI23J33_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_3_cry_3_c_RNI23J33_LC_14_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_countdown_3_cry_3_c_RNI23J33_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(N__7554),
            .in2(N__7547),
            .in3(N__7530),
            .lcout(\DUT.uart_inst0.tx_countdown_3_4 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_countdown_3_cry_3 ),
            .carryout(\DUT.uart_inst0.tx_countdown_3_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_3_cry_4_c_RNIQRFM2_LC_14_14_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_3_cry_4_c_RNIQRFM2_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_3_cry_4_c_RNIQRFM2_LC_14_14_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \DUT.uart_inst0.tx_countdown_3_cry_4_c_RNIQRFM2_LC_14_14_5  (
            .in0(N__7842),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7836),
            .lcout(\DUT.uart_inst0.tx_countdown_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNI4K692_1_LC_14_14_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNI4K692_1_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNI4K692_1_LC_14_14_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNI4K692_1_LC_14_14_6  (
            .in0(N__7717),
            .in1(N__7751),
            .in2(N__7832),
            .in3(N__7803),
            .lcout(\DUT.uart_inst0.tx_countdown_RNI4K692Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNI6M692_3_LC_14_14_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNI6M692_3_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNI6M692_3_LC_14_14_7 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNI6M692_3_LC_14_14_7  (
            .in0(N__7804),
            .in1(N__7775),
            .in2(N__7760),
            .in3(N__7718),
            .lcout(\DUT.uart_inst0.tx_countdown_RNI6M692Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.un1_tx_bits_remaining_cry_0_c_LC_14_15_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.un1_tx_bits_remaining_cry_0_c_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.un1_tx_bits_remaining_cry_0_c_LC_14_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.uart_inst0.un1_tx_bits_remaining_cry_0_c_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__8700),
            .in2(N__9219),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\DUT.uart_inst0.un1_tx_bits_remaining_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_1_LC_14_15_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_bits_remaining_1_LC_14_15_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_bits_remaining_1_LC_14_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_1_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(N__9246),
            .in2(N__9240),
            .in3(N__7683),
            .lcout(\DUT.uart_inst0.tx_bits_remainingZ0Z_1 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.un1_tx_bits_remaining_cry_0 ),
            .carryout(\DUT.uart_inst0.un1_tx_bits_remaining_cry_1 ),
            .clk(N__13459),
            .ce(),
            .sr(N__8973));
    defparam \DUT.uart_inst0.tx_bits_remaining_2_LC_14_15_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_bits_remaining_2_LC_14_15_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_bits_remaining_2_LC_14_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_2_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__9126),
            .in2(N__9144),
            .in3(N__7680),
            .lcout(\DUT.uart_inst0.tx_bits_remainingZ0Z_2 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.un1_tx_bits_remaining_cry_1 ),
            .carryout(\DUT.uart_inst0.un1_tx_bits_remaining_cry_2 ),
            .clk(N__13459),
            .ce(),
            .sr(N__8973));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_14_15_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_14_15_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_14_15_3  (
            .in0(_gnd_net_),
            .in1(N__9036),
            .in2(_gnd_net_),
            .in3(N__7677),
            .lcout(\DUT.uart_inst0.tx_bits_remaining_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ft2232h_inst.rRx_n_LC_14_16_0 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rRx_n_LC_14_16_0 .SEQ_MODE=4'b1001;
    defparam \fifo_inst.ft2232h_inst.rRx_n_LC_14_16_0 .LUT_INIT=16'b1100111010101110;
    LogicCell40 \fifo_inst.ft2232h_inst.rRx_n_LC_14_16_0  (
            .in0(N__9555),
            .in1(N__7646),
            .in2(N__9531),
            .in3(N__9460),
            .lcout(P1A3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13454),
            .ce(),
            .sr(N__13281));
    defparam rRxRead_LC_14_16_1.C_ON=1'b0;
    defparam rRxRead_LC_14_16_1.SEQ_MODE=4'b1000;
    defparam rRxRead_LC_14_16_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 rRxRead_LC_14_16_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7891),
            .lcout(rRxReadZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13454),
            .ce(),
            .sr(N__13281));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_LC_14_16_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_LC_14_16_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_LC_14_16_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_0_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(N__11078),
            .in2(_gnd_net_),
            .in3(N__13173),
            .lcout(\DUT.fifo_tx_inst.rFifoDataro_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13454),
            .ce(),
            .sr(N__13281));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI250E6_0_LC_14_17_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI250E6_0_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI250E6_0_LC_14_17_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNI250E6_0_LC_14_17_0  (
            .in0(_gnd_net_),
            .in1(N__9814),
            .in2(_gnd_net_),
            .in3(N__7908),
            .lcout(N_100_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_0_LC_14_17_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_0_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_0_LC_14_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_0_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7892),
            .lcout(N_100_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_14_17_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_14_17_2 .LUT_INIT=16'b0101111100111111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_14_17_2  (
            .in0(N__9578),
            .in1(N__9542),
            .in2(N__9945),
            .in3(N__9399),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rTxByte_52_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNIHJV05_LC_14_17_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNIHJV05_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNIHJV05_LC_14_17_3 .LUT_INIT=16'b0101010111010101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_0_RNIHJV05_LC_14_17_3  (
            .in0(N__12187),
            .in1(N__7902),
            .in2(N__7896),
            .in3(N__7893),
            .lcout(rFifoDatarff_0_RNIHJV05),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_14_17_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_14_17_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_14_17_7 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_14_17_7  (
            .in0(N__9400),
            .in1(N__7851),
            .in2(N__7872),
            .in3(N__9917),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_14_18_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_14_18_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_14_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10054),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13445),
            .ce(N__7965),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_14_18_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_14_18_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_14_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9718),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13445),
            .ce(N__7965),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_14_18_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_14_18_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_14_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9658),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13445),
            .ce(N__7965),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_14_18_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_14_18_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_14_18_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_14_18_3  (
            .in0(N__9614),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13445),
            .ce(N__7965),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_14_18_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_14_18_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_14_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10280),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13445),
            .ce(N__7965),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_14_18_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_14_18_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_14_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10229),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13445),
            .ce(N__7965),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_14_18_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_14_18_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_14_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_14_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10183),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13445),
            .ce(N__7965),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_14_18_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_14_18_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_14_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_14_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10136),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13445),
            .ce(N__7965),
            .sr(_gnd_net_));
    defparam rTxByte_esr_5_LC_14_19_0.C_ON=1'b0;
    defparam rTxByte_esr_5_LC_14_19_0.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_5_LC_14_19_0.LUT_INIT=16'b1010000011001111;
    LogicCell40 rTxByte_esr_5_LC_14_19_0 (
            .in0(N__10194),
            .in1(N__8547),
            .in2(N__9964),
            .in3(N__7914),
            .lcout(rTxByteZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13440),
            .ce(N__9849),
            .sr(N__9828));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_14_19_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_14_19_1 .LUT_INIT=16'b0011010000110111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_14_19_1  (
            .in0(N__7947),
            .in1(N__9413),
            .in2(N__9966),
            .in3(N__7938),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rTxByte_esr_4_LC_14_19_2.C_ON=1'b0;
    defparam rTxByte_esr_4_LC_14_19_2.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_4_LC_14_19_2.LUT_INIT=16'b1100101100001011;
    LogicCell40 rTxByte_esr_4_LC_14_19_2 (
            .in0(N__9780),
            .in1(N__9958),
            .in2(N__7932),
            .in3(N__10242),
            .lcout(rTxByteZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13440),
            .ce(N__9849),
            .sr(N__9828));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_14_19_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_14_19_3 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_14_19_3  (
            .in0(N__7929),
            .in1(N__9946),
            .in2(N__7923),
            .in3(N__9411),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_14_19_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_14_19_4 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_14_19_4  (
            .in0(N__9412),
            .in1(N__9954),
            .in2(N__8586),
            .in3(N__8577),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rTxByte_esr_3_LC_14_19_5.C_ON=1'b0;
    defparam rTxByte_esr_3_LC_14_19_5.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_3_LC_14_19_5.LUT_INIT=16'b1100101000001111;
    LogicCell40 rTxByte_esr_3_LC_14_19_5 (
            .in0(N__8556),
            .in1(N__10287),
            .in2(N__8571),
            .in3(N__9953),
            .lcout(rTxByteZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13440),
            .ce(N__9849),
            .sr(N__9828));
    defparam rTxByte_esr_6_LC_14_19_6.C_ON=1'b0;
    defparam rTxByte_esr_6_LC_14_19_6.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_6_LC_14_19_6.LUT_INIT=16'b1010000011001111;
    LogicCell40 rTxByte_esr_6_LC_14_19_6 (
            .in0(N__10143),
            .in1(N__8562),
            .in2(N__9965),
            .in3(N__8568),
            .lcout(rTxByteZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13440),
            .ce(N__9849),
            .sr(N__9828));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_14_20_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_14_20_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_14_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10137),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13438),
            .ce(N__9773),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_14_20_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_14_20_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_14_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_14_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10170),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13438),
            .ce(N__9773),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_14_20_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_14_20_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_14_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_14_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9607),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13438),
            .ce(N__9773),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_14_20_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_14_20_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_14_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_14_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10221),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13438),
            .ce(N__9773),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_15_9_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_15_9_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_15_9_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_15_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_4_LC_15_11_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_4_LC_15_11_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_4_LC_15_11_0 .LUT_INIT=16'b1000110000100011;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_4_LC_15_11_0  (
            .in0(N__8340),
            .in1(N__8160),
            .in2(N__8148),
            .in3(N__8002),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13486),
            .ce(N__12014),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_LC_15_11_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_LC_15_11_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_out_LC_15_11_1 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \DUT.uart_inst0.tx_out_LC_15_11_1  (
            .in0(N__8604),
            .in1(N__8592),
            .in2(N__8627),
            .in3(N__9069),
            .lcout(P1A7_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13486),
            .ce(N__12014),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIFI07_LC_15_11_2 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIFI07_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIFI07_LC_15_11_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIFI07_LC_15_11_2  (
            .in0(N__11628),
            .in1(N__12161),
            .in2(_gnd_net_),
            .in3(N__10797),
            .lcout(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_3 ),
            .ltout(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIFI07_2_LC_15_11_3 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIFI07_2_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIFI07_2_LC_15_11_3 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIFI07_2_LC_15_11_3  (
            .in0(N__11753),
            .in1(_gnd_net_),
            .in2(N__8643),
            .in3(N__10961),
            .lcout(\fifo_inst.tx_fifo_inst.un18_rRamWrAddr_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNIPNAVK_0_LC_15_12_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNIPNAVK_0_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNIPNAVK_0_LC_15_12_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \DUT.uart_inst0.tx_state_RNIPNAVK_0_LC_15_12_0  (
            .in0(N__12424),
            .in1(N__9108),
            .in2(_gnd_net_),
            .in3(N__9068),
            .lcout(\DUT.uart_inst0.N_71_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_RNO_0_LC_15_12_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_RNO_0_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_out_RNO_0_LC_15_12_1 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \DUT.uart_inst0.tx_out_RNO_0_LC_15_12_1  (
            .in0(N__8689),
            .in1(N__8620),
            .in2(N__9183),
            .in3(N__10316),
            .lcout(\DUT.uart_inst0.N_112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_RNO_3_LC_15_12_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_RNO_3_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_out_RNO_3_LC_15_12_2 .LUT_INIT=16'b0000000010101000;
    LogicCell40 \DUT.uart_inst0.tx_out_RNO_3_LC_15_12_2  (
            .in0(N__10468),
            .in1(N__9178),
            .in2(N__10317),
            .in3(N__8688),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_out_6_iv_0_a3_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_RNO_2_LC_15_12_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_RNO_2_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_out_RNO_2_LC_15_12_3 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \DUT.uart_inst0.tx_out_RNO_2_LC_15_12_3  (
            .in0(N__8832),
            .in1(N__8954),
            .in2(N__8598),
            .in3(N__8871),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_out_6_iv_0_a3_1_sx_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_RNO_1_LC_15_12_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_RNO_1_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_out_RNO_1_LC_15_12_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_out_RNO_1_LC_15_12_4  (
            .in0(N__8798),
            .in1(N__8753),
            .in2(N__8595),
            .in3(N__8909),
            .lcout(\DUT.uart_inst0.N_113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_0_LC_15_13_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_0_LC_15_13_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_bits_remaining_0_LC_15_13_4 .LUT_INIT=16'b1100110010011100;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_0_LC_15_13_4  (
            .in0(N__9106),
            .in1(N__9210),
            .in2(N__12455),
            .in3(N__9067),
            .lcout(\DUT.uart_inst0.tx_bits_remainingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13477),
            .ce(),
            .sr(N__8972));
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_15_13_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_15_13_6 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_15_13_6  (
            .in0(N__9177),
            .in1(N__8866),
            .in2(N__8955),
            .in3(N__10475),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_countdown_7_i_a3_0_sx_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_15_13_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_15_13_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_15_13_7  (
            .in0(N__8799),
            .in1(N__8747),
            .in2(N__8982),
            .in3(N__8903),
            .lcout(\DUT.uart_inst0.N_116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNI8CH01_0_0_LC_15_14_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNI8CH01_0_0_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNI8CH01_0_0_LC_15_14_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \DUT.uart_inst0.tx_state_RNI8CH01_0_0_LC_15_14_0  (
            .in0(N__10503),
            .in1(N__12175),
            .in2(_gnd_net_),
            .in3(N__9300),
            .lcout(\DUT.uart_inst0.N_76_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIMJ5EC_LC_15_14_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIMJ5EC_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIMJ5EC_LC_15_14_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIMJ5EC_LC_15_14_2  (
            .in0(N__8951),
            .in1(N__8894),
            .in2(N__8868),
            .in3(N__8820),
            .lcout(\DUT.uart_inst0.tx_countdown_3_cry_2_c_RNIMJ5ECZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNI6I8K_1_LC_15_14_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNI6I8K_1_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNI6I8K_1_LC_15_14_3 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \DUT.uart_inst0.tx_state_RNI6I8K_1_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(N__8693),
            .in2(_gnd_net_),
            .in3(N__13052),
            .lcout(\DUT.uart_inst0.N_77 ),
            .ltout(\DUT.uart_inst0.N_77_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNI9DTT5_0_LC_15_14_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNI9DTT5_0_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNI9DTT5_0_LC_15_14_4 .LUT_INIT=16'b1111101011011000;
    LogicCell40 \DUT.uart_inst0.tx_state_RNI9DTT5_0_LC_15_14_4  (
            .in0(N__10500),
            .in1(N__8789),
            .in2(N__8757),
            .in3(N__8738),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_state_RNI9DTT5Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNIBV9AJ_0_LC_15_14_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNIBV9AJ_0_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNIBV9AJ_0_LC_15_14_5 .LUT_INIT=16'b1111000011101110;
    LogicCell40 \DUT.uart_inst0.tx_state_RNIBV9AJ_0_LC_15_14_5  (
            .in0(N__9299),
            .in1(N__10501),
            .in2(N__8712),
            .in3(N__8709),
            .lcout(\DUT.uart_inst0.N_99 ),
            .ltout(\DUT.uart_inst0.N_99_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.un1_tx_bits_remaining_cry_0_c_RNO_LC_15_14_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.un1_tx_bits_remaining_cry_0_c_RNO_LC_15_14_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.un1_tx_bits_remaining_cry_0_c_RNO_LC_15_14_6 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \DUT.uart_inst0.un1_tx_bits_remaining_cry_0_c_RNO_LC_15_14_6  (
            .in0(N__9211),
            .in1(N__12381),
            .in2(N__8703),
            .in3(N__9099),
            .lcout(\DUT.uart_inst0.un1_tx_bits_remaining_cry_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNIIAMI1_1_LC_15_14_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNIIAMI1_1_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNIIAMI1_1_LC_15_14_7 .LUT_INIT=16'b1110111011001111;
    LogicCell40 \DUT.uart_inst0.tx_state_RNIIAMI1_1_LC_15_14_7  (
            .in0(N__9173),
            .in1(N__8694),
            .in2(N__13065),
            .in3(N__10502),
            .lcout(\DUT.uart_inst0.N_96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_3_LC_15_15_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_3_LC_15_15_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_bits_remaining_3_LC_15_15_0 .LUT_INIT=16'b1111111100010000;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_3_LC_15_15_0  (
            .in0(N__9295),
            .in1(N__10539),
            .in2(N__12417),
            .in3(N__9252),
            .lcout(\DUT.uart_inst0.tx_bits_remainingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13466),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNIAIE4L_1_LC_15_15_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNIAIE4L_1_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNIAIE4L_1_LC_15_15_1 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNIAIE4L_1_LC_15_15_1  (
            .in0(N__9239),
            .in1(N__9100),
            .in2(N__12418),
            .in3(N__9058),
            .lcout(\DUT.uart_inst0.tx_bits_remaining_RNIAIE4LZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_3_LC_15_15_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_3_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_3_LC_15_15_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_3_LC_15_15_3  (
            .in0(N__9139),
            .in1(N__9235),
            .in2(N__9120),
            .in3(N__9212),
            .lcout(\DUT.uart_inst0.N_124 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ft2232h_inst.rFifoState_RNIRPB71_0_LC_15_15_4 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rFifoState_RNIRPB71_0_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ft2232h_inst.rFifoState_RNIRPB71_0_LC_15_15_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \fifo_inst.ft2232h_inst.rFifoState_RNIRPB71_0_LC_15_15_4  (
            .in0(N__9461),
            .in1(N__9502),
            .in2(_gnd_net_),
            .in3(N__9524),
            .lcout(\fifo_inst.ft2232h_inst.rFifoStatec_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNIBJE4L_2_LC_15_15_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNIBJE4L_2_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNIBJE4L_2_LC_15_15_5 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNIBJE4L_2_LC_15_15_5  (
            .in0(N__9140),
            .in1(N__9101),
            .in2(N__12419),
            .in3(N__9059),
            .lcout(\DUT.uart_inst0.tx_bits_remaining_RNIBJE4LZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ft2232h_inst.rFifoState_RNO_0_0_LC_15_15_6 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rFifoState_RNO_0_0_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ft2232h_inst.rFifoState_RNO_0_0_LC_15_15_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \fifo_inst.ft2232h_inst.rFifoState_RNO_0_0_LC_15_15_6  (
            .in0(N__9462),
            .in1(N__9503),
            .in2(_gnd_net_),
            .in3(N__9525),
            .lcout(\fifo_inst.ft2232h_inst.N_103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_1_3_LC_15_15_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_1_3_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_1_3_LC_15_15_7 .LUT_INIT=16'b1010101010011010;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNO_1_3_LC_15_15_7  (
            .in0(N__9119),
            .in1(N__9102),
            .in2(N__12420),
            .in3(N__9060),
            .lcout(\DUT.uart_inst0.un1_tx_bits_remaining_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ft2232h_inst.rFifoState_1_LC_15_16_0 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rFifoState_1_LC_15_16_0 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rFifoState_1_LC_15_16_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_inst.ft2232h_inst.rFifoState_1_LC_15_16_0  (
            .in0(N__9453),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9527),
            .lcout(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13460),
            .ce(),
            .sr(N__13282));
    defparam \fifo_inst.ft2232h_inst.rTx_n_LC_15_16_1 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rTx_n_LC_15_16_1 .SEQ_MODE=4'b1001;
    defparam \fifo_inst.ft2232h_inst.rTx_n_LC_15_16_1 .LUT_INIT=16'b1100000011101010;
    LogicCell40 \fifo_inst.ft2232h_inst.rTx_n_LC_15_16_1  (
            .in0(N__8998),
            .in1(N__13920),
            .in2(N__13872),
            .in3(N__12959),
            .lcout(P1A4_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13460),
            .ce(),
            .sr(N__13282));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_3_LC_15_16_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_3_LC_15_16_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_3_LC_15_16_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_3_LC_15_16_2  (
            .in0(_gnd_net_),
            .in1(N__9774),
            .in2(_gnd_net_),
            .in3(N__9579),
            .lcout(\DUT.fifo_rx_inst.rFifoDataro_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13460),
            .ce(),
            .sr(N__13282));
    defparam \fifo_inst.ft2232h_inst.rFifoState_2_LC_15_16_4 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rFifoState_2_LC_15_16_4 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rFifoState_2_LC_15_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.ft2232h_inst.rFifoState_2_LC_15_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9567),
            .lcout(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13460),
            .ce(),
            .sr(N__13282));
    defparam \fifo_inst.ft2232h_inst.rFifoState_0_LC_15_16_5 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rFifoState_0_LC_15_16_5 .SEQ_MODE=4'b1001;
    defparam \fifo_inst.ft2232h_inst.rFifoState_0_LC_15_16_5 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \fifo_inst.ft2232h_inst.rFifoState_0_LC_15_16_5  (
            .in0(N__9561),
            .in1(N__13919),
            .in2(N__13871),
            .in3(N__9554),
            .lcout(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13460),
            .ce(),
            .sr(N__13282));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_LC_15_16_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_LC_15_16_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_LC_15_16_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_2_LC_15_16_6  (
            .in0(_gnd_net_),
            .in1(N__10082),
            .in2(_gnd_net_),
            .in3(N__9543),
            .lcout(\DUT.fifo_rx_inst.rFifoDataro_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13460),
            .ce(),
            .sr(N__13282));
    defparam \fifo_inst.ft2232h_inst.rFifoState_3_LC_15_16_7 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rFifoState_3_LC_15_16_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rFifoState_3_LC_15_16_7 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \fifo_inst.ft2232h_inst.rFifoState_3_LC_15_16_7  (
            .in0(N__9526),
            .in1(N__9504),
            .in2(_gnd_net_),
            .in3(N__9454),
            .lcout(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13460),
            .ce(),
            .sr(N__13282));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_15_17_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_15_17_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_15_17_0  (
            .in0(N__10023),
            .in1(N__9959),
            .in2(N__9423),
            .in3(N__9414),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rTxByte_esr_0_LC_15_17_1.C_ON=1'b0;
    defparam rTxByte_esr_0_LC_15_17_1.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_0_LC_15_17_1.LUT_INIT=16'b1010110100001101;
    LogicCell40 rTxByte_esr_0_LC_15_17_1 (
            .in0(N__9960),
            .in1(N__9792),
            .in2(N__9348),
            .in3(N__9735),
            .lcout(rTxByteZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13455),
            .ce(N__9845),
            .sr(N__9827));
    defparam rTxByte_esr_7_LC_15_17_2.C_ON=1'b0;
    defparam rTxByte_esr_7_LC_15_17_2.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_7_LC_15_17_2.LUT_INIT=16'b1000111110000011;
    LogicCell40 rTxByte_esr_7_LC_15_17_2 (
            .in0(N__10092),
            .in1(N__9963),
            .in2(N__9345),
            .in3(N__9330),
            .lcout(rTxByteZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13455),
            .ce(N__9845),
            .sr(N__9827));
    defparam rTxByte_esr_1_LC_15_17_4.C_ON=1'b0;
    defparam rTxByte_esr_1_LC_15_17_4.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_1_LC_15_17_4.LUT_INIT=16'b1100000010111011;
    LogicCell40 rTxByte_esr_1_LC_15_17_4 (
            .in0(N__9798),
            .in1(N__9961),
            .in2(N__9678),
            .in3(N__9318),
            .lcout(rTxByteZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13455),
            .ce(N__9845),
            .sr(N__9827));
    defparam rTxByte_esr_2_LC_15_17_6.C_ON=1'b0;
    defparam rTxByte_esr_2_LC_15_17_6.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_2_LC_15_17_6.LUT_INIT=16'b1000111110000011;
    LogicCell40 rTxByte_esr_2_LC_15_17_6 (
            .in0(N__9627),
            .in1(N__9962),
            .in2(N__9858),
            .in3(N__9786),
            .lcout(rTxByteZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13455),
            .ce(N__9845),
            .sr(N__9827));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_15_18_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_15_18_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_15_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_15_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9726),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13450),
            .ce(N__9772),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_15_18_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_15_18_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_15_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_15_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10058),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13450),
            .ce(N__9772),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_15_18_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_15_18_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_15_18_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(N__9666),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13450),
            .ce(N__9772),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_15_18_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_15_18_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_15_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_15_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10281),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13450),
            .ce(N__9772),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_15_19_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_15_19_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_15_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_15_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10059),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13446),
            .ce(N__10083),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_15_19_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_15_19_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_15_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_15_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9725),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13446),
            .ce(N__10083),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_15_19_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_15_19_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_15_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_15_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9665),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13446),
            .ce(N__10083),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_15_19_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_15_19_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_15_19_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_15_19_3  (
            .in0(N__9618),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13446),
            .ce(N__10083),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_15_19_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_15_19_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_15_19_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_15_19_4  (
            .in0(N__10273),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13446),
            .ce(N__10083),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_15_19_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_15_19_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_15_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_15_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10233),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13446),
            .ce(N__10083),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_15_19_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_15_19_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_15_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_15_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10188),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13446),
            .ce(N__10083),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_15_19_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_15_19_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_15_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_15_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10129),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13446),
            .ce(N__10083),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_15_20_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_15_20_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_15_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_15_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10044),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13441),
            .ce(N__10014),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIGLV01_2_LC_16_10_0 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIGLV01_2_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIGLV01_2_LC_16_10_0 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIGLV01_2_LC_16_10_0  (
            .in0(N__9972),
            .in1(N__11577),
            .in2(N__12476),
            .in3(N__10742),
            .lcout(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_2_LC_16_10_1 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_2_LC_16_10_1 .SEQ_MODE=4'b1010;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_2_LC_16_10_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_2_LC_16_10_1  (
            .in0(N__10743),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12160),
            .lcout(\fifo_inst.tx_fifo_inst.rRamRdAddr_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13491),
            .ce(N__11288),
            .sr(N__13289));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_1_LC_16_10_2 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_1_LC_16_10_2 .SEQ_MODE=4'b1010;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_1_LC_16_10_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_1_LC_16_10_2  (
            .in0(N__12159),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10359),
            .lcout(\fifo_inst.tx_fifo_inst.rRamRdAddr_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13491),
            .ce(N__11288),
            .sr(N__13289));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIFI07_0_LC_16_11_2 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIFI07_0_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIFI07_0_LC_16_11_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIFI07_0_LC_16_11_2  (
            .in0(N__10790),
            .in1(N__12164),
            .in2(_gnd_net_),
            .in3(N__11627),
            .lcout(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_0_1_LC_16_11_4 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_0_1_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_0_1_LC_16_11_4 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_0_1_LC_16_11_4  (
            .in0(N__10346),
            .in1(N__11575),
            .in2(N__12456),
            .in3(N__10358),
            .lcout(\fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_1_1 ),
            .ltout(\fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNI_1_LC_16_11_5 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNI_1_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNI_1_LC_16_11_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_RNI_1_LC_16_11_5  (
            .in0(N__11476),
            .in1(_gnd_net_),
            .in2(N__10362),
            .in3(_gnd_net_),
            .lcout(\fifo_inst.tx_fifo_inst.rRamRdAddr_RNIZ0Z_1 ),
            .ltout(\fifo_inst.tx_fifo_inst.rRamRdAddr_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_1_LC_16_11_6 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_1_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_1_LC_16_11_6 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_1_LC_16_11_6  (
            .in0(N__10347),
            .in1(N__12428),
            .in2(N__10338),
            .in3(N__11576),
            .lcout(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_1 ),
            .ltout(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_2_1_LC_16_11_7 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_2_1_LC_16_11_7 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_2_1_LC_16_11_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_2_1_LC_16_11_7  (
            .in0(N__11660),
            .in1(N__10762),
            .in2(N__10320),
            .in3(N__10724),
            .lcout(\fifo_inst.tx_fifo_inst.un15_rRamRdAddr_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_0_LC_16_12_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_0_LC_16_12_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_0_LC_16_12_0 .LUT_INIT=16'b1100110000001010;
    LogicCell40 \DUT.uart_inst0.tx_data_0_LC_16_12_0  (
            .in0(N__11016),
            .in1(N__10305),
            .in2(N__11061),
            .in3(N__10533),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13487),
            .ce(N__10376),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_3_LC_16_12_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_3_LC_16_12_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_3_LC_16_12_1 .LUT_INIT=16'b1010000010101100;
    LogicCell40 \DUT.uart_inst0.tx_data_3_LC_16_12_1  (
            .in0(N__10569),
            .in1(N__10926),
            .in2(N__10547),
            .in3(N__11060),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13487),
            .ce(N__10376),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_1_LC_16_12_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_1_LC_16_12_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_1_LC_16_12_2 .LUT_INIT=16'b1101110000010000;
    LogicCell40 \DUT.uart_inst0.tx_data_1_LC_16_12_2  (
            .in0(N__11055),
            .in1(N__10526),
            .in2(N__11094),
            .in3(N__10293),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13487),
            .ce(N__10376),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_2_LC_16_12_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_2_LC_16_12_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_2_LC_16_12_3 .LUT_INIT=16'b1010000010101100;
    LogicCell40 \DUT.uart_inst0.tx_data_2_LC_16_12_3  (
            .in0(N__10299),
            .in1(N__12648),
            .in2(N__10546),
            .in3(N__11059),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13487),
            .ce(N__10376),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_7_LC_16_13_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_7_LC_16_13_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_7_LC_16_13_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \DUT.uart_inst0.tx_data_7_LC_16_13_2  (
            .in0(N__11052),
            .in1(N__10908),
            .in2(_gnd_net_),
            .in3(N__10545),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13483),
            .ce(N__10383),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_4_LC_16_13_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_4_LC_16_13_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_4_LC_16_13_3 .LUT_INIT=16'b1010101000110000;
    LogicCell40 \DUT.uart_inst0.tx_data_4_LC_16_13_3  (
            .in0(N__10389),
            .in1(N__11053),
            .in2(N__10623),
            .in3(N__10543),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13483),
            .ce(N__10383),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_6_LC_16_13_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_6_LC_16_13_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_6_LC_16_13_4 .LUT_INIT=16'b1111010000000100;
    LogicCell40 \DUT.uart_inst0.tx_data_6_LC_16_13_4  (
            .in0(N__11051),
            .in1(N__10599),
            .in2(N__10548),
            .in3(N__10560),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13483),
            .ce(N__10383),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_5_LC_16_13_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_5_LC_16_13_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_5_LC_16_13_5 .LUT_INIT=16'b1010101000110000;
    LogicCell40 \DUT.uart_inst0.tx_data_5_LC_16_13_5  (
            .in0(N__10554),
            .in1(N__11054),
            .in2(N__11112),
            .in3(N__10544),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13483),
            .ce(N__10383),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_16_14_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_16_14_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_16_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_16_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12876),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13478),
            .ce(N__11157),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_16_14_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_16_14_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_16_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_16_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13231),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13478),
            .ce(N__11157),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_16_14_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_16_14_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_16_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_16_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12918),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13478),
            .ce(N__11157),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_16_14_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_16_14_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_16_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_16_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14012),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13478),
            .ce(N__11157),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_16_14_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_16_14_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_16_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_16_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12522),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13478),
            .ce(N__11157),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_16_15_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_16_15_0 .LUT_INIT=16'b0000010111110011;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_16_15_0  (
            .in0(N__10659),
            .in1(N__10608),
            .in2(N__12759),
            .in3(N__12849),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_16_15_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_16_15_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_16_15_1  (
            .in0(N__11202),
            .in1(N__10590),
            .in2(N__10626),
            .in3(N__12757),
            .lcout(\DUT.rFifoDatarx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_16_15_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_16_15_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_16_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_16_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11242),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13471),
            .ce(N__13181),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_16_15_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_16_15_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_16_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_16_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14004),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13471),
            .ce(N__13181),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_16_15_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_16_15_6 .LUT_INIT=16'b0000010111110011;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_16_15_6  (
            .in0(N__10578),
            .in1(N__12543),
            .in2(N__12758),
            .in3(N__12848),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_16_15_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_16_15_7 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_16_15_7  (
            .in0(N__11190),
            .in1(N__10584),
            .in2(N__10602),
            .in3(N__12756),
            .lcout(\DUT.rFifoDatarx_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_16_16_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_16_16_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_16_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_16_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12613),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13467),
            .ce(N__11156),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_16_16_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_16_16_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_16_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_16_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11243),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13467),
            .ce(N__11156),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_16_16_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_16_16_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_16_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_16_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12583),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13467),
            .ce(N__11156),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_16_17_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_16_17_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_16_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_16_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12582),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13461),
            .ce(N__13954),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_16_17_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_16_17_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_16_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_16_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11247),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13461),
            .ce(N__13954),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIDL6N_7_LC_17_9_0 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIDL6N_7_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIDL6N_7_LC_17_9_0 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIDL6N_7_LC_17_9_0  (
            .in0(N__10650),
            .in1(N__13854),
            .in2(N__12480),
            .in3(N__10673),
            .lcout(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_7_LC_17_9_1 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_7_LC_17_9_1 .SEQ_MODE=4'b1010;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_7_LC_17_9_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_7_LC_17_9_1  (
            .in0(N__10674),
            .in1(_gnd_net_),
            .in2(N__12477),
            .in3(_gnd_net_),
            .lcout(\fifo_inst.tx_fifo_inst.rRamRdAddr_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13497),
            .ce(N__11287),
            .sr(N__13292));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_4_LC_17_9_2 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_4_LC_17_9_2 .SEQ_MODE=4'b1010;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_4_LC_17_9_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_4_LC_17_9_2  (
            .in0(N__10701),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12462),
            .lcout(\fifo_inst.tx_fifo_inst.rRamRdAddr_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13497),
            .ce(N__11287),
            .sr(N__13292));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIKR111_4_LC_17_9_3 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIKR111_4_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIKR111_4_LC_17_9_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIKR111_4_LC_17_9_3  (
            .in0(N__11580),
            .in1(N__10644),
            .in2(N__12478),
            .in3(N__10700),
            .lcout(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_6_LC_17_9_4 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_6_LC_17_9_4 .SEQ_MODE=4'b1010;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_6_LC_17_9_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_6_LC_17_9_4  (
            .in0(N__10686),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12463),
            .lcout(\fifo_inst.tx_fifo_inst.rRamRdAddr_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13497),
            .ce(N__11287),
            .sr(N__13292));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIO1411_6_LC_17_9_5 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIO1411_6_LC_17_9_5 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIO1411_6_LC_17_9_5 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIO1411_6_LC_17_9_5  (
            .in0(N__11579),
            .in1(N__10638),
            .in2(N__12479),
            .in3(N__10685),
            .lcout(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_0_LC_17_9_7 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_0_LC_17_9_7 .SEQ_MODE=4'b1010;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_0_LC_17_9_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_0_LC_17_9_7  (
            .in0(N__12461),
            .in1(N__11494),
            .in2(_gnd_net_),
            .in3(N__11543),
            .lcout(\fifo_inst.tx_fifo_inst.rRamRdAddr_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13497),
            .ce(N__11287),
            .sr(N__13292));
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1_c_LC_17_10_0 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1_c_LC_17_10_0 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1_c_LC_17_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1_c_LC_17_10_0  (
            .in0(_gnd_net_),
            .in1(N__10632),
            .in2(N__11495),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1_c_RNI5G02_LC_17_10_1 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1_c_RNI5G02_LC_17_10_1 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1_c_RNI5G02_LC_17_10_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1_c_RNI5G02_LC_17_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10766),
            .in3(N__10734),
            .lcout(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1_c_RNI5GZ0Z02 ),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_1 ),
            .carryout(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI6I12_LC_17_10_2 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI6I12_LC_17_10_2 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI6I12_LC_17_10_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI6I12_LC_17_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11516),
            .in3(N__10731),
            .lcout(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI6IZ0Z12 ),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2 ),
            .carryout(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_3_c_RNI7K22_LC_17_10_3 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_3_c_RNI7K22_LC_17_10_3 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_3_c_RNI7K22_LC_17_10_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_3_c_RNI7K22_LC_17_10_3  (
            .in0(_gnd_net_),
            .in1(N__10720),
            .in2(_gnd_net_),
            .in3(N__10692),
            .lcout(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_3_c_RNI7KZ0Z22 ),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_3 ),
            .carryout(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_4_c_RNI44E4_LC_17_10_4 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_4_c_RNI44E4_LC_17_10_4 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_4_c_RNI44E4_LC_17_10_4 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_4_c_RNI44E4_LC_17_10_4  (
            .in0(N__12162),
            .in1(_gnd_net_),
            .in2(N__11659),
            .in3(N__10689),
            .lcout(\fifo_inst.tx_fifo_inst.rRamRdAddr_rst_4 ),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_4 ),
            .carryout(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_5_c_RNI9O42_LC_17_10_5 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_5_c_RNI9O42_LC_17_10_5 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_5_c_RNI9O42_LC_17_10_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_5_c_RNI9O42_LC_17_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10852),
            .in3(N__10677),
            .lcout(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_5_c_RNI9OZ0Z42 ),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_5 ),
            .carryout(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_6_c_RNIAQ52_LC_17_10_6 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_6_c_RNIAQ52_LC_17_10_6 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_6_c_RNIAQ52_LC_17_10_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_6_c_RNIAQ52_LC_17_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10882),
            .in3(N__10665),
            .lcout(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_6_c_RNIAQZ0Z52 ),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_6 ),
            .carryout(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_7_c_RNI7AH4_LC_17_10_7 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_7_c_RNI7AH4_LC_17_10_7 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_7_c_RNI7AH4_LC_17_10_7 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_7_c_RNI7AH4_LC_17_10_7  (
            .in0(N__11443),
            .in1(N__12163),
            .in2(_gnd_net_),
            .in3(N__10662),
            .lcout(\fifo_inst.tx_fifo_inst.rRamRdAddr_rst_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ft2232h_inst.rTxRdEn_RNIS0VN_LC_17_11_0 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rTxRdEn_RNIS0VN_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ft2232h_inst.rTxRdEn_RNIS0VN_LC_17_11_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fifo_inst.ft2232h_inst.rTxRdEn_RNIS0VN_LC_17_11_0  (
            .in0(_gnd_net_),
            .in1(N__10896),
            .in2(_gnd_net_),
            .in3(N__13828),
            .lcout(\fifo_inst.rTxRdEn_RNIS0VN ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNISDA2_LC_17_11_2 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNISDA2_LC_17_11_2 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNISDA2_LC_17_11_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNISDA2_LC_17_11_2  (
            .in0(N__12171),
            .in1(N__11620),
            .in2(_gnd_net_),
            .in3(N__11744),
            .lcout(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ft2232h_inst.rFifoState_RNIG8PK_4_LC_17_11_3 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rFifoState_RNIG8PK_4_LC_17_11_3 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ft2232h_inst.rFifoState_RNIG8PK_4_LC_17_11_3 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \fifo_inst.ft2232h_inst.rFifoState_RNIG8PK_4_LC_17_11_3  (
            .in0(N__13827),
            .in1(N__12169),
            .in2(_gnd_net_),
            .in3(N__13911),
            .lcout(\fifo_inst.ft2232h_inst.rFifoState_RNIG8PKZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_3_1_LC_17_11_4 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_3_1_LC_17_11_4 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_3_1_LC_17_11_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIA4VU_3_1_LC_17_11_4  (
            .in0(N__10889),
            .in1(N__10853),
            .in2(N__11421),
            .in3(N__10827),
            .lcout(\fifo_inst.tx_fifo_inst.un15_rRamRdAddr ),
            .ltout(\fifo_inst.tx_fifo_inst.un15_rRamRdAddr_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNISDA2_0_LC_17_11_5 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNISDA2_0_LC_17_11_5 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNISDA2_0_LC_17_11_5 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_RNISDA2_0_LC_17_11_5  (
            .in0(_gnd_net_),
            .in1(N__12453),
            .in2(N__10821),
            .in3(N__11486),
            .lcout(),
            .ltout(\fifo_inst.tx_fifo_inst.rRamRdAddr_rst_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNISJ0L_0_LC_17_11_6 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNISJ0L_0_LC_17_11_6 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNISJ0L_0_LC_17_11_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_RNISJ0L_0_LC_17_11_6  (
            .in0(_gnd_net_),
            .in1(N__10818),
            .in2(N__10809),
            .in3(N__13826),
            .lcout(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ft2232h_inst.rTxRdEn_fast_LC_17_11_7 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rTxRdEn_fast_LC_17_11_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rTxRdEn_fast_LC_17_11_7 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \fifo_inst.ft2232h_inst.rTxRdEn_fast_LC_17_11_7  (
            .in0(N__13829),
            .in1(N__12170),
            .in2(_gnd_net_),
            .in3(N__13912),
            .lcout(\fifo_inst.rTxRdEn_fast ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13492),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_LC_17_12_0 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_LC_17_12_0 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_LC_17_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_LC_17_12_0  (
            .in0(_gnd_net_),
            .in1(N__11745),
            .in2(N__11775),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_17_12_0_),
            .carryout(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNII2L4_LC_17_12_1 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNII2L4_LC_17_12_1 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNII2L4_LC_17_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNII2L4_LC_17_12_1  (
            .in0(_gnd_net_),
            .in1(N__11604),
            .in2(_gnd_net_),
            .in3(N__10806),
            .lcout(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNII2LZ0Z4 ),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1 ),
            .carryout(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIJ4M4_LC_17_12_2 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIJ4M4_LC_17_12_2 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIJ4M4_LC_17_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIJ4M4_LC_17_12_2  (
            .in0(_gnd_net_),
            .in1(N__10803),
            .in2(_gnd_net_),
            .in3(N__10779),
            .lcout(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2_c_RNIJ4MZ0Z4 ),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_2 ),
            .carryout(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIK6N4_LC_17_12_3 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIK6N4_LC_17_12_3 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIK6N4_LC_17_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIK6N4_LC_17_12_3  (
            .in0(_gnd_net_),
            .in1(N__10920),
            .in2(_gnd_net_),
            .in3(N__10776),
            .lcout(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIK6NZ0Z4 ),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3 ),
            .carryout(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_4_c_RNIHM27_LC_17_12_4 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_4_c_RNIHM27_LC_17_12_4 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_4_c_RNIHM27_LC_17_12_4 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_4_c_RNIHM27_LC_17_12_4  (
            .in0(N__12179),
            .in1(_gnd_net_),
            .in2(N__11822),
            .in3(N__10989),
            .lcout(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_5 ),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_4 ),
            .carryout(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNIIO37_LC_17_12_5 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNIIO37_LC_17_12_5 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNIIO37_LC_17_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNIIO37_LC_17_12_5  (
            .in0(_gnd_net_),
            .in1(N__11928),
            .in2(_gnd_net_),
            .in3(N__10986),
            .lcout(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNIIOZ0Z37 ),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5 ),
            .carryout(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNIJQ47_LC_17_12_6 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNIJQ47_LC_17_12_6 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNIJQ47_LC_17_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNIJQ47_LC_17_12_6  (
            .in0(_gnd_net_),
            .in1(N__10983),
            .in2(_gnd_net_),
            .in3(N__10971),
            .lcout(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNIJQZ0Z47 ),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6 ),
            .carryout(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_7_c_RNIKS57_LC_17_12_7 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_7_c_RNIKS57_LC_17_12_7 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_7_c_RNIKS57_LC_17_12_7 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_7_c_RNIKS57_LC_17_12_7  (
            .in0(N__10948),
            .in1(N__12180),
            .in2(_gnd_net_),
            .in3(N__10968),
            .lcout(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_17_13_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_17_13_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_17_13_2 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_17_13_2  (
            .in0(N__13194),
            .in1(N__12724),
            .in2(N__11904),
            .in3(N__12845),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_17_13_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_17_13_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_17_13_3 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_17_13_3  (
            .in0(N__12725),
            .in1(N__11256),
            .in2(N__10935),
            .in3(N__10932),
            .lcout(\DUT.rFifoDatarx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIGK17_0_LC_17_13_5 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIGK17_0_LC_17_13_5 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIGK17_0_LC_17_13_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIGK17_0_LC_17_13_5  (
            .in0(_gnd_net_),
            .in1(N__12186),
            .in2(_gnd_net_),
            .in3(N__11852),
            .lcout(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_17_13_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_17_13_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_17_13_6 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_17_13_6  (
            .in0(N__10914),
            .in1(N__12726),
            .in2(N__11184),
            .in3(N__11691),
            .lcout(\DUT.rFifoDatarx_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_17_14_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_17_14_0 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_17_14_0  (
            .in0(N__12837),
            .in1(N__13971),
            .in2(N__12748),
            .in3(N__10902),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_17_14_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_17_14_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_17_14_1  (
            .in0(N__12723),
            .in1(N__10998),
            .in2(N__11121),
            .in3(N__11118),
            .lcout(\DUT.rFifoDatarx_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_17_14_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_17_14_3 .LUT_INIT=16'b0000010111110011;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_17_14_3  (
            .in0(N__11910),
            .in1(N__12855),
            .in2(N__12747),
            .in3(N__12836),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_17_14_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_17_14_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_17_14_4 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_17_14_4  (
            .in0(N__11103),
            .in1(N__11196),
            .in2(N__11097),
            .in3(N__12722),
            .lcout(\DUT.rFifoDatarx_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_17_14_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_17_14_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_17_14_5 .LUT_INIT=16'b0101000000111111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_17_14_5  (
            .in0(N__13518),
            .in1(N__11136),
            .in2(N__12746),
            .in3(N__12835),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoDataror_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_RNIJBAM_LC_17_14_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_RNIJBAM_LC_17_14_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_RNIJBAM_LC_17_14_6 .LUT_INIT=16'b1111000000110101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_0_RNIJBAM_LC_17_14_6  (
            .in0(N__11172),
            .in1(N__11082),
            .in2(N__11064),
            .in3(N__12721),
            .lcout(\DUT.rFifoDataror_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_17_14_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_17_14_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_17_14_7 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_17_14_7  (
            .in0(N__12720),
            .in1(N__11025),
            .in2(N__11007),
            .in3(N__12939),
            .lcout(\DUT.rFifoDatarxZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_17_15_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_17_15_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_17_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_17_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12928),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13479),
            .ce(N__13538),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_17_15_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_17_15_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_17_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_17_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14005),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13479),
            .ce(N__13538),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_17_15_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_17_15_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_17_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_17_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12635),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13479),
            .ce(N__13538),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_17_15_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_17_15_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_17_15_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_17_15_3  (
            .in0(N__13238),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13479),
            .ce(N__13538),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_17_15_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_17_15_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_17_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_17_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11241),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13479),
            .ce(N__13538),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_17_15_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_17_15_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_17_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_17_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12886),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13479),
            .ce(N__13538),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_17_15_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_17_15_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_17_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_17_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12588),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13479),
            .ce(N__13538),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_17_15_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_17_15_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_17_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_17_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12530),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13479),
            .ce(N__13538),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_1_LC_17_16_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_1_LC_17_16_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_1_LC_17_16_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_1_LC_17_16_3  (
            .in0(_gnd_net_),
            .in1(N__11171),
            .in2(_gnd_net_),
            .in3(N__13945),
            .lcout(\DUT.fifo_tx_inst.rFifoDataro_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13472),
            .ce(),
            .sr(N__13284));
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_1_LC_17_16_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_1_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_1_LC_17_16_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_1_LC_17_16_4  (
            .in0(N__11337),
            .in1(N__11363),
            .in2(_gnd_net_),
            .in3(N__13139),
            .lcout(\DUT.fifo_tx_inst.N_105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_LC_17_16_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_LC_17_16_5 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_LC_17_16_5  (
            .in0(N__13140),
            .in1(N__11364),
            .in2(_gnd_net_),
            .in3(N__11338),
            .lcout(\DUT.fifo_tx_inst.rFifoData_awe2 ),
            .ltout(\DUT.fifo_tx_inst.rFifoData_awe2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_LC_17_16_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_LC_17_16_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_LC_17_16_6 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_2_LC_17_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11139),
            .in3(N__11135),
            .lcout(\DUT.fifo_tx_inst.rFifoDataro_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13472),
            .ce(),
            .sr(N__13284));
    defparam \DUT.fifo_tx_inst.rWritePtr_1_LC_17_17_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_1_LC_17_17_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rWritePtr_1_LC_17_17_0 .LUT_INIT=16'b0000101100000100;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_1_LC_17_17_0  (
            .in0(N__13138),
            .in1(N__11336),
            .in2(N__11376),
            .in3(N__11362),
            .lcout(\DUT.fifo_tx_inst.rWritePtrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13468),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_2_1_LC_17_17_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_2_1_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_2_1_LC_17_17_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_RNIN79A_2_1_LC_17_17_1  (
            .in0(N__11360),
            .in1(N__13022),
            .in2(N__11339),
            .in3(N__13573),
            .lcout(\DUT.fifo_tx_inst.rFifoData_awe3 ),
            .ltout(\DUT.fifo_tx_inst.rFifoData_awe3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIJLJC_1_LC_17_17_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIJLJC_1_LC_17_17_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIJLJC_1_LC_17_17_2 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_RNIJLJC_1_LC_17_17_2  (
            .in0(N__12190),
            .in1(_gnd_net_),
            .in2(N__11379),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_tx_inst.un1_i11_i ),
            .ltout(\DUT.fifo_tx_inst.un1_i11_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_0_LC_17_17_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_0_LC_17_17_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rWritePtr_0_LC_17_17_3 .LUT_INIT=16'b0000101000000101;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_0_LC_17_17_3  (
            .in0(N__11335),
            .in1(_gnd_net_),
            .in2(N__11367),
            .in3(N__13137),
            .lcout(\DUT.fifo_tx_inst.rWritePtrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13468),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_0_1_LC_17_17_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_0_1_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_0_1_LC_17_17_7 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_RNIN79A_0_1_LC_17_17_7  (
            .in0(N__11361),
            .in1(_gnd_net_),
            .in2(N__11340),
            .in3(N__13136),
            .lcout(\DUT.fifo_tx_inst.rFifoData_awe1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIFO7N_8_LC_18_9_1 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIFO7N_8_LC_18_9_1 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIFO7N_8_LC_18_9_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIFO7N_8_LC_18_9_1  (
            .in0(N__11298),
            .in1(N__13843),
            .in2(_gnd_net_),
            .in3(N__11309),
            .lcout(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_5_LC_18_10_0 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_5_LC_18_10_0 .SEQ_MODE=4'b1010;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_5_LC_18_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_5_LC_18_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11684),
            .lcout(\fifo_inst.tx_fifo_inst.rRamRdAddr_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13498),
            .ce(N__11292),
            .sr(N__13293));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_8_LC_18_10_1 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_8_LC_18_10_1 .SEQ_MODE=4'b1010;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_8_LC_18_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_8_LC_18_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11310),
            .lcout(\fifo_inst.tx_fifo_inst.rRamRdAddr_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13498),
            .ce(N__11292),
            .sr(N__13293));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_3_LC_18_10_6 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_3_LC_18_10_6 .SEQ_MODE=4'b1010;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_3_LC_18_10_6 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_3_LC_18_10_6  (
            .in0(N__12460),
            .in1(_gnd_net_),
            .in2(N__11544),
            .in3(N__11597),
            .lcout(\fifo_inst.tx_fifo_inst.rRamRdAddr_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13498),
            .ce(N__11292),
            .sr(N__13293));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNI9F4N_5_LC_18_11_0 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNI9F4N_5_LC_18_11_0 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNI9F4N_5_LC_18_11_0 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_RNI9F4N_5_LC_18_11_0  (
            .in0(N__11685),
            .in1(_gnd_net_),
            .in2(N__13838),
            .in3(N__11673),
            .lcout(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNI111S_LC_18_11_1 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNI111S_LC_18_11_1 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNI111S_LC_18_11_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNI111S_LC_18_11_1  (
            .in0(N__11864),
            .in1(N__11781),
            .in2(N__11402),
            .in3(N__11637),
            .lcout(\fifo_inst.tx_fifo_inst.un18_rRamWrAddr ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIEGV6_0_LC_18_11_2 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIEGV6_0_LC_18_11_2 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIEGV6_0_LC_18_11_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIEGV6_0_LC_18_11_2  (
            .in0(N__12177),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11411),
            .lcout(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI20C4_LC_18_11_3 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI20C4_LC_18_11_3 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI20C4_LC_18_11_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI20C4_LC_18_11_3  (
            .in0(N__12436),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11598),
            .lcout(),
            .ltout(\fifo_inst.tx_fifo_inst.un17_rRamRdAddr_1_cry_2_c_RNI20CZ0Z4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIIO011_3_LC_18_11_4 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIIO011_3_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIIO011_3_LC_18_11_4 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_RNIIO011_3_LC_18_11_4  (
            .in0(N__11586),
            .in1(N__11578),
            .in2(N__11547),
            .in3(N__11536),
            .lcout(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_3 ),
            .ltout(\fifo_inst.tx_fifo_inst.rRamRdAddrZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNI_8_LC_18_11_5 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNI_8_LC_18_11_5 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNI_8_LC_18_11_5 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_RNI_8_LC_18_11_5  (
            .in0(N__11487),
            .in1(_gnd_net_),
            .in2(N__11448),
            .in3(N__11444),
            .lcout(\fifo_inst.tx_fifo_inst.un15_rRamRdAddr_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ft2232h_inst.rTxRdEn_LC_18_11_6 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rTxRdEn_LC_18_11_6 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rTxRdEn_LC_18_11_6 .LUT_INIT=16'b0010100000101000;
    LogicCell40 \fifo_inst.ft2232h_inst.rTxRdEn_LC_18_11_6  (
            .in0(N__12176),
            .in1(N__13913),
            .in2(N__13839),
            .in3(_gnd_net_),
            .lcout(\fifo_inst.wTxRdEn ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13495),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIEGV6_LC_18_11_7 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIEGV6_LC_18_11_7 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIEGV6_LC_18_11_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIEGV6_LC_18_11_7  (
            .in0(N__11412),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12178),
            .lcout(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNISDA2_LC_18_12_0 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNISDA2_LC_18_12_0 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNISDA2_LC_18_12_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNISDA2_LC_18_12_0  (
            .in0(_gnd_net_),
            .in1(N__12184),
            .in2(_gnd_net_),
            .in3(N__11939),
            .lcout(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNISDA2_LC_18_12_1 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNISDA2_LC_18_12_1 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNISDA2_LC_18_12_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_6_c_RNISDA2_LC_18_12_1  (
            .in0(N__12185),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11882),
            .lcout(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIGK17_LC_18_12_2 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIGK17_LC_18_12_2 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIGK17_LC_18_12_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_3_c_RNIGK17_LC_18_12_2  (
            .in0(N__11853),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12183),
            .lcout(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_4 ),
            .ltout(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIQIBG_LC_18_12_3 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIQIBG_LC_18_12_3 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIQIBG_LC_18_12_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIQIBG_LC_18_12_3  (
            .in0(N__11818),
            .in1(N__11795),
            .in2(N__11784),
            .in3(N__11702),
            .lcout(\fifo_inst.tx_fifo_inst.un18_rRamWrAddr_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNISDA2_2_LC_18_12_4 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNISDA2_2_LC_18_12_4 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNISDA2_2_LC_18_12_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNISDA2_2_LC_18_12_4  (
            .in0(N__11718),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12182),
            .lcout(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_1 ),
            .ltout(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNI_LC_18_12_5 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNI_LC_18_12_5 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNI_LC_18_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNI_LC_18_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11763),
            .in3(N__11749),
            .lcout(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIZ0 ),
            .ltout(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNIZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNISDA2_1_LC_18_12_6 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNISDA2_1_LC_18_12_6 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNISDA2_1_LC_18_12_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_1_c_RNISDA2_1_LC_18_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11712),
            .in3(N__12181),
            .lcout(\fifo_inst.tx_fifo_inst.rRamWrAddrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_18_13_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_18_13_0 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_18_13_0  (
            .in0(N__12834),
            .in1(N__11895),
            .in2(N__12745),
            .in3(N__12492),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rReadPtr_RNINFEP_0_LC_18_13_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rReadPtr_RNINFEP_0_LC_18_13_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rReadPtr_RNINFEP_0_LC_18_13_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \DUT.fifo_tx_inst.rReadPtr_RNINFEP_0_LC_18_13_1  (
            .in0(N__12846),
            .in1(N__13114),
            .in2(_gnd_net_),
            .in3(N__13082),
            .lcout(\DUT.fifo_tx_inst.N_101 ),
            .ltout(\DUT.fifo_tx_inst.N_101_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rReadPtr_RNILV421_1_LC_18_13_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rReadPtr_RNILV421_1_LC_18_13_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rReadPtr_RNILV421_1_LC_18_13_2 .LUT_INIT=16'b1010000011111111;
    LogicCell40 \DUT.fifo_tx_inst.rReadPtr_RNILV421_1_LC_18_13_2  (
            .in0(N__12713),
            .in1(_gnd_net_),
            .in2(N__12483),
            .in3(N__12435),
            .lcout(\DUT.fifo_tx_inst.un1_i11_2_i ),
            .ltout(\DUT.fifo_tx_inst.un1_i11_2_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rReadPtr_0_LC_18_13_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rReadPtr_0_LC_18_13_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rReadPtr_0_LC_18_13_3 .LUT_INIT=16'b0000011000001010;
    LogicCell40 \DUT.fifo_tx_inst.rReadPtr_0_LC_18_13_3  (
            .in0(N__12847),
            .in1(N__13115),
            .in2(N__12195),
            .in3(N__13083),
            .lcout(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13489),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNISDA2_0_LC_18_13_6 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNISDA2_0_LC_18_13_6 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNISDA2_0_LC_18_13_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_cry_5_c_RNISDA2_0_LC_18_13_6  (
            .in0(_gnd_net_),
            .in1(N__12189),
            .in2(_gnd_net_),
            .in3(N__11940),
            .lcout(\fifo_inst.tx_fifo_inst.un20_rRamWrAddr_1_axb_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rReadPtr_1_LC_18_13_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rReadPtr_1_LC_18_13_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rReadPtr_1_LC_18_13_7 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \DUT.fifo_tx_inst.rReadPtr_1_LC_18_13_7  (
            .in0(N__12730),
            .in1(N__11922),
            .in2(_gnd_net_),
            .in3(N__11916),
            .lcout(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13489),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_18_14_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_18_14_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_18_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_18_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12933),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13488),
            .ce(N__13961),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_18_14_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_18_14_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_18_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_18_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12891),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13488),
            .ce(N__13961),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_18_14_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_18_14_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_18_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_18_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13239),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13488),
            .ce(N__13961),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_18_14_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_18_14_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_18_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_18_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12531),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13488),
            .ce(N__13961),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_18_14_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_18_14_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_18_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_18_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12636),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13488),
            .ce(N__13961),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_18_15_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_18_15_0 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_18_15_0  (
            .in0(N__12838),
            .in1(N__12945),
            .in2(N__12749),
            .in3(N__12897),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_18_15_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_18_15_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_18_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_18_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12929),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13484),
            .ce(N__13185),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_18_15_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_18_15_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_18_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_18_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12887),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13484),
            .ce(N__13185),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_18_15_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_18_15_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_18_15_6 .LUT_INIT=16'b0010001101100111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_18_15_6  (
            .in0(N__12734),
            .in1(N__12839),
            .in2(N__12597),
            .in3(N__12786),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_18_15_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_18_15_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_18_15_7 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_18_15_7  (
            .in0(N__12780),
            .in1(N__12774),
            .in2(N__12762),
            .in3(N__12735),
            .lcout(\DUT.rFifoDatarx_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_18_16_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_18_16_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_18_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_18_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12631),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13480),
            .ce(N__13174),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_18_16_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_18_16_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_18_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_18_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12584),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13480),
            .ce(N__13174),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_18_16_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_18_16_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_18_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_18_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12529),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13480),
            .ce(N__13174),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_18_16_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_18_16_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_18_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_18_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13221),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13480),
            .ce(N__13174),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIN9O8_0_LC_18_17_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIN9O8_0_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIN9O8_0_LC_18_17_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNIN9O8_0_LC_18_17_0  (
            .in0(N__13567),
            .in1(N__13610),
            .in2(_gnd_net_),
            .in3(N__13656),
            .lcout(\DUT.N_93 ),
            .ltout(\DUT.N_93_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIEBIJ_0_LC_18_17_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIEBIJ_0_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIEBIJ_0_LC_18_17_1 .LUT_INIT=16'b1100111100110011;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNIEBIJ_0_LC_18_17_1  (
            .in0(_gnd_net_),
            .in1(N__13017),
            .in2(N__13146),
            .in3(N__13079),
            .lcout(\DUT.fifo_tx_inst.N_98 ),
            .ltout(\DUT.fifo_tx_inst.N_98_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_18_17_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_18_17_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_18_17_2 .LUT_INIT=16'b0000011100000111;
    LogicCell40 \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_18_17_2  (
            .in0(N__13569),
            .in1(N__13019),
            .in2(N__13143),
            .in3(N__13657),
            .lcout(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIMBD3_2_LC_18_17_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIMBD3_2_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIMBD3_2_LC_18_17_4 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNIMBD3_2_LC_18_17_4  (
            .in0(N__13568),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13018),
            .lcout(\DUT.fifo_tx_inst.N_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNO_0_2_LC_18_17_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNO_0_2_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNO_0_2_LC_18_17_6 .LUT_INIT=16'b1101001011110000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNO_0_2_LC_18_17_6  (
            .in0(N__13081),
            .in1(N__13021),
            .in2(N__13577),
            .in3(N__13110),
            .lcout(\DUT.fifo_tx_inst.un1_rFifoCount_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIBPFM_1_LC_18_17_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIBPFM_1_LC_18_17_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIBPFM_1_LC_18_17_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNIBPFM_1_LC_18_17_7  (
            .in0(N__13020),
            .in1(N__13109),
            .in2(N__13614),
            .in3(N__13080),
            .lcout(\DUT.fifo_tx_inst.rFifoCount_RNIBPFMZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_0_LC_18_18_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_0_LC_18_18_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoCount_0_LC_18_18_5 .LUT_INIT=16'b1111000010000111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_0_LC_18_18_5  (
            .in0(N__13026),
            .in1(N__13578),
            .in2(N__13667),
            .in3(N__12972),
            .lcout(\DUT.fifo_tx_inst.rFifoCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13469),
            .ce(),
            .sr(N__13283));
    defparam \fifo_inst.ft2232h_inst.rFifoState_4_LC_20_13_6 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rFifoState_4_LC_20_13_6 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rFifoState_4_LC_20_13_6 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \fifo_inst.ft2232h_inst.rFifoState_4_LC_20_13_6  (
            .in0(N__12966),
            .in1(N__13898),
            .in2(_gnd_net_),
            .in3(N__13863),
            .lcout(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13496),
            .ce(),
            .sr(N__13291));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_20_14_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_20_14_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_20_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_20_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14016),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13493),
            .ce(N__13962),
            .sr(_gnd_net_));
    defparam \fifo_inst.ft2232h_inst.rTxBusReady_LC_20_15_7 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rTxBusReady_LC_20_15_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rTxBusReady_LC_20_15_7 .LUT_INIT=16'b1011111110101010;
    LogicCell40 \fifo_inst.ft2232h_inst.rTxBusReady_LC_20_15_7  (
            .in0(N__13929),
            .in1(N__13907),
            .in2(N__13870),
            .in3(N__13686),
            .lcout(rTxBusReady),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13490),
            .ce(),
            .sr(N__13288));
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_20_17_0 .C_ON=1'b1;
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_20_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_20_17_0  (
            .in0(_gnd_net_),
            .in1(N__13668),
            .in2(N__13638),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_20_17_0_),
            .carryout(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_1_LC_20_17_1 .C_ON=1'b1;
    defparam \DUT.fifo_tx_inst.rFifoCount_1_LC_20_17_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoCount_1_LC_20_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_1_LC_20_17_1  (
            .in0(_gnd_net_),
            .in1(N__13609),
            .in2(N__13626),
            .in3(N__13593),
            .lcout(\DUT.fifo_tx_inst.rFifoCountZ0Z_1 ),
            .ltout(),
            .carryin(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0 ),
            .carryout(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1 ),
            .clk(N__13485),
            .ce(),
            .sr(N__13287));
    defparam \DUT.fifo_tx_inst.rFifoCount_2_LC_20_17_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_2_LC_20_17_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoCount_2_LC_20_17_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_2_LC_20_17_2  (
            .in0(_gnd_net_),
            .in1(N__13590),
            .in2(_gnd_net_),
            .in3(N__13581),
            .lcout(\DUT.fifo_tx_inst.rFifoCountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13485),
            .ce(),
            .sr(N__13287));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_3_LC_21_15_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_3_LC_21_15_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_3_LC_21_15_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_3_LC_21_15_5  (
            .in0(_gnd_net_),
            .in1(N__13539),
            .in2(_gnd_net_),
            .in3(N__13514),
            .lcout(\DUT.fifo_tx_inst.rFifoDataro_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13494),
            .ce(),
            .sr(N__13290));
endmodule // top
