// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Mar 29 2020 23:01:15

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    ioFifoData,
    P1A9,
    P1A1,
    P1A8,
    oRx_n,
    P1A7,
    P1A3,
    iTxE_n,
    iRxF_n,
    iClk,
    P1A2,
    BTN_N,
    BTN1,
    oTx_n,
    P1A4);

    output [7:0] ioFifoData;
    output P1A9;
    input P1A1;
    output P1A8;
    output oRx_n;
    output P1A7;
    output P1A3;
    input iTxE_n;
    input iRxF_n;
    input iClk;
    output P1A2;
    input BTN_N;
    input BTN1;
    output oTx_n;
    output P1A4;

    wire N__13526;
    wire N__13512;
    wire N__13511;
    wire N__13510;
    wire N__13503;
    wire N__13502;
    wire N__13501;
    wire N__13494;
    wire N__13493;
    wire N__13492;
    wire N__13485;
    wire N__13484;
    wire N__13483;
    wire N__13476;
    wire N__13475;
    wire N__13474;
    wire N__13467;
    wire N__13466;
    wire N__13465;
    wire N__13458;
    wire N__13457;
    wire N__13456;
    wire N__13449;
    wire N__13448;
    wire N__13447;
    wire N__13440;
    wire N__13439;
    wire N__13438;
    wire N__13431;
    wire N__13430;
    wire N__13429;
    wire N__13422;
    wire N__13421;
    wire N__13420;
    wire N__13413;
    wire N__13412;
    wire N__13411;
    wire N__13404;
    wire N__13403;
    wire N__13402;
    wire N__13395;
    wire N__13394;
    wire N__13393;
    wire N__13386;
    wire N__13385;
    wire N__13384;
    wire N__13377;
    wire N__13376;
    wire N__13375;
    wire N__13368;
    wire N__13367;
    wire N__13366;
    wire N__13359;
    wire N__13358;
    wire N__13357;
    wire N__13350;
    wire N__13349;
    wire N__13348;
    wire N__13341;
    wire N__13340;
    wire N__13339;
    wire N__13322;
    wire N__13321;
    wire N__13320;
    wire N__13319;
    wire N__13316;
    wire N__13313;
    wire N__13310;
    wire N__13307;
    wire N__13302;
    wire N__13299;
    wire N__13296;
    wire N__13293;
    wire N__13288;
    wire N__13283;
    wire N__13280;
    wire N__13277;
    wire N__13276;
    wire N__13275;
    wire N__13274;
    wire N__13271;
    wire N__13268;
    wire N__13265;
    wire N__13262;
    wire N__13259;
    wire N__13254;
    wire N__13251;
    wire N__13248;
    wire N__13245;
    wire N__13242;
    wire N__13235;
    wire N__13232;
    wire N__13229;
    wire N__13228;
    wire N__13225;
    wire N__13222;
    wire N__13217;
    wire N__13216;
    wire N__13213;
    wire N__13210;
    wire N__13209;
    wire N__13204;
    wire N__13201;
    wire N__13196;
    wire N__13193;
    wire N__13190;
    wire N__13189;
    wire N__13188;
    wire N__13187;
    wire N__13184;
    wire N__13181;
    wire N__13178;
    wire N__13175;
    wire N__13172;
    wire N__13169;
    wire N__13164;
    wire N__13161;
    wire N__13158;
    wire N__13153;
    wire N__13148;
    wire N__13147;
    wire N__13144;
    wire N__13141;
    wire N__13140;
    wire N__13137;
    wire N__13134;
    wire N__13131;
    wire N__13130;
    wire N__13123;
    wire N__13120;
    wire N__13115;
    wire N__13112;
    wire N__13109;
    wire N__13106;
    wire N__13105;
    wire N__13102;
    wire N__13099;
    wire N__13098;
    wire N__13095;
    wire N__13092;
    wire N__13089;
    wire N__13088;
    wire N__13081;
    wire N__13078;
    wire N__13075;
    wire N__13072;
    wire N__13067;
    wire N__13064;
    wire N__13061;
    wire N__13058;
    wire N__13055;
    wire N__13054;
    wire N__13053;
    wire N__13052;
    wire N__13051;
    wire N__13050;
    wire N__13049;
    wire N__13048;
    wire N__13047;
    wire N__13046;
    wire N__13045;
    wire N__13044;
    wire N__13043;
    wire N__13042;
    wire N__13041;
    wire N__13040;
    wire N__13039;
    wire N__13038;
    wire N__13037;
    wire N__13036;
    wire N__13035;
    wire N__13034;
    wire N__13033;
    wire N__13032;
    wire N__13031;
    wire N__13030;
    wire N__13029;
    wire N__13028;
    wire N__13027;
    wire N__13026;
    wire N__13025;
    wire N__13024;
    wire N__13023;
    wire N__13022;
    wire N__13021;
    wire N__13020;
    wire N__13019;
    wire N__13018;
    wire N__13017;
    wire N__13016;
    wire N__13015;
    wire N__13014;
    wire N__13013;
    wire N__13012;
    wire N__13011;
    wire N__13010;
    wire N__13009;
    wire N__13008;
    wire N__13007;
    wire N__13006;
    wire N__13005;
    wire N__13004;
    wire N__13003;
    wire N__13002;
    wire N__13001;
    wire N__13000;
    wire N__12887;
    wire N__12884;
    wire N__12883;
    wire N__12880;
    wire N__12879;
    wire N__12876;
    wire N__12873;
    wire N__12870;
    wire N__12867;
    wire N__12862;
    wire N__12861;
    wire N__12856;
    wire N__12853;
    wire N__12848;
    wire N__12847;
    wire N__12846;
    wire N__12845;
    wire N__12844;
    wire N__12843;
    wire N__12842;
    wire N__12841;
    wire N__12840;
    wire N__12837;
    wire N__12834;
    wire N__12831;
    wire N__12828;
    wire N__12825;
    wire N__12822;
    wire N__12819;
    wire N__12818;
    wire N__12817;
    wire N__12816;
    wire N__12815;
    wire N__12814;
    wire N__12813;
    wire N__12812;
    wire N__12811;
    wire N__12808;
    wire N__12807;
    wire N__12804;
    wire N__12797;
    wire N__12788;
    wire N__12785;
    wire N__12782;
    wire N__12779;
    wire N__12776;
    wire N__12773;
    wire N__12770;
    wire N__12767;
    wire N__12764;
    wire N__12763;
    wire N__12762;
    wire N__12761;
    wire N__12760;
    wire N__12759;
    wire N__12758;
    wire N__12757;
    wire N__12756;
    wire N__12753;
    wire N__12752;
    wire N__12751;
    wire N__12748;
    wire N__12747;
    wire N__12744;
    wire N__12743;
    wire N__12742;
    wire N__12741;
    wire N__12736;
    wire N__12727;
    wire N__12718;
    wire N__12715;
    wire N__12712;
    wire N__12709;
    wire N__12706;
    wire N__12703;
    wire N__12702;
    wire N__12699;
    wire N__12696;
    wire N__12695;
    wire N__12692;
    wire N__12689;
    wire N__12686;
    wire N__12679;
    wire N__12676;
    wire N__12673;
    wire N__12670;
    wire N__12667;
    wire N__12660;
    wire N__12657;
    wire N__12648;
    wire N__12637;
    wire N__12636;
    wire N__12633;
    wire N__12628;
    wire N__12625;
    wire N__12618;
    wire N__12611;
    wire N__12608;
    wire N__12605;
    wire N__12602;
    wire N__12599;
    wire N__12596;
    wire N__12587;
    wire N__12584;
    wire N__12581;
    wire N__12576;
    wire N__12569;
    wire N__12566;
    wire N__12563;
    wire N__12560;
    wire N__12557;
    wire N__12554;
    wire N__12551;
    wire N__12548;
    wire N__12545;
    wire N__12542;
    wire N__12539;
    wire N__12536;
    wire N__12533;
    wire N__12530;
    wire N__12527;
    wire N__12524;
    wire N__12523;
    wire N__12520;
    wire N__12517;
    wire N__12514;
    wire N__12511;
    wire N__12506;
    wire N__12503;
    wire N__12500;
    wire N__12499;
    wire N__12498;
    wire N__12497;
    wire N__12494;
    wire N__12491;
    wire N__12488;
    wire N__12485;
    wire N__12480;
    wire N__12477;
    wire N__12474;
    wire N__12471;
    wire N__12466;
    wire N__12461;
    wire N__12458;
    wire N__12455;
    wire N__12452;
    wire N__12449;
    wire N__12446;
    wire N__12445;
    wire N__12442;
    wire N__12439;
    wire N__12438;
    wire N__12435;
    wire N__12432;
    wire N__12429;
    wire N__12422;
    wire N__12421;
    wire N__12418;
    wire N__12415;
    wire N__12410;
    wire N__12407;
    wire N__12404;
    wire N__12401;
    wire N__12398;
    wire N__12397;
    wire N__12394;
    wire N__12391;
    wire N__12390;
    wire N__12385;
    wire N__12382;
    wire N__12381;
    wire N__12376;
    wire N__12373;
    wire N__12368;
    wire N__12365;
    wire N__12362;
    wire N__12359;
    wire N__12356;
    wire N__12353;
    wire N__12350;
    wire N__12349;
    wire N__12346;
    wire N__12343;
    wire N__12338;
    wire N__12337;
    wire N__12334;
    wire N__12331;
    wire N__12326;
    wire N__12325;
    wire N__12322;
    wire N__12319;
    wire N__12316;
    wire N__12311;
    wire N__12310;
    wire N__12307;
    wire N__12304;
    wire N__12299;
    wire N__12298;
    wire N__12295;
    wire N__12292;
    wire N__12287;
    wire N__12286;
    wire N__12283;
    wire N__12280;
    wire N__12275;
    wire N__12274;
    wire N__12271;
    wire N__12268;
    wire N__12265;
    wire N__12260;
    wire N__12259;
    wire N__12256;
    wire N__12253;
    wire N__12248;
    wire N__12245;
    wire N__12242;
    wire N__12239;
    wire N__12236;
    wire N__12233;
    wire N__12230;
    wire N__12227;
    wire N__12226;
    wire N__12225;
    wire N__12224;
    wire N__12223;
    wire N__12222;
    wire N__12221;
    wire N__12218;
    wire N__12217;
    wire N__12216;
    wire N__12215;
    wire N__12208;
    wire N__12205;
    wire N__12200;
    wire N__12199;
    wire N__12196;
    wire N__12189;
    wire N__12182;
    wire N__12179;
    wire N__12170;
    wire N__12169;
    wire N__12168;
    wire N__12167;
    wire N__12166;
    wire N__12159;
    wire N__12158;
    wire N__12157;
    wire N__12156;
    wire N__12155;
    wire N__12154;
    wire N__12153;
    wire N__12148;
    wire N__12145;
    wire N__12142;
    wire N__12137;
    wire N__12130;
    wire N__12119;
    wire N__12116;
    wire N__12113;
    wire N__12110;
    wire N__12107;
    wire N__12104;
    wire N__12101;
    wire N__12098;
    wire N__12095;
    wire N__12092;
    wire N__12089;
    wire N__12086;
    wire N__12083;
    wire N__12080;
    wire N__12077;
    wire N__12074;
    wire N__12073;
    wire N__12072;
    wire N__12071;
    wire N__12070;
    wire N__12067;
    wire N__12066;
    wire N__12065;
    wire N__12064;
    wire N__12063;
    wire N__12062;
    wire N__12061;
    wire N__12060;
    wire N__12059;
    wire N__12056;
    wire N__12053;
    wire N__12050;
    wire N__12047;
    wire N__12044;
    wire N__12041;
    wire N__12036;
    wire N__12031;
    wire N__12028;
    wire N__12025;
    wire N__12022;
    wire N__12019;
    wire N__12016;
    wire N__12013;
    wire N__12010;
    wire N__12007;
    wire N__12004;
    wire N__12001;
    wire N__12000;
    wire N__11997;
    wire N__11994;
    wire N__11993;
    wire N__11990;
    wire N__11989;
    wire N__11986;
    wire N__11985;
    wire N__11982;
    wire N__11981;
    wire N__11980;
    wire N__11979;
    wire N__11978;
    wire N__11977;
    wire N__11976;
    wire N__11975;
    wire N__11930;
    wire N__11927;
    wire N__11924;
    wire N__11921;
    wire N__11920;
    wire N__11919;
    wire N__11918;
    wire N__11915;
    wire N__11912;
    wire N__11911;
    wire N__11910;
    wire N__11907;
    wire N__11904;
    wire N__11901;
    wire N__11894;
    wire N__11885;
    wire N__11884;
    wire N__11883;
    wire N__11882;
    wire N__11881;
    wire N__11880;
    wire N__11879;
    wire N__11878;
    wire N__11875;
    wire N__11872;
    wire N__11869;
    wire N__11868;
    wire N__11861;
    wire N__11856;
    wire N__11853;
    wire N__11850;
    wire N__11845;
    wire N__11834;
    wire N__11833;
    wire N__11830;
    wire N__11829;
    wire N__11826;
    wire N__11823;
    wire N__11822;
    wire N__11821;
    wire N__11818;
    wire N__11815;
    wire N__11812;
    wire N__11809;
    wire N__11804;
    wire N__11795;
    wire N__11792;
    wire N__11789;
    wire N__11786;
    wire N__11783;
    wire N__11780;
    wire N__11777;
    wire N__11774;
    wire N__11773;
    wire N__11772;
    wire N__11769;
    wire N__11768;
    wire N__11767;
    wire N__11766;
    wire N__11765;
    wire N__11764;
    wire N__11763;
    wire N__11760;
    wire N__11757;
    wire N__11754;
    wire N__11745;
    wire N__11740;
    wire N__11729;
    wire N__11728;
    wire N__11725;
    wire N__11724;
    wire N__11723;
    wire N__11720;
    wire N__11719;
    wire N__11718;
    wire N__11717;
    wire N__11714;
    wire N__11705;
    wire N__11700;
    wire N__11693;
    wire N__11690;
    wire N__11687;
    wire N__11686;
    wire N__11685;
    wire N__11684;
    wire N__11681;
    wire N__11680;
    wire N__11677;
    wire N__11672;
    wire N__11669;
    wire N__11666;
    wire N__11665;
    wire N__11664;
    wire N__11663;
    wire N__11662;
    wire N__11661;
    wire N__11660;
    wire N__11657;
    wire N__11652;
    wire N__11649;
    wire N__11638;
    wire N__11637;
    wire N__11636;
    wire N__11633;
    wire N__11628;
    wire N__11623;
    wire N__11618;
    wire N__11609;
    wire N__11608;
    wire N__11607;
    wire N__11606;
    wire N__11605;
    wire N__11604;
    wire N__11603;
    wire N__11602;
    wire N__11601;
    wire N__11600;
    wire N__11599;
    wire N__11598;
    wire N__11597;
    wire N__11596;
    wire N__11595;
    wire N__11594;
    wire N__11593;
    wire N__11590;
    wire N__11585;
    wire N__11582;
    wire N__11577;
    wire N__11576;
    wire N__11573;
    wire N__11570;
    wire N__11567;
    wire N__11566;
    wire N__11565;
    wire N__11564;
    wire N__11561;
    wire N__11558;
    wire N__11555;
    wire N__11552;
    wire N__11549;
    wire N__11548;
    wire N__11547;
    wire N__11546;
    wire N__11545;
    wire N__11542;
    wire N__11541;
    wire N__11538;
    wire N__11537;
    wire N__11536;
    wire N__11533;
    wire N__11530;
    wire N__11527;
    wire N__11524;
    wire N__11521;
    wire N__11508;
    wire N__11505;
    wire N__11500;
    wire N__11483;
    wire N__11480;
    wire N__11477;
    wire N__11472;
    wire N__11469;
    wire N__11462;
    wire N__11457;
    wire N__11438;
    wire N__11437;
    wire N__11434;
    wire N__11433;
    wire N__11432;
    wire N__11431;
    wire N__11428;
    wire N__11425;
    wire N__11420;
    wire N__11417;
    wire N__11416;
    wire N__11415;
    wire N__11414;
    wire N__11413;
    wire N__11412;
    wire N__11411;
    wire N__11410;
    wire N__11409;
    wire N__11408;
    wire N__11407;
    wire N__11406;
    wire N__11403;
    wire N__11398;
    wire N__11395;
    wire N__11388;
    wire N__11377;
    wire N__11374;
    wire N__11371;
    wire N__11368;
    wire N__11361;
    wire N__11358;
    wire N__11355;
    wire N__11342;
    wire N__11339;
    wire N__11336;
    wire N__11333;
    wire N__11330;
    wire N__11329;
    wire N__11326;
    wire N__11323;
    wire N__11318;
    wire N__11317;
    wire N__11314;
    wire N__11311;
    wire N__11306;
    wire N__11305;
    wire N__11302;
    wire N__11299;
    wire N__11296;
    wire N__11293;
    wire N__11288;
    wire N__11287;
    wire N__11284;
    wire N__11281;
    wire N__11276;
    wire N__11273;
    wire N__11272;
    wire N__11269;
    wire N__11268;
    wire N__11265;
    wire N__11262;
    wire N__11259;
    wire N__11252;
    wire N__11251;
    wire N__11248;
    wire N__11245;
    wire N__11240;
    wire N__11239;
    wire N__11238;
    wire N__11235;
    wire N__11230;
    wire N__11225;
    wire N__11222;
    wire N__11221;
    wire N__11218;
    wire N__11215;
    wire N__11210;
    wire N__11207;
    wire N__11204;
    wire N__11201;
    wire N__11198;
    wire N__11195;
    wire N__11192;
    wire N__11189;
    wire N__11186;
    wire N__11183;
    wire N__11180;
    wire N__11177;
    wire N__11174;
    wire N__11171;
    wire N__11168;
    wire N__11165;
    wire N__11162;
    wire N__11159;
    wire N__11156;
    wire N__11153;
    wire N__11150;
    wire N__11149;
    wire N__11146;
    wire N__11143;
    wire N__11138;
    wire N__11135;
    wire N__11132;
    wire N__11129;
    wire N__11126;
    wire N__11123;
    wire N__11122;
    wire N__11121;
    wire N__11120;
    wire N__11117;
    wire N__11112;
    wire N__11109;
    wire N__11108;
    wire N__11105;
    wire N__11100;
    wire N__11097;
    wire N__11094;
    wire N__11089;
    wire N__11086;
    wire N__11083;
    wire N__11080;
    wire N__11077;
    wire N__11074;
    wire N__11071;
    wire N__11066;
    wire N__11065;
    wire N__11062;
    wire N__11061;
    wire N__11058;
    wire N__11055;
    wire N__11052;
    wire N__11049;
    wire N__11044;
    wire N__11041;
    wire N__11038;
    wire N__11035;
    wire N__11032;
    wire N__11029;
    wire N__11026;
    wire N__11023;
    wire N__11020;
    wire N__11015;
    wire N__11012;
    wire N__11011;
    wire N__11010;
    wire N__11009;
    wire N__11006;
    wire N__11005;
    wire N__11000;
    wire N__10997;
    wire N__10994;
    wire N__10991;
    wire N__10982;
    wire N__10979;
    wire N__10976;
    wire N__10973;
    wire N__10970;
    wire N__10967;
    wire N__10964;
    wire N__10961;
    wire N__10958;
    wire N__10955;
    wire N__10952;
    wire N__10949;
    wire N__10946;
    wire N__10943;
    wire N__10940;
    wire N__10937;
    wire N__10934;
    wire N__10931;
    wire N__10928;
    wire N__10925;
    wire N__10922;
    wire N__10919;
    wire N__10916;
    wire N__10915;
    wire N__10914;
    wire N__10911;
    wire N__10910;
    wire N__10909;
    wire N__10908;
    wire N__10907;
    wire N__10906;
    wire N__10905;
    wire N__10904;
    wire N__10903;
    wire N__10902;
    wire N__10901;
    wire N__10896;
    wire N__10893;
    wire N__10886;
    wire N__10879;
    wire N__10872;
    wire N__10869;
    wire N__10856;
    wire N__10855;
    wire N__10854;
    wire N__10853;
    wire N__10852;
    wire N__10851;
    wire N__10850;
    wire N__10849;
    wire N__10848;
    wire N__10847;
    wire N__10846;
    wire N__10843;
    wire N__10842;
    wire N__10841;
    wire N__10840;
    wire N__10839;
    wire N__10836;
    wire N__10833;
    wire N__10832;
    wire N__10831;
    wire N__10830;
    wire N__10827;
    wire N__10826;
    wire N__10825;
    wire N__10822;
    wire N__10819;
    wire N__10816;
    wire N__10803;
    wire N__10790;
    wire N__10779;
    wire N__10776;
    wire N__10763;
    wire N__10760;
    wire N__10757;
    wire N__10754;
    wire N__10751;
    wire N__10748;
    wire N__10745;
    wire N__10742;
    wire N__10739;
    wire N__10736;
    wire N__10735;
    wire N__10734;
    wire N__10731;
    wire N__10730;
    wire N__10729;
    wire N__10726;
    wire N__10723;
    wire N__10718;
    wire N__10715;
    wire N__10710;
    wire N__10703;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10691;
    wire N__10688;
    wire N__10685;
    wire N__10684;
    wire N__10683;
    wire N__10682;
    wire N__10679;
    wire N__10672;
    wire N__10667;
    wire N__10664;
    wire N__10663;
    wire N__10660;
    wire N__10659;
    wire N__10658;
    wire N__10657;
    wire N__10656;
    wire N__10655;
    wire N__10654;
    wire N__10653;
    wire N__10652;
    wire N__10649;
    wire N__10648;
    wire N__10647;
    wire N__10644;
    wire N__10633;
    wire N__10630;
    wire N__10627;
    wire N__10624;
    wire N__10621;
    wire N__10616;
    wire N__10611;
    wire N__10598;
    wire N__10597;
    wire N__10596;
    wire N__10595;
    wire N__10594;
    wire N__10589;
    wire N__10586;
    wire N__10581;
    wire N__10574;
    wire N__10571;
    wire N__10568;
    wire N__10567;
    wire N__10564;
    wire N__10561;
    wire N__10558;
    wire N__10557;
    wire N__10556;
    wire N__10555;
    wire N__10554;
    wire N__10553;
    wire N__10550;
    wire N__10547;
    wire N__10536;
    wire N__10529;
    wire N__10528;
    wire N__10527;
    wire N__10526;
    wire N__10525;
    wire N__10524;
    wire N__10523;
    wire N__10522;
    wire N__10521;
    wire N__10502;
    wire N__10499;
    wire N__10496;
    wire N__10493;
    wire N__10492;
    wire N__10491;
    wire N__10490;
    wire N__10487;
    wire N__10484;
    wire N__10481;
    wire N__10478;
    wire N__10473;
    wire N__10470;
    wire N__10469;
    wire N__10466;
    wire N__10461;
    wire N__10458;
    wire N__10451;
    wire N__10448;
    wire N__10445;
    wire N__10442;
    wire N__10441;
    wire N__10438;
    wire N__10437;
    wire N__10434;
    wire N__10431;
    wire N__10428;
    wire N__10425;
    wire N__10424;
    wire N__10421;
    wire N__10418;
    wire N__10415;
    wire N__10412;
    wire N__10403;
    wire N__10400;
    wire N__10397;
    wire N__10394;
    wire N__10391;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10379;
    wire N__10376;
    wire N__10373;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10352;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10340;
    wire N__10337;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10322;
    wire N__10319;
    wire N__10316;
    wire N__10313;
    wire N__10310;
    wire N__10307;
    wire N__10304;
    wire N__10301;
    wire N__10298;
    wire N__10295;
    wire N__10292;
    wire N__10289;
    wire N__10286;
    wire N__10283;
    wire N__10280;
    wire N__10277;
    wire N__10274;
    wire N__10271;
    wire N__10268;
    wire N__10265;
    wire N__10262;
    wire N__10259;
    wire N__10256;
    wire N__10253;
    wire N__10250;
    wire N__10247;
    wire N__10246;
    wire N__10243;
    wire N__10240;
    wire N__10235;
    wire N__10234;
    wire N__10233;
    wire N__10232;
    wire N__10229;
    wire N__10226;
    wire N__10223;
    wire N__10220;
    wire N__10211;
    wire N__10208;
    wire N__10205;
    wire N__10202;
    wire N__10199;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10187;
    wire N__10184;
    wire N__10181;
    wire N__10180;
    wire N__10175;
    wire N__10172;
    wire N__10171;
    wire N__10170;
    wire N__10169;
    wire N__10166;
    wire N__10165;
    wire N__10162;
    wire N__10161;
    wire N__10158;
    wire N__10155;
    wire N__10150;
    wire N__10147;
    wire N__10146;
    wire N__10145;
    wire N__10142;
    wire N__10141;
    wire N__10140;
    wire N__10137;
    wire N__10134;
    wire N__10129;
    wire N__10126;
    wire N__10123;
    wire N__10120;
    wire N__10117;
    wire N__10116;
    wire N__10115;
    wire N__10112;
    wire N__10111;
    wire N__10108;
    wire N__10105;
    wire N__10102;
    wire N__10095;
    wire N__10092;
    wire N__10085;
    wire N__10082;
    wire N__10075;
    wire N__10072;
    wire N__10067;
    wire N__10064;
    wire N__10061;
    wire N__10056;
    wire N__10049;
    wire N__10046;
    wire N__10045;
    wire N__10042;
    wire N__10041;
    wire N__10040;
    wire N__10039;
    wire N__10036;
    wire N__10035;
    wire N__10032;
    wire N__10029;
    wire N__10026;
    wire N__10023;
    wire N__10020;
    wire N__10019;
    wire N__10016;
    wire N__10013;
    wire N__10010;
    wire N__10007;
    wire N__10004;
    wire N__10001;
    wire N__9998;
    wire N__9995;
    wire N__9988;
    wire N__9977;
    wire N__9976;
    wire N__9973;
    wire N__9970;
    wire N__9969;
    wire N__9968;
    wire N__9965;
    wire N__9962;
    wire N__9959;
    wire N__9956;
    wire N__9953;
    wire N__9950;
    wire N__9947;
    wire N__9938;
    wire N__9937;
    wire N__9936;
    wire N__9933;
    wire N__9928;
    wire N__9925;
    wire N__9922;
    wire N__9919;
    wire N__9916;
    wire N__9911;
    wire N__9908;
    wire N__9905;
    wire N__9902;
    wire N__9901;
    wire N__9898;
    wire N__9897;
    wire N__9896;
    wire N__9893;
    wire N__9890;
    wire N__9883;
    wire N__9880;
    wire N__9875;
    wire N__9874;
    wire N__9873;
    wire N__9872;
    wire N__9865;
    wire N__9862;
    wire N__9857;
    wire N__9856;
    wire N__9853;
    wire N__9852;
    wire N__9845;
    wire N__9844;
    wire N__9843;
    wire N__9840;
    wire N__9835;
    wire N__9830;
    wire N__9829;
    wire N__9826;
    wire N__9825;
    wire N__9822;
    wire N__9819;
    wire N__9816;
    wire N__9809;
    wire N__9806;
    wire N__9803;
    wire N__9802;
    wire N__9801;
    wire N__9798;
    wire N__9795;
    wire N__9792;
    wire N__9785;
    wire N__9782;
    wire N__9781;
    wire N__9780;
    wire N__9773;
    wire N__9772;
    wire N__9771;
    wire N__9770;
    wire N__9769;
    wire N__9766;
    wire N__9757;
    wire N__9752;
    wire N__9749;
    wire N__9748;
    wire N__9747;
    wire N__9744;
    wire N__9739;
    wire N__9734;
    wire N__9733;
    wire N__9732;
    wire N__9731;
    wire N__9730;
    wire N__9723;
    wire N__9720;
    wire N__9717;
    wire N__9716;
    wire N__9713;
    wire N__9706;
    wire N__9701;
    wire N__9698;
    wire N__9697;
    wire N__9694;
    wire N__9691;
    wire N__9688;
    wire N__9683;
    wire N__9680;
    wire N__9677;
    wire N__9676;
    wire N__9675;
    wire N__9672;
    wire N__9669;
    wire N__9666;
    wire N__9661;
    wire N__9656;
    wire N__9653;
    wire N__9650;
    wire N__9647;
    wire N__9646;
    wire N__9645;
    wire N__9642;
    wire N__9639;
    wire N__9636;
    wire N__9633;
    wire N__9630;
    wire N__9623;
    wire N__9620;
    wire N__9617;
    wire N__9614;
    wire N__9613;
    wire N__9612;
    wire N__9611;
    wire N__9610;
    wire N__9609;
    wire N__9608;
    wire N__9607;
    wire N__9606;
    wire N__9605;
    wire N__9602;
    wire N__9601;
    wire N__9600;
    wire N__9599;
    wire N__9596;
    wire N__9595;
    wire N__9592;
    wire N__9591;
    wire N__9590;
    wire N__9581;
    wire N__9580;
    wire N__9567;
    wire N__9566;
    wire N__9565;
    wire N__9564;
    wire N__9551;
    wire N__9548;
    wire N__9545;
    wire N__9542;
    wire N__9541;
    wire N__9540;
    wire N__9539;
    wire N__9536;
    wire N__9533;
    wire N__9530;
    wire N__9527;
    wire N__9524;
    wire N__9519;
    wire N__9516;
    wire N__9511;
    wire N__9506;
    wire N__9491;
    wire N__9490;
    wire N__9487;
    wire N__9486;
    wire N__9483;
    wire N__9480;
    wire N__9477;
    wire N__9474;
    wire N__9471;
    wire N__9464;
    wire N__9461;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9448;
    wire N__9445;
    wire N__9442;
    wire N__9439;
    wire N__9436;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9424;
    wire N__9419;
    wire N__9416;
    wire N__9415;
    wire N__9414;
    wire N__9411;
    wire N__9408;
    wire N__9403;
    wire N__9398;
    wire N__9395;
    wire N__9392;
    wire N__9389;
    wire N__9386;
    wire N__9385;
    wire N__9384;
    wire N__9381;
    wire N__9378;
    wire N__9375;
    wire N__9368;
    wire N__9365;
    wire N__9362;
    wire N__9359;
    wire N__9358;
    wire N__9357;
    wire N__9354;
    wire N__9351;
    wire N__9348;
    wire N__9341;
    wire N__9338;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9328;
    wire N__9327;
    wire N__9324;
    wire N__9319;
    wire N__9314;
    wire N__9311;
    wire N__9308;
    wire N__9305;
    wire N__9304;
    wire N__9303;
    wire N__9300;
    wire N__9297;
    wire N__9294;
    wire N__9287;
    wire N__9284;
    wire N__9281;
    wire N__9278;
    wire N__9277;
    wire N__9276;
    wire N__9273;
    wire N__9268;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9254;
    wire N__9253;
    wire N__9252;
    wire N__9249;
    wire N__9246;
    wire N__9243;
    wire N__9236;
    wire N__9233;
    wire N__9230;
    wire N__9227;
    wire N__9224;
    wire N__9221;
    wire N__9220;
    wire N__9219;
    wire N__9216;
    wire N__9211;
    wire N__9206;
    wire N__9203;
    wire N__9200;
    wire N__9197;
    wire N__9194;
    wire N__9191;
    wire N__9188;
    wire N__9185;
    wire N__9182;
    wire N__9181;
    wire N__9180;
    wire N__9177;
    wire N__9172;
    wire N__9167;
    wire N__9164;
    wire N__9161;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9146;
    wire N__9143;
    wire N__9142;
    wire N__9141;
    wire N__9138;
    wire N__9133;
    wire N__9128;
    wire N__9125;
    wire N__9122;
    wire N__9119;
    wire N__9118;
    wire N__9115;
    wire N__9114;
    wire N__9111;
    wire N__9106;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9092;
    wire N__9091;
    wire N__9090;
    wire N__9087;
    wire N__9084;
    wire N__9081;
    wire N__9074;
    wire N__9071;
    wire N__9068;
    wire N__9065;
    wire N__9064;
    wire N__9063;
    wire N__9060;
    wire N__9057;
    wire N__9052;
    wire N__9047;
    wire N__9044;
    wire N__9041;
    wire N__9038;
    wire N__9035;
    wire N__9034;
    wire N__9029;
    wire N__9026;
    wire N__9025;
    wire N__9024;
    wire N__9021;
    wire N__9020;
    wire N__9019;
    wire N__9018;
    wire N__9017;
    wire N__9016;
    wire N__9015;
    wire N__9012;
    wire N__9011;
    wire N__9010;
    wire N__9009;
    wire N__9006;
    wire N__9005;
    wire N__9004;
    wire N__9003;
    wire N__9000;
    wire N__8995;
    wire N__8978;
    wire N__8977;
    wire N__8976;
    wire N__8969;
    wire N__8968;
    wire N__8965;
    wire N__8964;
    wire N__8961;
    wire N__8956;
    wire N__8953;
    wire N__8950;
    wire N__8947;
    wire N__8946;
    wire N__8943;
    wire N__8938;
    wire N__8935;
    wire N__8930;
    wire N__8925;
    wire N__8920;
    wire N__8909;
    wire N__8906;
    wire N__8903;
    wire N__8900;
    wire N__8897;
    wire N__8894;
    wire N__8891;
    wire N__8888;
    wire N__8885;
    wire N__8882;
    wire N__8879;
    wire N__8878;
    wire N__8877;
    wire N__8874;
    wire N__8871;
    wire N__8868;
    wire N__8865;
    wire N__8862;
    wire N__8859;
    wire N__8852;
    wire N__8851;
    wire N__8848;
    wire N__8845;
    wire N__8844;
    wire N__8841;
    wire N__8838;
    wire N__8835;
    wire N__8832;
    wire N__8829;
    wire N__8826;
    wire N__8819;
    wire N__8816;
    wire N__8815;
    wire N__8812;
    wire N__8809;
    wire N__8804;
    wire N__8801;
    wire N__8800;
    wire N__8797;
    wire N__8794;
    wire N__8791;
    wire N__8788;
    wire N__8785;
    wire N__8782;
    wire N__8779;
    wire N__8776;
    wire N__8775;
    wire N__8770;
    wire N__8767;
    wire N__8762;
    wire N__8761;
    wire N__8756;
    wire N__8753;
    wire N__8752;
    wire N__8751;
    wire N__8750;
    wire N__8747;
    wire N__8744;
    wire N__8743;
    wire N__8740;
    wire N__8737;
    wire N__8732;
    wire N__8729;
    wire N__8728;
    wire N__8723;
    wire N__8722;
    wire N__8717;
    wire N__8714;
    wire N__8711;
    wire N__8708;
    wire N__8705;
    wire N__8702;
    wire N__8699;
    wire N__8698;
    wire N__8695;
    wire N__8692;
    wire N__8689;
    wire N__8686;
    wire N__8683;
    wire N__8680;
    wire N__8679;
    wire N__8674;
    wire N__8671;
    wire N__8668;
    wire N__8665;
    wire N__8662;
    wire N__8659;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8639;
    wire N__8638;
    wire N__8637;
    wire N__8636;
    wire N__8635;
    wire N__8632;
    wire N__8623;
    wire N__8618;
    wire N__8617;
    wire N__8614;
    wire N__8613;
    wire N__8612;
    wire N__8609;
    wire N__8608;
    wire N__8601;
    wire N__8596;
    wire N__8591;
    wire N__8590;
    wire N__8589;
    wire N__8586;
    wire N__8581;
    wire N__8576;
    wire N__8575;
    wire N__8574;
    wire N__8571;
    wire N__8570;
    wire N__8569;
    wire N__8568;
    wire N__8563;
    wire N__8560;
    wire N__8557;
    wire N__8552;
    wire N__8549;
    wire N__8546;
    wire N__8543;
    wire N__8534;
    wire N__8533;
    wire N__8532;
    wire N__8531;
    wire N__8530;
    wire N__8525;
    wire N__8522;
    wire N__8519;
    wire N__8516;
    wire N__8511;
    wire N__8504;
    wire N__8501;
    wire N__8498;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8485;
    wire N__8480;
    wire N__8477;
    wire N__8476;
    wire N__8475;
    wire N__8474;
    wire N__8471;
    wire N__8466;
    wire N__8463;
    wire N__8456;
    wire N__8453;
    wire N__8450;
    wire N__8449;
    wire N__8446;
    wire N__8443;
    wire N__8438;
    wire N__8437;
    wire N__8434;
    wire N__8431;
    wire N__8428;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8407;
    wire N__8404;
    wire N__8401;
    wire N__8396;
    wire N__8395;
    wire N__8392;
    wire N__8391;
    wire N__8390;
    wire N__8389;
    wire N__8388;
    wire N__8387;
    wire N__8382;
    wire N__8371;
    wire N__8366;
    wire N__8363;
    wire N__8362;
    wire N__8359;
    wire N__8358;
    wire N__8357;
    wire N__8354;
    wire N__8353;
    wire N__8352;
    wire N__8349;
    wire N__8348;
    wire N__8343;
    wire N__8340;
    wire N__8337;
    wire N__8336;
    wire N__8333;
    wire N__8332;
    wire N__8329;
    wire N__8328;
    wire N__8325;
    wire N__8320;
    wire N__8317;
    wire N__8314;
    wire N__8311;
    wire N__8308;
    wire N__8305;
    wire N__8300;
    wire N__8293;
    wire N__8290;
    wire N__8287;
    wire N__8284;
    wire N__8281;
    wire N__8278;
    wire N__8273;
    wire N__8268;
    wire N__8265;
    wire N__8262;
    wire N__8259;
    wire N__8256;
    wire N__8253;
    wire N__8246;
    wire N__8245;
    wire N__8240;
    wire N__8237;
    wire N__8234;
    wire N__8231;
    wire N__8228;
    wire N__8227;
    wire N__8224;
    wire N__8223;
    wire N__8222;
    wire N__8221;
    wire N__8218;
    wire N__8215;
    wire N__8210;
    wire N__8207;
    wire N__8198;
    wire N__8197;
    wire N__8196;
    wire N__8195;
    wire N__8194;
    wire N__8193;
    wire N__8192;
    wire N__8183;
    wire N__8182;
    wire N__8177;
    wire N__8176;
    wire N__8173;
    wire N__8170;
    wire N__8167;
    wire N__8164;
    wire N__8163;
    wire N__8162;
    wire N__8161;
    wire N__8158;
    wire N__8155;
    wire N__8150;
    wire N__8147;
    wire N__8144;
    wire N__8139;
    wire N__8126;
    wire N__8123;
    wire N__8120;
    wire N__8117;
    wire N__8114;
    wire N__8111;
    wire N__8108;
    wire N__8105;
    wire N__8102;
    wire N__8099;
    wire N__8096;
    wire N__8093;
    wire N__8090;
    wire N__8087;
    wire N__8084;
    wire N__8081;
    wire N__8078;
    wire N__8075;
    wire N__8072;
    wire N__8069;
    wire N__8066;
    wire N__8063;
    wire N__8060;
    wire N__8057;
    wire N__8054;
    wire N__8051;
    wire N__8048;
    wire N__8045;
    wire N__8042;
    wire N__8039;
    wire N__8036;
    wire N__8033;
    wire N__8030;
    wire N__8027;
    wire N__8024;
    wire N__8021;
    wire N__8018;
    wire N__8015;
    wire N__8012;
    wire N__8009;
    wire N__8006;
    wire N__8003;
    wire N__8002;
    wire N__7999;
    wire N__7996;
    wire N__7993;
    wire N__7990;
    wire N__7987;
    wire N__7982;
    wire N__7979;
    wire N__7976;
    wire N__7973;
    wire N__7970;
    wire N__7967;
    wire N__7964;
    wire N__7961;
    wire N__7958;
    wire N__7955;
    wire N__7952;
    wire N__7949;
    wire N__7946;
    wire N__7943;
    wire N__7940;
    wire N__7937;
    wire N__7936;
    wire N__7935;
    wire N__7930;
    wire N__7927;
    wire N__7926;
    wire N__7925;
    wire N__7924;
    wire N__7923;
    wire N__7922;
    wire N__7921;
    wire N__7920;
    wire N__7919;
    wire N__7918;
    wire N__7917;
    wire N__7914;
    wire N__7913;
    wire N__7910;
    wire N__7907;
    wire N__7904;
    wire N__7901;
    wire N__7900;
    wire N__7899;
    wire N__7896;
    wire N__7895;
    wire N__7894;
    wire N__7893;
    wire N__7888;
    wire N__7881;
    wire N__7878;
    wire N__7875;
    wire N__7872;
    wire N__7863;
    wire N__7858;
    wire N__7851;
    wire N__7848;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7814;
    wire N__7811;
    wire N__7810;
    wire N__7809;
    wire N__7806;
    wire N__7803;
    wire N__7802;
    wire N__7799;
    wire N__7794;
    wire N__7791;
    wire N__7788;
    wire N__7787;
    wire N__7784;
    wire N__7781;
    wire N__7778;
    wire N__7775;
    wire N__7766;
    wire N__7763;
    wire N__7760;
    wire N__7759;
    wire N__7758;
    wire N__7755;
    wire N__7754;
    wire N__7751;
    wire N__7748;
    wire N__7745;
    wire N__7742;
    wire N__7739;
    wire N__7732;
    wire N__7731;
    wire N__7728;
    wire N__7725;
    wire N__7722;
    wire N__7715;
    wire N__7712;
    wire N__7709;
    wire N__7708;
    wire N__7707;
    wire N__7704;
    wire N__7703;
    wire N__7700;
    wire N__7697;
    wire N__7694;
    wire N__7691;
    wire N__7688;
    wire N__7681;
    wire N__7680;
    wire N__7677;
    wire N__7674;
    wire N__7671;
    wire N__7664;
    wire N__7661;
    wire N__7658;
    wire N__7655;
    wire N__7654;
    wire N__7653;
    wire N__7652;
    wire N__7649;
    wire N__7646;
    wire N__7643;
    wire N__7640;
    wire N__7637;
    wire N__7632;
    wire N__7629;
    wire N__7628;
    wire N__7625;
    wire N__7620;
    wire N__7617;
    wire N__7610;
    wire N__7607;
    wire N__7604;
    wire N__7601;
    wire N__7598;
    wire N__7595;
    wire N__7592;
    wire N__7589;
    wire N__7586;
    wire N__7585;
    wire N__7582;
    wire N__7579;
    wire N__7576;
    wire N__7573;
    wire N__7570;
    wire N__7567;
    wire N__7562;
    wire N__7559;
    wire N__7556;
    wire N__7553;
    wire N__7550;
    wire N__7547;
    wire N__7546;
    wire N__7543;
    wire N__7540;
    wire N__7537;
    wire N__7534;
    wire N__7531;
    wire N__7528;
    wire N__7523;
    wire N__7522;
    wire N__7519;
    wire N__7516;
    wire N__7511;
    wire N__7508;
    wire N__7507;
    wire N__7504;
    wire N__7501;
    wire N__7496;
    wire N__7495;
    wire N__7490;
    wire N__7487;
    wire N__7484;
    wire N__7481;
    wire N__7480;
    wire N__7477;
    wire N__7474;
    wire N__7469;
    wire N__7468;
    wire N__7463;
    wire N__7460;
    wire N__7459;
    wire N__7456;
    wire N__7451;
    wire N__7448;
    wire N__7445;
    wire N__7442;
    wire N__7439;
    wire N__7436;
    wire N__7433;
    wire N__7430;
    wire N__7427;
    wire N__7426;
    wire N__7423;
    wire N__7422;
    wire N__7419;
    wire N__7418;
    wire N__7415;
    wire N__7412;
    wire N__7409;
    wire N__7406;
    wire N__7401;
    wire N__7396;
    wire N__7393;
    wire N__7390;
    wire N__7385;
    wire N__7382;
    wire N__7379;
    wire N__7376;
    wire N__7375;
    wire N__7374;
    wire N__7371;
    wire N__7370;
    wire N__7367;
    wire N__7364;
    wire N__7361;
    wire N__7358;
    wire N__7355;
    wire N__7352;
    wire N__7351;
    wire N__7348;
    wire N__7345;
    wire N__7340;
    wire N__7337;
    wire N__7328;
    wire N__7327;
    wire N__7326;
    wire N__7323;
    wire N__7320;
    wire N__7319;
    wire N__7316;
    wire N__7313;
    wire N__7310;
    wire N__7307;
    wire N__7304;
    wire N__7303;
    wire N__7298;
    wire N__7295;
    wire N__7292;
    wire N__7289;
    wire N__7280;
    wire N__7277;
    wire N__7274;
    wire N__7273;
    wire N__7272;
    wire N__7271;
    wire N__7268;
    wire N__7267;
    wire N__7266;
    wire N__7265;
    wire N__7264;
    wire N__7259;
    wire N__7256;
    wire N__7253;
    wire N__7244;
    wire N__7235;
    wire N__7234;
    wire N__7233;
    wire N__7230;
    wire N__7229;
    wire N__7228;
    wire N__7225;
    wire N__7222;
    wire N__7217;
    wire N__7214;
    wire N__7205;
    wire N__7202;
    wire N__7199;
    wire N__7196;
    wire N__7193;
    wire N__7190;
    wire N__7189;
    wire N__7184;
    wire N__7181;
    wire N__7180;
    wire N__7175;
    wire N__7172;
    wire N__7169;
    wire N__7168;
    wire N__7163;
    wire N__7160;
    wire N__7157;
    wire N__7154;
    wire N__7151;
    wire N__7148;
    wire N__7145;
    wire N__7142;
    wire N__7141;
    wire N__7140;
    wire N__7139;
    wire N__7138;
    wire N__7135;
    wire N__7132;
    wire N__7131;
    wire N__7130;
    wire N__7127;
    wire N__7122;
    wire N__7119;
    wire N__7112;
    wire N__7107;
    wire N__7106;
    wire N__7099;
    wire N__7096;
    wire N__7091;
    wire N__7088;
    wire N__7085;
    wire N__7082;
    wire N__7079;
    wire N__7076;
    wire N__7073;
    wire N__7072;
    wire N__7071;
    wire N__7070;
    wire N__7069;
    wire N__7068;
    wire N__7065;
    wire N__7062;
    wire N__7053;
    wire N__7046;
    wire N__7043;
    wire N__7040;
    wire N__7037;
    wire N__7034;
    wire N__7033;
    wire N__7032;
    wire N__7031;
    wire N__7030;
    wire N__7029;
    wire N__7026;
    wire N__7023;
    wire N__7020;
    wire N__7019;
    wire N__7018;
    wire N__7013;
    wire N__7010;
    wire N__7003;
    wire N__7002;
    wire N__6999;
    wire N__6998;
    wire N__6995;
    wire N__6994;
    wire N__6993;
    wire N__6986;
    wire N__6981;
    wire N__6974;
    wire N__6971;
    wire N__6966;
    wire N__6959;
    wire N__6956;
    wire N__6955;
    wire N__6954;
    wire N__6953;
    wire N__6948;
    wire N__6947;
    wire N__6942;
    wire N__6941;
    wire N__6940;
    wire N__6939;
    wire N__6938;
    wire N__6937;
    wire N__6936;
    wire N__6935;
    wire N__6932;
    wire N__6929;
    wire N__6926;
    wire N__6923;
    wire N__6918;
    wire N__6909;
    wire N__6906;
    wire N__6903;
    wire N__6890;
    wire N__6889;
    wire N__6886;
    wire N__6883;
    wire N__6880;
    wire N__6877;
    wire N__6872;
    wire N__6871;
    wire N__6870;
    wire N__6869;
    wire N__6864;
    wire N__6863;
    wire N__6862;
    wire N__6859;
    wire N__6858;
    wire N__6855;
    wire N__6854;
    wire N__6853;
    wire N__6852;
    wire N__6851;
    wire N__6848;
    wire N__6843;
    wire N__6840;
    wire N__6837;
    wire N__6834;
    wire N__6831;
    wire N__6828;
    wire N__6823;
    wire N__6818;
    wire N__6813;
    wire N__6800;
    wire N__6797;
    wire N__6796;
    wire N__6795;
    wire N__6794;
    wire N__6793;
    wire N__6792;
    wire N__6791;
    wire N__6790;
    wire N__6789;
    wire N__6788;
    wire N__6785;
    wire N__6782;
    wire N__6781;
    wire N__6780;
    wire N__6777;
    wire N__6768;
    wire N__6765;
    wire N__6760;
    wire N__6757;
    wire N__6754;
    wire N__6749;
    wire N__6734;
    wire N__6733;
    wire N__6732;
    wire N__6731;
    wire N__6730;
    wire N__6729;
    wire N__6726;
    wire N__6723;
    wire N__6720;
    wire N__6719;
    wire N__6714;
    wire N__6713;
    wire N__6712;
    wire N__6711;
    wire N__6708;
    wire N__6705;
    wire N__6700;
    wire N__6699;
    wire N__6698;
    wire N__6697;
    wire N__6696;
    wire N__6695;
    wire N__6692;
    wire N__6689;
    wire N__6688;
    wire N__6687;
    wire N__6686;
    wire N__6685;
    wire N__6680;
    wire N__6679;
    wire N__6678;
    wire N__6675;
    wire N__6672;
    wire N__6669;
    wire N__6666;
    wire N__6659;
    wire N__6654;
    wire N__6649;
    wire N__6644;
    wire N__6639;
    wire N__6636;
    wire N__6631;
    wire N__6628;
    wire N__6605;
    wire N__6602;
    wire N__6599;
    wire N__6596;
    wire N__6593;
    wire N__6590;
    wire N__6587;
    wire N__6584;
    wire N__6581;
    wire N__6578;
    wire N__6575;
    wire N__6572;
    wire N__6569;
    wire N__6566;
    wire N__6565;
    wire N__6564;
    wire N__6563;
    wire N__6562;
    wire N__6561;
    wire N__6560;
    wire N__6559;
    wire N__6558;
    wire N__6555;
    wire N__6554;
    wire N__6553;
    wire N__6550;
    wire N__6547;
    wire N__6542;
    wire N__6537;
    wire N__6532;
    wire N__6525;
    wire N__6522;
    wire N__6509;
    wire N__6506;
    wire N__6503;
    wire N__6500;
    wire N__6497;
    wire N__6494;
    wire N__6493;
    wire N__6492;
    wire N__6491;
    wire N__6488;
    wire N__6487;
    wire N__6484;
    wire N__6483;
    wire N__6482;
    wire N__6481;
    wire N__6480;
    wire N__6479;
    wire N__6478;
    wire N__6477;
    wire N__6474;
    wire N__6471;
    wire N__6468;
    wire N__6465;
    wire N__6462;
    wire N__6455;
    wire N__6446;
    wire N__6443;
    wire N__6428;
    wire N__6427;
    wire N__6426;
    wire N__6425;
    wire N__6424;
    wire N__6421;
    wire N__6420;
    wire N__6419;
    wire N__6416;
    wire N__6413;
    wire N__6412;
    wire N__6409;
    wire N__6406;
    wire N__6405;
    wire N__6404;
    wire N__6401;
    wire N__6400;
    wire N__6397;
    wire N__6396;
    wire N__6393;
    wire N__6390;
    wire N__6385;
    wire N__6382;
    wire N__6379;
    wire N__6374;
    wire N__6371;
    wire N__6368;
    wire N__6363;
    wire N__6344;
    wire N__6341;
    wire N__6338;
    wire N__6335;
    wire N__6334;
    wire N__6333;
    wire N__6332;
    wire N__6329;
    wire N__6326;
    wire N__6325;
    wire N__6322;
    wire N__6321;
    wire N__6320;
    wire N__6317;
    wire N__6316;
    wire N__6315;
    wire N__6314;
    wire N__6311;
    wire N__6308;
    wire N__6305;
    wire N__6302;
    wire N__6297;
    wire N__6294;
    wire N__6287;
    wire N__6284;
    wire N__6269;
    wire N__6266;
    wire N__6263;
    wire N__6260;
    wire N__6257;
    wire N__6254;
    wire N__6253;
    wire N__6252;
    wire N__6251;
    wire N__6250;
    wire N__6249;
    wire N__6248;
    wire N__6245;
    wire N__6244;
    wire N__6243;
    wire N__6242;
    wire N__6239;
    wire N__6238;
    wire N__6235;
    wire N__6234;
    wire N__6231;
    wire N__6228;
    wire N__6225;
    wire N__6220;
    wire N__6213;
    wire N__6208;
    wire N__6205;
    wire N__6202;
    wire N__6197;
    wire N__6182;
    wire N__6179;
    wire N__6176;
    wire N__6173;
    wire N__6170;
    wire N__6167;
    wire N__6164;
    wire N__6161;
    wire N__6158;
    wire N__6155;
    wire N__6152;
    wire N__6149;
    wire N__6146;
    wire N__6143;
    wire N__6142;
    wire N__6141;
    wire N__6140;
    wire N__6137;
    wire N__6136;
    wire N__6133;
    wire N__6132;
    wire N__6131;
    wire N__6130;
    wire N__6127;
    wire N__6126;
    wire N__6125;
    wire N__6124;
    wire N__6121;
    wire N__6118;
    wire N__6113;
    wire N__6108;
    wire N__6103;
    wire N__6100;
    wire N__6095;
    wire N__6092;
    wire N__6077;
    wire N__6074;
    wire N__6071;
    wire N__6068;
    wire N__6065;
    wire N__6062;
    wire N__6059;
    wire N__6058;
    wire N__6055;
    wire N__6052;
    wire N__6047;
    wire N__6046;
    wire N__6043;
    wire N__6042;
    wire N__6039;
    wire N__6034;
    wire N__6029;
    wire N__6026;
    wire N__6023;
    wire N__6020;
    wire N__6017;
    wire N__6014;
    wire N__6011;
    wire N__6008;
    wire N__6005;
    wire N__6002;
    wire N__5999;
    wire N__5996;
    wire N__5993;
    wire N__5990;
    wire N__5987;
    wire N__5984;
    wire N__5981;
    wire N__5978;
    wire N__5975;
    wire N__5972;
    wire N__5969;
    wire N__5966;
    wire N__5963;
    wire N__5960;
    wire N__5957;
    wire N__5954;
    wire N__5951;
    wire N__5948;
    wire N__5945;
    wire N__5942;
    wire N__5939;
    wire N__5936;
    wire N__5933;
    wire N__5930;
    wire N__5927;
    wire N__5924;
    wire N__5921;
    wire N__5918;
    wire N__5915;
    wire N__5912;
    wire N__5909;
    wire N__5906;
    wire N__5903;
    wire N__5900;
    wire N__5897;
    wire N__5894;
    wire N__5891;
    wire N__5888;
    wire N__5885;
    wire N__5882;
    wire N__5879;
    wire N__5876;
    wire N__5873;
    wire N__5870;
    wire N__5867;
    wire N__5864;
    wire N__5861;
    wire N__5858;
    wire N__5857;
    wire N__5856;
    wire N__5855;
    wire N__5850;
    wire N__5845;
    wire N__5840;
    wire N__5839;
    wire N__5836;
    wire N__5835;
    wire N__5834;
    wire N__5833;
    wire N__5826;
    wire N__5823;
    wire N__5822;
    wire N__5819;
    wire N__5816;
    wire N__5809;
    wire N__5804;
    wire N__5803;
    wire N__5802;
    wire N__5801;
    wire N__5800;
    wire N__5793;
    wire N__5788;
    wire N__5783;
    wire N__5780;
    wire N__5777;
    wire N__5774;
    wire N__5771;
    wire N__5768;
    wire N__5765;
    wire N__5762;
    wire N__5759;
    wire N__5756;
    wire N__5753;
    wire N__5750;
    wire N__5747;
    wire N__5744;
    wire N__5741;
    wire N__5738;
    wire N__5735;
    wire N__5732;
    wire N__5729;
    wire N__5726;
    wire N__5723;
    wire N__5720;
    wire N__5717;
    wire N__5714;
    wire N__5711;
    wire N__5708;
    wire N__5705;
    wire N__5702;
    wire N__5699;
    wire N__5696;
    wire N__5693;
    wire N__5690;
    wire N__5687;
    wire N__5684;
    wire N__5681;
    wire N__5678;
    wire N__5675;
    wire N__5672;
    wire N__5669;
    wire N__5666;
    wire N__5663;
    wire N__5660;
    wire N__5659;
    wire N__5658;
    wire N__5657;
    wire N__5654;
    wire N__5651;
    wire N__5646;
    wire N__5645;
    wire N__5644;
    wire N__5643;
    wire N__5642;
    wire N__5639;
    wire N__5634;
    wire N__5629;
    wire N__5626;
    wire N__5623;
    wire N__5612;
    wire N__5609;
    wire N__5606;
    wire N__5603;
    wire N__5600;
    wire N__5597;
    wire N__5594;
    wire N__5591;
    wire N__5588;
    wire N__5585;
    wire N__5582;
    wire N__5579;
    wire N__5576;
    wire N__5573;
    wire N__5570;
    wire N__5567;
    wire N__5564;
    wire N__5561;
    wire N__5558;
    wire N__5555;
    wire N__5552;
    wire N__5549;
    wire N__5546;
    wire N__5543;
    wire N__5540;
    wire N__5537;
    wire N__5534;
    wire N__5533;
    wire N__5532;
    wire N__5531;
    wire N__5530;
    wire N__5529;
    wire N__5528;
    wire N__5523;
    wire N__5522;
    wire N__5517;
    wire N__5512;
    wire N__5511;
    wire N__5508;
    wire N__5507;
    wire N__5506;
    wire N__5503;
    wire N__5500;
    wire N__5495;
    wire N__5492;
    wire N__5489;
    wire N__5486;
    wire N__5483;
    wire N__5468;
    wire N__5465;
    wire N__5462;
    wire N__5459;
    wire N__5456;
    wire N__5453;
    wire N__5450;
    wire N__5447;
    wire N__5444;
    wire N__5441;
    wire N__5438;
    wire N__5435;
    wire N__5432;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5411;
    wire N__5408;
    wire N__5407;
    wire N__5406;
    wire N__5405;
    wire N__5404;
    wire N__5403;
    wire N__5402;
    wire N__5401;
    wire N__5398;
    wire N__5395;
    wire N__5384;
    wire N__5381;
    wire N__5378;
    wire N__5375;
    wire N__5366;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5354;
    wire N__5351;
    wire N__5348;
    wire N__5347;
    wire N__5346;
    wire N__5339;
    wire N__5336;
    wire N__5333;
    wire N__5330;
    wire N__5327;
    wire N__5324;
    wire N__5321;
    wire N__5318;
    wire N__5315;
    wire N__5312;
    wire N__5311;
    wire N__5310;
    wire N__5307;
    wire N__5306;
    wire N__5303;
    wire N__5300;
    wire N__5299;
    wire N__5296;
    wire N__5295;
    wire N__5292;
    wire N__5287;
    wire N__5284;
    wire N__5281;
    wire N__5278;
    wire N__5273;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5255;
    wire N__5252;
    wire N__5249;
    wire N__5246;
    wire N__5243;
    wire N__5240;
    wire N__5237;
    wire N__5236;
    wire N__5235;
    wire N__5234;
    wire N__5231;
    wire N__5226;
    wire N__5223;
    wire N__5220;
    wire N__5217;
    wire N__5210;
    wire N__5209;
    wire N__5208;
    wire N__5205;
    wire N__5204;
    wire N__5203;
    wire N__5200;
    wire N__5197;
    wire N__5192;
    wire N__5189;
    wire N__5188;
    wire N__5187;
    wire N__5180;
    wire N__5177;
    wire N__5174;
    wire N__5171;
    wire N__5166;
    wire N__5159;
    wire N__5156;
    wire N__5153;
    wire N__5150;
    wire N__5147;
    wire N__5144;
    wire N__5141;
    wire N__5138;
    wire N__5135;
    wire N__5132;
    wire N__5129;
    wire N__5126;
    wire N__5123;
    wire N__5120;
    wire N__5117;
    wire N__5114;
    wire N__5111;
    wire N__5108;
    wire N__5105;
    wire N__5102;
    wire N__5099;
    wire N__5096;
    wire N__5093;
    wire N__5090;
    wire N__5087;
    wire N__5084;
    wire N__5081;
    wire N__5078;
    wire N__5075;
    wire N__5072;
    wire N__5069;
    wire BTN_N_c;
    wire VCCG0;
    wire GNDG0;
    wire \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO ;
    wire \DUT.uart_inst0.rx_bits_remaining_RNO_1Z0Z_1_cascade_ ;
    wire \DUT.uart_inst0.m5_1_1_cascade_ ;
    wire \DUT.uart_inst0.N_6_0_0 ;
    wire \DUT.uart_inst0.N_6_0_0_cascade_ ;
    wire \DUT.uart_inst0.N_15_mux_0 ;
    wire \DUT.uart_inst0.recv_state_ns_0_i_a2_0_2_3_cascade_ ;
    wire \DUT.uart_inst0.m16_N_3L3_1_cascade_ ;
    wire \DUT.uart_inst0.rx_bits_remaining_RNO_4Z0Z_1 ;
    wire \DUT.uart_inst0.g0_i_a3_5_cascade_ ;
    wire \DUT.uart_inst0.g0_0_i_a3_0_3 ;
    wire \DUT.uart_inst0.g0_0_i_a3_0_4_cascade_ ;
    wire \DUT.uart_inst0.g0_0 ;
    wire \DUT.uart_inst0.g0_i_a3_0_5_cascade_ ;
    wire \DUT.uart_inst0.g0_i_a3_8 ;
    wire \DUT.uart_inst0.g0_i_a3_0_6 ;
    wire \DUT.uart_inst0.g0_i_a3_0_7_cascade_ ;
    wire \DUT.uart_inst0.N_6_0_cascade_ ;
    wire \DUT.uart_inst0.N_40 ;
    wire \DUT.uart_inst0.rx_bits_remainingZ0Z_3 ;
    wire \DUT.uart_inst0.rx_bits_remainingZ0Z_0 ;
    wire \DUT.uart_inst0.recv_state_RNIL139CZ0Z_2 ;
    wire \DUT.uart_inst0.N_35_0 ;
    wire \DUT.uart_inst0.g0_0_2_cascade_ ;
    wire \DUT.uart_inst0.rx_bits_remainingZ0Z_2 ;
    wire \DUT.uart_inst0.m8_e_3 ;
    wire \DUT.uart_inst0.rx_bits_remainingZ0Z_1 ;
    wire \DUT.uart_inst0.g0_i_a3_6 ;
    wire \DUT.uart_inst0.recv_state_ns_0_i_a2_0_0_3 ;
    wire \DUT.uart_inst0.recv_stateZ0Z_3 ;
    wire \DUT.uart_inst0.g0_0_0 ;
    wire \DUT.uart_inst0.g0_0_1 ;
    wire \DUT.uart_inst0.N_81_mux_i_i_a5_0_4_0_cascade_ ;
    wire \DUT.uart_inst0.N_81_mux_i_i_a5_0_4 ;
    wire \DUT.uart_inst0.N_81_mux_i_i_0 ;
    wire \DUT.uart_inst0.N_81_mux_i_i_a5_0_5_cascade_ ;
    wire \DUT.uart_inst0.N_81_mux_i_i_a5_1_5 ;
    wire \DUT.uart_inst0.m8_e_2 ;
    wire bfn_8_15_0_;
    wire \DUT.uart_inst0.rx_countdown_3_cry_0_s1 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_1_s1 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_2_s1 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_3_s1 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_4_s1 ;
    wire \DUT.uart_inst0.m9_3 ;
    wire \DUT.uart_inst0.m9_4 ;
    wire \DUT.uart_inst0.N_8 ;
    wire \DUT.uart_inst0.N_81_mux_i_i_0_0 ;
    wire \DUT.uart_inst0.N_81_mux_i_i_a5_0_5_0 ;
    wire \DUT.uart_inst0.m4_3_cascade_ ;
    wire \DUT.uart_inst0.N_18_mux ;
    wire \DUT.uart_inst0.N_297_cascade_ ;
    wire \DUT.uart_inst0.recv_stateZ0Z_1 ;
    wire \DUT.uart_inst0.N_15_3 ;
    wire \DUT.uart_inst0.g0_0_i_a3_3_cascade_ ;
    wire \DUT.uart_inst0.g0_0_i_a3_4 ;
    wire \DUT.uart_inst0.recv_stateZ0Z_2 ;
    wire wPllLocked_i;
    wire bfn_8_18_0_;
    wire \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0 ;
    wire \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_awe3_cascade_ ;
    wire \DUT.fifo_rx_inst.un1_i11_i_cascade_ ;
    wire \DUT.fifo_rx_inst.un1_rFifoCount_1_axb_2 ;
    wire \DUT.fifo_rx_inst.un1_i11_i ;
    wire \DUT.fifo_rx_inst.rFifoCount_RNIK3G92Z0Z_1 ;
    wire \DUT.fifo_rx_inst.rWritePtr16_cascade_ ;
    wire \DUT.fifo_rx_inst.rWritePtr16 ;
    wire \DUT.fifo_rx_inst.rWritePtrZ0Z_0 ;
    wire \DUT.fifo_rx_inst.rWritePtrZ0Z_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_2 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_6 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_4 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_4 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_5 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_5 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_6 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_3 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_3 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_7 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_2 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_2 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_3 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_4 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_5 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_6 ;
    wire \DUT.uart_inst0.N_81_mux_i_i_a5_1_4 ;
    wire \DUT.uart_inst0.N_13_0 ;
    wire \DUT.uart_inst0.rx_countdown_RNO_2Z0Z_2 ;
    wire \DUT.uart_inst0.G_21_0_1_0_cascade_ ;
    wire \DUT.uart_inst0.G_9_i_o4_0 ;
    wire \DUT.uart_inst0.g0_0_3 ;
    wire \DUT.uart_inst0.G_16_i_a3_0_2_cascade_ ;
    wire \DUT.uart_inst0.N_45_cascade_ ;
    wire \DUT.uart_inst0.N_55 ;
    wire \DUT.uart_inst0.rx_countdown_3_s1_4 ;
    wire \DUT.uart_inst0.N_10 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_0_cascade_ ;
    wire \DUT.uart_inst0.G_21_0_1 ;
    wire \DUT.uart_inst0.recv_stateZ0Z_4 ;
    wire \DUT.uart_inst0.N_45 ;
    wire \DUT.uart_inst0.recv_state_ns_0_0_0 ;
    wire \DUT.uart_inst0.rx_countdown_3_s1_2 ;
    wire \DUT.uart_inst0.G_16_i_a3_0_3 ;
    wire \DUT.uart_inst0.g1_1 ;
    wire \DUT.uart_inst0.rx_countdown_3_s1_1 ;
    wire \DUT.uart_inst0.N_81_mux_i_i_a5_1_5_0 ;
    wire \DUT.uart_inst0.N_81_mux_i_i_a5_1_3 ;
    wire \DUT.uart_inst0.rx_countdown_3_s1_3 ;
    wire \DUT.uart_inst0.N_300_cascade_ ;
    wire \DUT.uart_inst0.G_16_i_a3_3_cascade_ ;
    wire \DUT.uart_inst0.G_16_i_a3_4 ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_1 ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_5 ;
    wire \DUT.uart_inst0.N_11_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_awe3_cascade_ ;
    wire \DUT.fifo_tx_inst.un1_i11_i ;
    wire \DUT.fifo_tx_inst.un1_i11_i_cascade_ ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_4 ;
    wire \DUT.uart_inst0.rx_countdownZ1Z_3 ;
    wire \DUT.uart_inst0.N_13_mux ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_2 ;
    wire \DUT.uart_inst0.rx_countdown_3_s1_5 ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_3 ;
    wire \DUT.uart_inst0.N_8_0_cascade_ ;
    wire \DUT.uart_inst0.m10_0_1 ;
    wire \DUT.uart_inst0.m11_0 ;
    wire \DUT.uart_inst0.N_15_mux ;
    wire \DUT.uart_inst0.N_11_0_cascade_ ;
    wire \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa ;
    wire \DUT.fifo_rx_inst.N_87_cascade_ ;
    wire \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0 ;
    wire \DUT.wRcvd ;
    wire \DUT.fifo_rx_inst.N_87 ;
    wire \DUT.fifo_rx_inst.N_92_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoCountZ0Z_0 ;
    wire \DUT.fifo_rx_inst.rFifoCountZ0Z_2 ;
    wire \DUT.fifo_rx_inst.rFifoCountZ0Z_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_awe2 ;
    wire \DUT.fifo_tx_inst.rFifoData_awe2_cascade_ ;
    wire \DUT.fifo_tx_inst.rFifoDataro_3 ;
    wire \DUT.fifo_tx_inst.rFifoDataro_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_awe0_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoDataro_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_awe1 ;
    wire \DUT.fifo_rx_inst.rFifoDataro_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_awe2 ;
    wire \DUT.fifo_rx_inst.rFifoDataro_3 ;
    wire \DUT.fifo_rx_inst.rFifoDataro_2 ;
    wire \DUT.fifo_rx_inst.rTxByte_42_1 ;
    wire \DUT.fifo_rx_inst.rTxByte_42_0_cascade_ ;
    wire N_92_i;
    wire rFifoDatarff_0_RNIHJV05_cascade_;
    wire \DUT.wRxByte_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_0 ;
    wire \DUT.wRxByte_1 ;
    wire \DUT.wRxByte_2 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_2 ;
    wire \DUT.wRxByte_3 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_3 ;
    wire \DUT.wRxByte_4 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_4 ;
    wire \DUT.wRxByte_5 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_5 ;
    wire \DUT.wRxByte_6 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_6 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_7 ;
    wire \DUT.fifo_rx_inst.rFifoData_awe3 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_7 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7 ;
    wire P1A3_c;
    wire \fifo_inst.ft2232h_inst.rFifoStateZ0Z_1 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_10 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_0 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_11 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_12 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_9 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_13 ;
    wire \DUT.uart_inst0.un1_N_5_mux_cascade_ ;
    wire \DUT.uart_inst0.g0_i_o6_0_4_cascade_ ;
    wire \DUT.uart_inst0.g0_i_o6_0_5 ;
    wire \DUT.uart_inst0.N_139_0_cascade_ ;
    wire \DUT.uart_inst0.tx_bits_remaining_RNO_1Z0Z_3 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_1 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_2 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_3 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_4 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_5 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_6 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_7 ;
    wire \DUT.uart_inst0.N_22_i ;
    wire \DUT.uart_inst0.N_79_cascade_ ;
    wire \DUT.uart_inst0.tx_state_ns_i_i_0_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_ ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_2 ;
    wire \DUT.rFifoDatarx_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_3 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ;
    wire \DUT.rFifoDatarx_3 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_3 ;
    wire \DUT.fifo_tx_inst.rFifoDataro_0 ;
    wire \DUT.fifo_tx_inst.rFifoDataro_1 ;
    wire \DUT.rFifoDataror_1 ;
    wire \DUT.rFifoDataror_1_cascade_ ;
    wire \DUT.rFifoDataror_0_0 ;
    wire \DUT.rFifoDataror_0 ;
    wire wPllLocked;
    wire \DUT.fifo_rx_inst.CO0 ;
    wire \DUT.fifo_rx_inst.un1_i11_2_i ;
    wire \DUT.fifo_rx_inst.un1_i11_2_i_cascade_ ;
    wire \DUT.fifo_rx_inst.N_92 ;
    wire \DUT.fifo_rx_inst.rReadPtrZ0Z_0 ;
    wire \DUT.fifo_tx_inst.rWritePtrZ0Z_0 ;
    wire \DUT.fifo_tx_inst.rWritePtrZ0Z_1 ;
    wire \DUT.fifo_tx_inst.N_83_cascade_ ;
    wire \DUT.fifo_tx_inst.N_88 ;
    wire \DUT.fifo_tx_inst.N_88_cascade_ ;
    wire \DUT.rTransmitc ;
    wire \DUT.fifo_tx_inst.rWritePtr16 ;
    wire \DUT.fifo_tx_inst.un1_i11_2_i ;
    wire \DUT.fifo_rx_inst.rReadPtrZ0Z_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1 ;
    wire N_92_i_0;
    wire rFifoDatarff_0_RNIHJV05;
    wire \fifo_inst.ft2232h_inst.rFifoStateZ0Z_2 ;
    wire P1A4_c;
    wire \fifo_inst.ft2232h_inst.rFifoStateZ0Z_3 ;
    wire rTxBusReady;
    wire \fifo_inst.ft2232h_inst.rFifoStateZ0Z_4 ;
    wire \fifo_inst.ft2232h_inst.rTxRdEnZ0 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_1 ;
    wire bfn_11_13_0_;
    wire \DUT.uart_inst0.rx_clk_dividerZ1Z_1 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_0 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_1 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_3 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_2_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_2 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_3 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_5 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_4_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_4 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_6 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_5_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_5 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_7 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_6 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_7 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_8 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO ;
    wire bfn_11_14_0_;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_9 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_8 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_10 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_9 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_11 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_10 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_11 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_13 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_12 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_14 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_13 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_15 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_14 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_15 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_16 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO ;
    wire bfn_11_15_0_;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_16 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_17 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_12 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_2 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO ;
    wire \DUT.uart_inst0.N_50 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_4 ;
    wire \DUT.uart_inst0.N_98_cascade_ ;
    wire P1A7_c;
    wire \DUT.uart_inst0.N_82 ;
    wire \DUT.uart_inst0.N_99 ;
    wire \DUT.uart_inst0.N_100 ;
    wire P1A1_c;
    wire \DUT.uart_inst0.recv_stateZ0Z_5 ;
    wire \DUT.uart_inst0.recv_stateZ0Z_0 ;
    wire \DUT.uart_inst0.N_49 ;
    wire \fifo_inst.ft2232h_inst.rFifoStatec_0 ;
    wire \DUT.uart_inst0.tx_bits_remainingZ0Z_3 ;
    wire \DUT.uart_inst0.N_139 ;
    wire \DUT.uart_inst0.tx_bits_remainingZ0Z_2 ;
    wire \DUT.rTransmitc_0 ;
    wire \DUT.uart_inst0.N_85_cascade_ ;
    wire \DUT.uart_inst0.N_66 ;
    wire \DUT.uart_inst0.N_22_cascade_ ;
    wire \DUT.uart_inst0.tx_bits_remainingZ0Z_0 ;
    wire \DUT.uart_inst0.N_22 ;
    wire \DUT.uart_inst0.tx_bits_remainingZ0Z_1 ;
    wire \DUT.uart_inst0.N_65_i ;
    wire \DUT.uart_inst0.tx_dataZ0Z_0 ;
    wire \DUT.uart_inst0.N_85 ;
    wire \DUT.uart_inst0.N_89 ;
    wire bfn_11_18_0_;
    wire \DUT.uart_inst0.tx_clk_divider_cry_0 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_1 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_2 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_3 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_4 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_5 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_6 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_7 ;
    wire bfn_11_19_0_;
    wire \DUT.uart_inst0.tx_clk_divider_cry_8 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_9 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_10 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_11 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_12 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_7 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_ ;
    wire \DUT.rFifoDatarx_7 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_7 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_0 ;
    wire \DUT.rFifoDatarxZ0Z_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1_cascade_ ;
    wire \DUT.rFifoDatarx_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_ ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_4 ;
    wire \DUT.rFifoDatarx_4 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_4 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_5 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ;
    wire \DUT.rFifoDatarx_5 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_5 ;
    wire \DUT.fifo_tx_inst.rReadPtrZ0Z_0 ;
    wire \DUT.fifo_tx_inst.rReadPtrZ0Z_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_ ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_6 ;
    wire \DUT.rFifoDatarx_6 ;
    wire \DUT.rFifoCount_0 ;
    wire \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0 ;
    wire bfn_11_22_0_;
    wire \DUT.fifo_tx_inst.rFifoCount_RNIBPFMZ0Z_1 ;
    wire \DUT.rFifoCount_1 ;
    wire \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0 ;
    wire rRxReadZ0;
    wire \DUT.fifo_tx_inst.N_83 ;
    wire \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1 ;
    wire \DUT.rFifoCount_2 ;
    wire wPllLocked_i_g;
    wire \DUT.wRxByte_7 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_7 ;
    wire \DUT.fifo_rx_inst.rFifoData_awe0 ;
    wire iRxF_n_c;
    wire iTxE_n_c;
    wire \fifo_inst.ft2232h_inst.rFifoStateZ0Z_0 ;
    wire \fifo_inst.ft2232h_inst.N_101 ;
    wire \DUT.uart_inst0.N_13_cascade_ ;
    wire \DUT.uart_inst0.g0_i_0_cascade_ ;
    wire \DUT.uart_inst0.g0_i_a6_0 ;
    wire \DUT.uart_inst0.g0_i_1_cascade_ ;
    wire \DUT.uart_inst0.g0_i_a6_3_0 ;
    wire \DUT.uart_inst0.g0_i_o2_1_cascade_ ;
    wire \DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0_cascade_ ;
    wire \DUT.uart_inst0.N_77 ;
    wire \DUT.uart_inst0.g0_i_o2_2 ;
    wire \DUT.uart_inst0.g0_i_o2_3 ;
    wire \DUT.uart_inst0.N_11 ;
    wire \DUT.uart_inst0.g0_11_a4_2 ;
    wire \DUT.uart_inst0.N_9 ;
    wire \DUT.uart_inst0.tx_state_ns_i_i_o2_a0_2_0_cascade_ ;
    wire \DUT.uart_inst0.N_71_i ;
    wire \DUT.uart_inst0.N_8_1 ;
    wire \DUT.uart_inst0.g0_i_a3_0_cascade_ ;
    wire wPllLocked_g;
    wire \DUT.uart_inst0.tx_countdownZ0Z_4 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_3 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_5 ;
    wire \DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0 ;
    wire \DUT.uart_inst0.g0_11_a3_2_cascade_ ;
    wire \DUT.uart_inst0.N_7 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_1 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_2 ;
    wire \DUT.uart_inst0.N_6_i ;
    wire \DUT.rTransmitZ0 ;
    wire \DUT.tx_state_0 ;
    wire \DUT.uart_inst0.tx_stateZ0Z_1 ;
    wire \DUT.uart_inst0.N_11_1 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_9 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_10 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_11 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_8 ;
    wire \DUT.uart_inst0.N_20 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_1 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_0 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_2 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_4 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_5 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_3 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_12 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_7 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_13 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_6 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_9 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_7 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_8_cascade_ ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_6 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_0 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_0 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_0_cascade_ ;
    wire \DUT.uart_inst0.N_5_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_3 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_4 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_5 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_6 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_7 ;
    wire \DUT.fifo_tx_inst.rFifoData_awe3 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_1 ;
    wire rTxByteZ0Z_2;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_2 ;
    wire rTxByteZ0Z_3;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_3 ;
    wire rTxByteZ0Z_4;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_4 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_6 ;
    wire rTxByteZ0Z_7;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_7 ;
    wire rTxByteZ0Z_1;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_1 ;
    wire rTxByteZ0Z_6;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_6 ;
    wire \DUT.fifo_tx_inst.rFifoData_awe0 ;
    wire rTxByteZ0Z_5;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_5 ;
    wire rTxByteZ0Z_0;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_0 ;
    wire clk_48mhz;
    wire \DUT.fifo_tx_inst.rFifoData_awe1 ;
    wire CONSTANT_ONE_NET;
    wire _gnd_net_;

    defparam \top_pll_inst.top_pll_inst_pll .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \top_pll_inst.top_pll_inst_pll .TEST_MODE=1'b0;
    defparam \top_pll_inst.top_pll_inst_pll .SHIFTREG_DIV_MODE=2'b00;
    defparam \top_pll_inst.top_pll_inst_pll .PLLOUT_SELECT="GENCLK";
    defparam \top_pll_inst.top_pll_inst_pll .FILTER_RANGE=3'b001;
    defparam \top_pll_inst.top_pll_inst_pll .FEEDBACK_PATH="SIMPLE";
    defparam \top_pll_inst.top_pll_inst_pll .FDA_RELATIVE=4'b0000;
    defparam \top_pll_inst.top_pll_inst_pll .FDA_FEEDBACK=4'b0000;
    defparam \top_pll_inst.top_pll_inst_pll .ENABLE_ICEGATE=1'b0;
    defparam \top_pll_inst.top_pll_inst_pll .DIVR=4'b0000;
    defparam \top_pll_inst.top_pll_inst_pll .DIVQ=3'b100;
    defparam \top_pll_inst.top_pll_inst_pll .DIVF=7'b0111111;
    defparam \top_pll_inst.top_pll_inst_pll .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    PLL40 \top_pll_inst.top_pll_inst_pll  (
            .PLLOUTGLOBAL(clk_48mhz),
            .SDI(GNDG0),
            .BYPASS(GNDG0),
            .RESETB(N__5081),
            .PLLOUTCORE(),
            .LOCK(\PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO ),
            .SDO(),
            .SCLK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .EXTFEEDBACK(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLIN(N__13526));
    IO_PAD \top_pll_inst.top_pll_inst_iopad  (
            .OE(VCCG0),
            .DIN(),
            .DOUT(N__13526),
            .PACKAGEPIN(iClk));
    IO_PAD P1A8_obuft_iopad (
            .OE(N__13512),
            .DIN(N__13511),
            .DOUT(N__13510),
            .PACKAGEPIN(P1A8));
    defparam P1A8_obuft_preio.NEG_TRIGGER=1'b0;
    defparam P1A8_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO P1A8_obuft_preio (
            .PADOEN(N__13512),
            .PADOUT(N__13511),
            .PADIN(N__13510),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_1_iopad (
            .OE(N__13503),
            .DIN(N__13502),
            .DOUT(N__13501),
            .PACKAGEPIN(ioFifoData[1]));
    defparam ioFifoData_obuft_1_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_1_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_1_preio (
            .PADOEN(N__13503),
            .PADOUT(N__13502),
            .PADIN(N__13501),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8698),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A9_obuft_iopad (
            .OE(N__13494),
            .DIN(N__13493),
            .DOUT(N__13492),
            .PACKAGEPIN(P1A9));
    defparam P1A9_obuft_preio.NEG_TRIGGER=1'b0;
    defparam P1A9_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO P1A9_obuft_preio (
            .PADOEN(N__13494),
            .PADOUT(N__13493),
            .PADIN(N__13492),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_4_iopad (
            .OE(N__13485),
            .DIN(N__13484),
            .DOUT(N__13483),
            .PACKAGEPIN(ioFifoData[4]));
    defparam ioFifoData_obuft_4_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_4_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_4_preio (
            .PADOEN(N__13485),
            .PADOUT(N__13484),
            .PADIN(N__13483),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8743),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A2_obuft_iopad (
            .OE(N__13476),
            .DIN(N__13475),
            .DOUT(N__13474),
            .PACKAGEPIN(P1A2));
    defparam P1A2_obuft_preio.NEG_TRIGGER=1'b0;
    defparam P1A2_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO P1A2_obuft_preio (
            .PADOEN(N__13476),
            .PADOUT(N__13475),
            .PADIN(N__13474),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A4_obuf_iopad (
            .OE(N__13467),
            .DIN(N__13466),
            .DOUT(N__13465),
            .PACKAGEPIN(P1A4));
    defparam P1A4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO P1A4_obuf_preio (
            .PADOEN(N__13467),
            .PADOUT(N__13466),
            .PADIN(N__13465),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8800),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_0_iopad (
            .OE(N__13458),
            .DIN(N__13457),
            .DOUT(N__13456),
            .PACKAGEPIN(ioFifoData[0]));
    defparam ioFifoData_obuft_0_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_0_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_0_preio (
            .PADOEN(N__13458),
            .PADOUT(N__13457),
            .PADIN(N__13456),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8722),
            .DIN0(),
            .DOUT0(N__12841),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD oRx_n_obuf_iopad (
            .OE(N__13449),
            .DIN(N__13448),
            .DOUT(N__13447),
            .PACKAGEPIN(oRx_n));
    defparam oRx_n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam oRx_n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO oRx_n_obuf_preio (
            .PADOEN(N__13449),
            .PADOUT(N__13448),
            .PADIN(N__13447),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7550),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_7_iopad (
            .OE(N__13440),
            .DIN(N__13439),
            .DOUT(N__13438),
            .PACKAGEPIN(ioFifoData[7]));
    defparam ioFifoData_obuft_7_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_7_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_7_preio (
            .PADOEN(N__13440),
            .PADOUT(N__13439),
            .PADIN(N__13438),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8751),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD iRxF_n_ibuf_iopad (
            .OE(N__13431),
            .DIN(N__13430),
            .DOUT(N__13429),
            .PACKAGEPIN(iRxF_n));
    defparam iRxF_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam iRxF_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO iRxF_n_ibuf_preio (
            .PADOEN(N__13431),
            .PADOUT(N__13430),
            .PADIN(N__13429),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(iRxF_n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A3_obuf_iopad (
            .OE(N__13422),
            .DIN(N__13421),
            .DOUT(N__13420),
            .PACKAGEPIN(P1A3));
    defparam P1A3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO P1A3_obuf_preio (
            .PADOEN(N__13422),
            .PADOUT(N__13421),
            .PADIN(N__13420),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7546),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A7_obuf_iopad (
            .OE(N__13413),
            .DIN(N__13412),
            .DOUT(N__13411),
            .PACKAGEPIN(P1A7));
    defparam P1A7_obuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A7_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO P1A7_obuf_preio (
            .PADOEN(N__13413),
            .PADOUT(N__13412),
            .PADIN(N__13411),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9461),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BTN_N_ibuf_iopad (
            .OE(N__13404),
            .DIN(N__13403),
            .DOUT(N__13402),
            .PACKAGEPIN(BTN_N));
    defparam BTN_N_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam BTN_N_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO BTN_N_ibuf_preio (
            .PADOEN(N__13404),
            .PADOUT(N__13403),
            .PADIN(N__13402),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(BTN_N_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_3_iopad (
            .OE(N__13395),
            .DIN(N__13394),
            .DOUT(N__13393),
            .PACKAGEPIN(ioFifoData[3]));
    defparam ioFifoData_obuft_3_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_3_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_3_preio (
            .PADOEN(N__13395),
            .PADOUT(N__13394),
            .PADIN(N__13393),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8752),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_6_iopad (
            .OE(N__13386),
            .DIN(N__13385),
            .DOUT(N__13384),
            .PACKAGEPIN(ioFifoData[6]));
    defparam ioFifoData_obuft_6_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_6_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_6_preio (
            .PADOEN(N__13386),
            .PADOUT(N__13385),
            .PADIN(N__13384),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8750),
            .DIN0(),
            .DOUT0(N__12840),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_5_iopad (
            .OE(N__13377),
            .DIN(N__13376),
            .DOUT(N__13375),
            .PACKAGEPIN(ioFifoData[5]));
    defparam ioFifoData_obuft_5_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_5_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_5_preio (
            .PADOEN(N__13377),
            .PADOUT(N__13376),
            .PADIN(N__13375),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8728),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD oTx_n_obuf_iopad (
            .OE(N__13368),
            .DIN(N__13367),
            .DOUT(N__13366),
            .PACKAGEPIN(oTx_n));
    defparam oTx_n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam oTx_n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO oTx_n_obuf_preio (
            .PADOEN(N__13368),
            .PADOUT(N__13367),
            .PADIN(N__13366),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8804),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD iTxE_n_ibuf_iopad (
            .OE(N__13359),
            .DIN(N__13358),
            .DOUT(N__13357),
            .PACKAGEPIN(iTxE_n));
    defparam iTxE_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam iTxE_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO iTxE_n_ibuf_preio (
            .PADOEN(N__13359),
            .PADOUT(N__13358),
            .PADIN(N__13357),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(iTxE_n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_2_iopad (
            .OE(N__13350),
            .DIN(N__13349),
            .DOUT(N__13348),
            .PACKAGEPIN(ioFifoData[2]));
    defparam ioFifoData_obuft_2_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_2_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_2_preio (
            .PADOEN(N__13350),
            .PADOUT(N__13349),
            .PADIN(N__13348),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8753),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A1_ibuf_iopad (
            .OE(N__13341),
            .DIN(N__13340),
            .DOUT(N__13339),
            .PACKAGEPIN(P1A1));
    defparam P1A1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO P1A1_ibuf_preio (
            .PADOEN(N__13341),
            .PADOUT(N__13340),
            .PADIN(N__13339),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(P1A1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__3179 (
            .O(N__13322),
            .I(N__13316));
    InMux I__3178 (
            .O(N__13321),
            .I(N__13313));
    InMux I__3177 (
            .O(N__13320),
            .I(N__13310));
    InMux I__3176 (
            .O(N__13319),
            .I(N__13307));
    LocalMux I__3175 (
            .O(N__13316),
            .I(N__13302));
    LocalMux I__3174 (
            .O(N__13313),
            .I(N__13302));
    LocalMux I__3173 (
            .O(N__13310),
            .I(N__13299));
    LocalMux I__3172 (
            .O(N__13307),
            .I(N__13296));
    Span4Mux_v I__3171 (
            .O(N__13302),
            .I(N__13293));
    Span4Mux_v I__3170 (
            .O(N__13299),
            .I(N__13288));
    Span4Mux_v I__3169 (
            .O(N__13296),
            .I(N__13288));
    Odrv4 I__3168 (
            .O(N__13293),
            .I(rTxByteZ0Z_7));
    Odrv4 I__3167 (
            .O(N__13288),
            .I(rTxByteZ0Z_7));
    InMux I__3166 (
            .O(N__13283),
            .I(N__13280));
    LocalMux I__3165 (
            .O(N__13280),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_7 ));
    InMux I__3164 (
            .O(N__13277),
            .I(N__13271));
    InMux I__3163 (
            .O(N__13276),
            .I(N__13268));
    InMux I__3162 (
            .O(N__13275),
            .I(N__13265));
    InMux I__3161 (
            .O(N__13274),
            .I(N__13262));
    LocalMux I__3160 (
            .O(N__13271),
            .I(N__13259));
    LocalMux I__3159 (
            .O(N__13268),
            .I(N__13254));
    LocalMux I__3158 (
            .O(N__13265),
            .I(N__13254));
    LocalMux I__3157 (
            .O(N__13262),
            .I(N__13251));
    Span4Mux_v I__3156 (
            .O(N__13259),
            .I(N__13248));
    Span4Mux_v I__3155 (
            .O(N__13254),
            .I(N__13245));
    Span4Mux_h I__3154 (
            .O(N__13251),
            .I(N__13242));
    Odrv4 I__3153 (
            .O(N__13248),
            .I(rTxByteZ0Z_1));
    Odrv4 I__3152 (
            .O(N__13245),
            .I(rTxByteZ0Z_1));
    Odrv4 I__3151 (
            .O(N__13242),
            .I(rTxByteZ0Z_1));
    InMux I__3150 (
            .O(N__13235),
            .I(N__13232));
    LocalMux I__3149 (
            .O(N__13232),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_1 ));
    InMux I__3148 (
            .O(N__13229),
            .I(N__13225));
    InMux I__3147 (
            .O(N__13228),
            .I(N__13222));
    LocalMux I__3146 (
            .O(N__13225),
            .I(N__13217));
    LocalMux I__3145 (
            .O(N__13222),
            .I(N__13217));
    Span4Mux_v I__3144 (
            .O(N__13217),
            .I(N__13213));
    InMux I__3143 (
            .O(N__13216),
            .I(N__13210));
    Sp12to4 I__3142 (
            .O(N__13213),
            .I(N__13204));
    LocalMux I__3141 (
            .O(N__13210),
            .I(N__13204));
    InMux I__3140 (
            .O(N__13209),
            .I(N__13201));
    Odrv12 I__3139 (
            .O(N__13204),
            .I(rTxByteZ0Z_6));
    LocalMux I__3138 (
            .O(N__13201),
            .I(rTxByteZ0Z_6));
    InMux I__3137 (
            .O(N__13196),
            .I(N__13193));
    LocalMux I__3136 (
            .O(N__13193),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_6 ));
    CEMux I__3135 (
            .O(N__13190),
            .I(N__13184));
    CEMux I__3134 (
            .O(N__13189),
            .I(N__13181));
    CEMux I__3133 (
            .O(N__13188),
            .I(N__13178));
    CEMux I__3132 (
            .O(N__13187),
            .I(N__13175));
    LocalMux I__3131 (
            .O(N__13184),
            .I(N__13172));
    LocalMux I__3130 (
            .O(N__13181),
            .I(N__13169));
    LocalMux I__3129 (
            .O(N__13178),
            .I(N__13164));
    LocalMux I__3128 (
            .O(N__13175),
            .I(N__13164));
    Span4Mux_h I__3127 (
            .O(N__13172),
            .I(N__13161));
    Span4Mux_v I__3126 (
            .O(N__13169),
            .I(N__13158));
    Span4Mux_v I__3125 (
            .O(N__13164),
            .I(N__13153));
    Span4Mux_h I__3124 (
            .O(N__13161),
            .I(N__13153));
    Odrv4 I__3123 (
            .O(N__13158),
            .I(\DUT.fifo_tx_inst.rFifoData_awe0 ));
    Odrv4 I__3122 (
            .O(N__13153),
            .I(\DUT.fifo_tx_inst.rFifoData_awe0 ));
    InMux I__3121 (
            .O(N__13148),
            .I(N__13144));
    InMux I__3120 (
            .O(N__13147),
            .I(N__13141));
    LocalMux I__3119 (
            .O(N__13144),
            .I(N__13137));
    LocalMux I__3118 (
            .O(N__13141),
            .I(N__13134));
    InMux I__3117 (
            .O(N__13140),
            .I(N__13131));
    Span4Mux_v I__3116 (
            .O(N__13137),
            .I(N__13123));
    Span4Mux_v I__3115 (
            .O(N__13134),
            .I(N__13123));
    LocalMux I__3114 (
            .O(N__13131),
            .I(N__13123));
    InMux I__3113 (
            .O(N__13130),
            .I(N__13120));
    Odrv4 I__3112 (
            .O(N__13123),
            .I(rTxByteZ0Z_5));
    LocalMux I__3111 (
            .O(N__13120),
            .I(rTxByteZ0Z_5));
    InMux I__3110 (
            .O(N__13115),
            .I(N__13112));
    LocalMux I__3109 (
            .O(N__13112),
            .I(N__13109));
    Odrv4 I__3108 (
            .O(N__13109),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_5 ));
    InMux I__3107 (
            .O(N__13106),
            .I(N__13102));
    InMux I__3106 (
            .O(N__13105),
            .I(N__13099));
    LocalMux I__3105 (
            .O(N__13102),
            .I(N__13095));
    LocalMux I__3104 (
            .O(N__13099),
            .I(N__13092));
    InMux I__3103 (
            .O(N__13098),
            .I(N__13089));
    Span4Mux_v I__3102 (
            .O(N__13095),
            .I(N__13081));
    Span4Mux_h I__3101 (
            .O(N__13092),
            .I(N__13081));
    LocalMux I__3100 (
            .O(N__13089),
            .I(N__13081));
    InMux I__3099 (
            .O(N__13088),
            .I(N__13078));
    Span4Mux_h I__3098 (
            .O(N__13081),
            .I(N__13075));
    LocalMux I__3097 (
            .O(N__13078),
            .I(N__13072));
    Odrv4 I__3096 (
            .O(N__13075),
            .I(rTxByteZ0Z_0));
    Odrv4 I__3095 (
            .O(N__13072),
            .I(rTxByteZ0Z_0));
    CascadeMux I__3094 (
            .O(N__13067),
            .I(N__13064));
    InMux I__3093 (
            .O(N__13064),
            .I(N__13061));
    LocalMux I__3092 (
            .O(N__13061),
            .I(N__13058));
    Odrv4 I__3091 (
            .O(N__13058),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_0 ));
    ClkMux I__3090 (
            .O(N__13055),
            .I(N__12887));
    ClkMux I__3089 (
            .O(N__13054),
            .I(N__12887));
    ClkMux I__3088 (
            .O(N__13053),
            .I(N__12887));
    ClkMux I__3087 (
            .O(N__13052),
            .I(N__12887));
    ClkMux I__3086 (
            .O(N__13051),
            .I(N__12887));
    ClkMux I__3085 (
            .O(N__13050),
            .I(N__12887));
    ClkMux I__3084 (
            .O(N__13049),
            .I(N__12887));
    ClkMux I__3083 (
            .O(N__13048),
            .I(N__12887));
    ClkMux I__3082 (
            .O(N__13047),
            .I(N__12887));
    ClkMux I__3081 (
            .O(N__13046),
            .I(N__12887));
    ClkMux I__3080 (
            .O(N__13045),
            .I(N__12887));
    ClkMux I__3079 (
            .O(N__13044),
            .I(N__12887));
    ClkMux I__3078 (
            .O(N__13043),
            .I(N__12887));
    ClkMux I__3077 (
            .O(N__13042),
            .I(N__12887));
    ClkMux I__3076 (
            .O(N__13041),
            .I(N__12887));
    ClkMux I__3075 (
            .O(N__13040),
            .I(N__12887));
    ClkMux I__3074 (
            .O(N__13039),
            .I(N__12887));
    ClkMux I__3073 (
            .O(N__13038),
            .I(N__12887));
    ClkMux I__3072 (
            .O(N__13037),
            .I(N__12887));
    ClkMux I__3071 (
            .O(N__13036),
            .I(N__12887));
    ClkMux I__3070 (
            .O(N__13035),
            .I(N__12887));
    ClkMux I__3069 (
            .O(N__13034),
            .I(N__12887));
    ClkMux I__3068 (
            .O(N__13033),
            .I(N__12887));
    ClkMux I__3067 (
            .O(N__13032),
            .I(N__12887));
    ClkMux I__3066 (
            .O(N__13031),
            .I(N__12887));
    ClkMux I__3065 (
            .O(N__13030),
            .I(N__12887));
    ClkMux I__3064 (
            .O(N__13029),
            .I(N__12887));
    ClkMux I__3063 (
            .O(N__13028),
            .I(N__12887));
    ClkMux I__3062 (
            .O(N__13027),
            .I(N__12887));
    ClkMux I__3061 (
            .O(N__13026),
            .I(N__12887));
    ClkMux I__3060 (
            .O(N__13025),
            .I(N__12887));
    ClkMux I__3059 (
            .O(N__13024),
            .I(N__12887));
    ClkMux I__3058 (
            .O(N__13023),
            .I(N__12887));
    ClkMux I__3057 (
            .O(N__13022),
            .I(N__12887));
    ClkMux I__3056 (
            .O(N__13021),
            .I(N__12887));
    ClkMux I__3055 (
            .O(N__13020),
            .I(N__12887));
    ClkMux I__3054 (
            .O(N__13019),
            .I(N__12887));
    ClkMux I__3053 (
            .O(N__13018),
            .I(N__12887));
    ClkMux I__3052 (
            .O(N__13017),
            .I(N__12887));
    ClkMux I__3051 (
            .O(N__13016),
            .I(N__12887));
    ClkMux I__3050 (
            .O(N__13015),
            .I(N__12887));
    ClkMux I__3049 (
            .O(N__13014),
            .I(N__12887));
    ClkMux I__3048 (
            .O(N__13013),
            .I(N__12887));
    ClkMux I__3047 (
            .O(N__13012),
            .I(N__12887));
    ClkMux I__3046 (
            .O(N__13011),
            .I(N__12887));
    ClkMux I__3045 (
            .O(N__13010),
            .I(N__12887));
    ClkMux I__3044 (
            .O(N__13009),
            .I(N__12887));
    ClkMux I__3043 (
            .O(N__13008),
            .I(N__12887));
    ClkMux I__3042 (
            .O(N__13007),
            .I(N__12887));
    ClkMux I__3041 (
            .O(N__13006),
            .I(N__12887));
    ClkMux I__3040 (
            .O(N__13005),
            .I(N__12887));
    ClkMux I__3039 (
            .O(N__13004),
            .I(N__12887));
    ClkMux I__3038 (
            .O(N__13003),
            .I(N__12887));
    ClkMux I__3037 (
            .O(N__13002),
            .I(N__12887));
    ClkMux I__3036 (
            .O(N__13001),
            .I(N__12887));
    ClkMux I__3035 (
            .O(N__13000),
            .I(N__12887));
    GlobalMux I__3034 (
            .O(N__12887),
            .I(clk_48mhz));
    CEMux I__3033 (
            .O(N__12884),
            .I(N__12880));
    CEMux I__3032 (
            .O(N__12883),
            .I(N__12876));
    LocalMux I__3031 (
            .O(N__12880),
            .I(N__12873));
    CEMux I__3030 (
            .O(N__12879),
            .I(N__12870));
    LocalMux I__3029 (
            .O(N__12876),
            .I(N__12867));
    Span4Mux_v I__3028 (
            .O(N__12873),
            .I(N__12862));
    LocalMux I__3027 (
            .O(N__12870),
            .I(N__12862));
    Span4Mux_h I__3026 (
            .O(N__12867),
            .I(N__12856));
    Span4Mux_v I__3025 (
            .O(N__12862),
            .I(N__12856));
    InMux I__3024 (
            .O(N__12861),
            .I(N__12853));
    Odrv4 I__3023 (
            .O(N__12856),
            .I(\DUT.fifo_tx_inst.rFifoData_awe1 ));
    LocalMux I__3022 (
            .O(N__12853),
            .I(\DUT.fifo_tx_inst.rFifoData_awe1 ));
    CascadeMux I__3021 (
            .O(N__12848),
            .I(N__12837));
    CascadeMux I__3020 (
            .O(N__12847),
            .I(N__12834));
    CascadeMux I__3019 (
            .O(N__12846),
            .I(N__12831));
    CascadeMux I__3018 (
            .O(N__12845),
            .I(N__12828));
    CascadeMux I__3017 (
            .O(N__12844),
            .I(N__12825));
    CascadeMux I__3016 (
            .O(N__12843),
            .I(N__12822));
    CascadeMux I__3015 (
            .O(N__12842),
            .I(N__12819));
    IoInMux I__3014 (
            .O(N__12841),
            .I(N__12808));
    IoInMux I__3013 (
            .O(N__12840),
            .I(N__12804));
    InMux I__3012 (
            .O(N__12837),
            .I(N__12797));
    InMux I__3011 (
            .O(N__12834),
            .I(N__12797));
    InMux I__3010 (
            .O(N__12831),
            .I(N__12797));
    InMux I__3009 (
            .O(N__12828),
            .I(N__12788));
    InMux I__3008 (
            .O(N__12825),
            .I(N__12788));
    InMux I__3007 (
            .O(N__12822),
            .I(N__12788));
    InMux I__3006 (
            .O(N__12819),
            .I(N__12788));
    CascadeMux I__3005 (
            .O(N__12818),
            .I(N__12785));
    CascadeMux I__3004 (
            .O(N__12817),
            .I(N__12782));
    CascadeMux I__3003 (
            .O(N__12816),
            .I(N__12779));
    CascadeMux I__3002 (
            .O(N__12815),
            .I(N__12776));
    CascadeMux I__3001 (
            .O(N__12814),
            .I(N__12773));
    CascadeMux I__3000 (
            .O(N__12813),
            .I(N__12770));
    CascadeMux I__2999 (
            .O(N__12812),
            .I(N__12767));
    CascadeMux I__2998 (
            .O(N__12811),
            .I(N__12764));
    LocalMux I__2997 (
            .O(N__12808),
            .I(N__12753));
    CascadeMux I__2996 (
            .O(N__12807),
            .I(N__12748));
    LocalMux I__2995 (
            .O(N__12804),
            .I(N__12744));
    LocalMux I__2994 (
            .O(N__12797),
            .I(N__12736));
    LocalMux I__2993 (
            .O(N__12788),
            .I(N__12736));
    InMux I__2992 (
            .O(N__12785),
            .I(N__12727));
    InMux I__2991 (
            .O(N__12782),
            .I(N__12727));
    InMux I__2990 (
            .O(N__12779),
            .I(N__12727));
    InMux I__2989 (
            .O(N__12776),
            .I(N__12727));
    InMux I__2988 (
            .O(N__12773),
            .I(N__12718));
    InMux I__2987 (
            .O(N__12770),
            .I(N__12718));
    InMux I__2986 (
            .O(N__12767),
            .I(N__12718));
    InMux I__2985 (
            .O(N__12764),
            .I(N__12718));
    CascadeMux I__2984 (
            .O(N__12763),
            .I(N__12715));
    CascadeMux I__2983 (
            .O(N__12762),
            .I(N__12712));
    CascadeMux I__2982 (
            .O(N__12761),
            .I(N__12709));
    CascadeMux I__2981 (
            .O(N__12760),
            .I(N__12706));
    CascadeMux I__2980 (
            .O(N__12759),
            .I(N__12703));
    CascadeMux I__2979 (
            .O(N__12758),
            .I(N__12699));
    CascadeMux I__2978 (
            .O(N__12757),
            .I(N__12696));
    CascadeMux I__2977 (
            .O(N__12756),
            .I(N__12692));
    IoSpan4Mux I__2976 (
            .O(N__12753),
            .I(N__12689));
    InMux I__2975 (
            .O(N__12752),
            .I(N__12686));
    InMux I__2974 (
            .O(N__12751),
            .I(N__12679));
    InMux I__2973 (
            .O(N__12748),
            .I(N__12679));
    InMux I__2972 (
            .O(N__12747),
            .I(N__12679));
    Span4Mux_s0_v I__2971 (
            .O(N__12744),
            .I(N__12676));
    CascadeMux I__2970 (
            .O(N__12743),
            .I(N__12673));
    CascadeMux I__2969 (
            .O(N__12742),
            .I(N__12670));
    CascadeMux I__2968 (
            .O(N__12741),
            .I(N__12667));
    Span4Mux_v I__2967 (
            .O(N__12736),
            .I(N__12660));
    LocalMux I__2966 (
            .O(N__12727),
            .I(N__12660));
    LocalMux I__2965 (
            .O(N__12718),
            .I(N__12660));
    InMux I__2964 (
            .O(N__12715),
            .I(N__12657));
    InMux I__2963 (
            .O(N__12712),
            .I(N__12648));
    InMux I__2962 (
            .O(N__12709),
            .I(N__12648));
    InMux I__2961 (
            .O(N__12706),
            .I(N__12648));
    InMux I__2960 (
            .O(N__12703),
            .I(N__12648));
    InMux I__2959 (
            .O(N__12702),
            .I(N__12637));
    InMux I__2958 (
            .O(N__12699),
            .I(N__12637));
    InMux I__2957 (
            .O(N__12696),
            .I(N__12637));
    InMux I__2956 (
            .O(N__12695),
            .I(N__12637));
    InMux I__2955 (
            .O(N__12692),
            .I(N__12637));
    Span4Mux_s2_v I__2954 (
            .O(N__12689),
            .I(N__12633));
    LocalMux I__2953 (
            .O(N__12686),
            .I(N__12628));
    LocalMux I__2952 (
            .O(N__12679),
            .I(N__12628));
    Span4Mux_h I__2951 (
            .O(N__12676),
            .I(N__12625));
    InMux I__2950 (
            .O(N__12673),
            .I(N__12618));
    InMux I__2949 (
            .O(N__12670),
            .I(N__12618));
    InMux I__2948 (
            .O(N__12667),
            .I(N__12618));
    Span4Mux_h I__2947 (
            .O(N__12660),
            .I(N__12611));
    LocalMux I__2946 (
            .O(N__12657),
            .I(N__12611));
    LocalMux I__2945 (
            .O(N__12648),
            .I(N__12611));
    LocalMux I__2944 (
            .O(N__12637),
            .I(N__12608));
    InMux I__2943 (
            .O(N__12636),
            .I(N__12605));
    Sp12to4 I__2942 (
            .O(N__12633),
            .I(N__12602));
    Sp12to4 I__2941 (
            .O(N__12628),
            .I(N__12599));
    Span4Mux_v I__2940 (
            .O(N__12625),
            .I(N__12596));
    LocalMux I__2939 (
            .O(N__12618),
            .I(N__12587));
    Span4Mux_v I__2938 (
            .O(N__12611),
            .I(N__12587));
    Span4Mux_v I__2937 (
            .O(N__12608),
            .I(N__12587));
    LocalMux I__2936 (
            .O(N__12605),
            .I(N__12587));
    Span12Mux_s10_v I__2935 (
            .O(N__12602),
            .I(N__12584));
    Span12Mux_v I__2934 (
            .O(N__12599),
            .I(N__12581));
    Span4Mux_v I__2933 (
            .O(N__12596),
            .I(N__12576));
    Span4Mux_h I__2932 (
            .O(N__12587),
            .I(N__12576));
    Odrv12 I__2931 (
            .O(N__12584),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__2930 (
            .O(N__12581),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2929 (
            .O(N__12576),
            .I(CONSTANT_ONE_NET));
    InMux I__2928 (
            .O(N__12569),
            .I(N__12566));
    LocalMux I__2927 (
            .O(N__12566),
            .I(N__12563));
    Span4Mux_h I__2926 (
            .O(N__12563),
            .I(N__12560));
    Odrv4 I__2925 (
            .O(N__12560),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_4 ));
    InMux I__2924 (
            .O(N__12557),
            .I(N__12554));
    LocalMux I__2923 (
            .O(N__12554),
            .I(N__12551));
    Span4Mux_h I__2922 (
            .O(N__12551),
            .I(N__12548));
    Odrv4 I__2921 (
            .O(N__12548),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_5 ));
    InMux I__2920 (
            .O(N__12545),
            .I(N__12542));
    LocalMux I__2919 (
            .O(N__12542),
            .I(N__12539));
    Span4Mux_h I__2918 (
            .O(N__12539),
            .I(N__12536));
    Odrv4 I__2917 (
            .O(N__12536),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_6 ));
    InMux I__2916 (
            .O(N__12533),
            .I(N__12530));
    LocalMux I__2915 (
            .O(N__12530),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_7 ));
    CEMux I__2914 (
            .O(N__12527),
            .I(N__12524));
    LocalMux I__2913 (
            .O(N__12524),
            .I(N__12520));
    InMux I__2912 (
            .O(N__12523),
            .I(N__12517));
    Span4Mux_v I__2911 (
            .O(N__12520),
            .I(N__12514));
    LocalMux I__2910 (
            .O(N__12517),
            .I(N__12511));
    Odrv4 I__2909 (
            .O(N__12514),
            .I(\DUT.fifo_tx_inst.rFifoData_awe3 ));
    Odrv12 I__2908 (
            .O(N__12511),
            .I(\DUT.fifo_tx_inst.rFifoData_awe3 ));
    InMux I__2907 (
            .O(N__12506),
            .I(N__12503));
    LocalMux I__2906 (
            .O(N__12503),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_1 ));
    InMux I__2905 (
            .O(N__12500),
            .I(N__12494));
    InMux I__2904 (
            .O(N__12499),
            .I(N__12491));
    InMux I__2903 (
            .O(N__12498),
            .I(N__12488));
    InMux I__2902 (
            .O(N__12497),
            .I(N__12485));
    LocalMux I__2901 (
            .O(N__12494),
            .I(N__12480));
    LocalMux I__2900 (
            .O(N__12491),
            .I(N__12480));
    LocalMux I__2899 (
            .O(N__12488),
            .I(N__12477));
    LocalMux I__2898 (
            .O(N__12485),
            .I(N__12474));
    Span4Mux_h I__2897 (
            .O(N__12480),
            .I(N__12471));
    Span4Mux_h I__2896 (
            .O(N__12477),
            .I(N__12466));
    Span4Mux_h I__2895 (
            .O(N__12474),
            .I(N__12466));
    Odrv4 I__2894 (
            .O(N__12471),
            .I(rTxByteZ0Z_2));
    Odrv4 I__2893 (
            .O(N__12466),
            .I(rTxByteZ0Z_2));
    CascadeMux I__2892 (
            .O(N__12461),
            .I(N__12458));
    InMux I__2891 (
            .O(N__12458),
            .I(N__12455));
    LocalMux I__2890 (
            .O(N__12455),
            .I(N__12452));
    Span4Mux_h I__2889 (
            .O(N__12452),
            .I(N__12449));
    Odrv4 I__2888 (
            .O(N__12449),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_2 ));
    InMux I__2887 (
            .O(N__12446),
            .I(N__12442));
    InMux I__2886 (
            .O(N__12445),
            .I(N__12439));
    LocalMux I__2885 (
            .O(N__12442),
            .I(N__12435));
    LocalMux I__2884 (
            .O(N__12439),
            .I(N__12432));
    InMux I__2883 (
            .O(N__12438),
            .I(N__12429));
    Span4Mux_h I__2882 (
            .O(N__12435),
            .I(N__12422));
    Span4Mux_v I__2881 (
            .O(N__12432),
            .I(N__12422));
    LocalMux I__2880 (
            .O(N__12429),
            .I(N__12422));
    Span4Mux_h I__2879 (
            .O(N__12422),
            .I(N__12418));
    InMux I__2878 (
            .O(N__12421),
            .I(N__12415));
    Odrv4 I__2877 (
            .O(N__12418),
            .I(rTxByteZ0Z_3));
    LocalMux I__2876 (
            .O(N__12415),
            .I(rTxByteZ0Z_3));
    InMux I__2875 (
            .O(N__12410),
            .I(N__12407));
    LocalMux I__2874 (
            .O(N__12407),
            .I(N__12404));
    Span4Mux_h I__2873 (
            .O(N__12404),
            .I(N__12401));
    Odrv4 I__2872 (
            .O(N__12401),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_3 ));
    InMux I__2871 (
            .O(N__12398),
            .I(N__12394));
    InMux I__2870 (
            .O(N__12397),
            .I(N__12391));
    LocalMux I__2869 (
            .O(N__12394),
            .I(N__12385));
    LocalMux I__2868 (
            .O(N__12391),
            .I(N__12385));
    InMux I__2867 (
            .O(N__12390),
            .I(N__12382));
    Span4Mux_v I__2866 (
            .O(N__12385),
            .I(N__12376));
    LocalMux I__2865 (
            .O(N__12382),
            .I(N__12376));
    InMux I__2864 (
            .O(N__12381),
            .I(N__12373));
    Odrv4 I__2863 (
            .O(N__12376),
            .I(rTxByteZ0Z_4));
    LocalMux I__2862 (
            .O(N__12373),
            .I(rTxByteZ0Z_4));
    CascadeMux I__2861 (
            .O(N__12368),
            .I(N__12365));
    InMux I__2860 (
            .O(N__12365),
            .I(N__12362));
    LocalMux I__2859 (
            .O(N__12362),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_4 ));
    CascadeMux I__2858 (
            .O(N__12359),
            .I(N__12356));
    InMux I__2857 (
            .O(N__12356),
            .I(N__12353));
    LocalMux I__2856 (
            .O(N__12353),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_6 ));
    InMux I__2855 (
            .O(N__12350),
            .I(N__12346));
    InMux I__2854 (
            .O(N__12349),
            .I(N__12343));
    LocalMux I__2853 (
            .O(N__12346),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_2 ));
    LocalMux I__2852 (
            .O(N__12343),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_2 ));
    InMux I__2851 (
            .O(N__12338),
            .I(N__12334));
    InMux I__2850 (
            .O(N__12337),
            .I(N__12331));
    LocalMux I__2849 (
            .O(N__12334),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_4 ));
    LocalMux I__2848 (
            .O(N__12331),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_4 ));
    CascadeMux I__2847 (
            .O(N__12326),
            .I(N__12322));
    InMux I__2846 (
            .O(N__12325),
            .I(N__12319));
    InMux I__2845 (
            .O(N__12322),
            .I(N__12316));
    LocalMux I__2844 (
            .O(N__12319),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_5 ));
    LocalMux I__2843 (
            .O(N__12316),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_5 ));
    InMux I__2842 (
            .O(N__12311),
            .I(N__12307));
    InMux I__2841 (
            .O(N__12310),
            .I(N__12304));
    LocalMux I__2840 (
            .O(N__12307),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_3 ));
    LocalMux I__2839 (
            .O(N__12304),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_3 ));
    InMux I__2838 (
            .O(N__12299),
            .I(N__12295));
    InMux I__2837 (
            .O(N__12298),
            .I(N__12292));
    LocalMux I__2836 (
            .O(N__12295),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_12 ));
    LocalMux I__2835 (
            .O(N__12292),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_12 ));
    InMux I__2834 (
            .O(N__12287),
            .I(N__12283));
    InMux I__2833 (
            .O(N__12286),
            .I(N__12280));
    LocalMux I__2832 (
            .O(N__12283),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_7 ));
    LocalMux I__2831 (
            .O(N__12280),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_7 ));
    CascadeMux I__2830 (
            .O(N__12275),
            .I(N__12271));
    InMux I__2829 (
            .O(N__12274),
            .I(N__12268));
    InMux I__2828 (
            .O(N__12271),
            .I(N__12265));
    LocalMux I__2827 (
            .O(N__12268),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_13 ));
    LocalMux I__2826 (
            .O(N__12265),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_13 ));
    InMux I__2825 (
            .O(N__12260),
            .I(N__12256));
    InMux I__2824 (
            .O(N__12259),
            .I(N__12253));
    LocalMux I__2823 (
            .O(N__12256),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_6 ));
    LocalMux I__2822 (
            .O(N__12253),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_6 ));
    InMux I__2821 (
            .O(N__12248),
            .I(N__12245));
    LocalMux I__2820 (
            .O(N__12245),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_9 ));
    InMux I__2819 (
            .O(N__12242),
            .I(N__12239));
    LocalMux I__2818 (
            .O(N__12239),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_7 ));
    CascadeMux I__2817 (
            .O(N__12236),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_8_cascade_ ));
    InMux I__2816 (
            .O(N__12233),
            .I(N__12230));
    LocalMux I__2815 (
            .O(N__12230),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_6 ));
    InMux I__2814 (
            .O(N__12227),
            .I(N__12218));
    InMux I__2813 (
            .O(N__12226),
            .I(N__12208));
    InMux I__2812 (
            .O(N__12225),
            .I(N__12208));
    InMux I__2811 (
            .O(N__12224),
            .I(N__12208));
    InMux I__2810 (
            .O(N__12223),
            .I(N__12205));
    InMux I__2809 (
            .O(N__12222),
            .I(N__12200));
    InMux I__2808 (
            .O(N__12221),
            .I(N__12200));
    LocalMux I__2807 (
            .O(N__12218),
            .I(N__12196));
    InMux I__2806 (
            .O(N__12217),
            .I(N__12189));
    InMux I__2805 (
            .O(N__12216),
            .I(N__12189));
    InMux I__2804 (
            .O(N__12215),
            .I(N__12189));
    LocalMux I__2803 (
            .O(N__12208),
            .I(N__12182));
    LocalMux I__2802 (
            .O(N__12205),
            .I(N__12182));
    LocalMux I__2801 (
            .O(N__12200),
            .I(N__12182));
    InMux I__2800 (
            .O(N__12199),
            .I(N__12179));
    Odrv4 I__2799 (
            .O(N__12196),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0 ));
    LocalMux I__2798 (
            .O(N__12189),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0 ));
    Odrv4 I__2797 (
            .O(N__12182),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0 ));
    LocalMux I__2796 (
            .O(N__12179),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0 ));
    InMux I__2795 (
            .O(N__12170),
            .I(N__12159));
    InMux I__2794 (
            .O(N__12169),
            .I(N__12159));
    InMux I__2793 (
            .O(N__12168),
            .I(N__12159));
    InMux I__2792 (
            .O(N__12167),
            .I(N__12148));
    InMux I__2791 (
            .O(N__12166),
            .I(N__12148));
    LocalMux I__2790 (
            .O(N__12159),
            .I(N__12145));
    InMux I__2789 (
            .O(N__12158),
            .I(N__12142));
    InMux I__2788 (
            .O(N__12157),
            .I(N__12137));
    InMux I__2787 (
            .O(N__12156),
            .I(N__12137));
    InMux I__2786 (
            .O(N__12155),
            .I(N__12130));
    InMux I__2785 (
            .O(N__12154),
            .I(N__12130));
    InMux I__2784 (
            .O(N__12153),
            .I(N__12130));
    LocalMux I__2783 (
            .O(N__12148),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_0 ));
    Odrv4 I__2782 (
            .O(N__12145),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_0 ));
    LocalMux I__2781 (
            .O(N__12142),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_0 ));
    LocalMux I__2780 (
            .O(N__12137),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_0 ));
    LocalMux I__2779 (
            .O(N__12130),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_0 ));
    CascadeMux I__2778 (
            .O(N__12119),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0_cascade_ ));
    InMux I__2777 (
            .O(N__12116),
            .I(N__12113));
    LocalMux I__2776 (
            .O(N__12113),
            .I(N__12110));
    Odrv12 I__2775 (
            .O(N__12110),
            .I(\DUT.uart_inst0.N_5_0 ));
    InMux I__2774 (
            .O(N__12107),
            .I(N__12104));
    LocalMux I__2773 (
            .O(N__12104),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_0 ));
    InMux I__2772 (
            .O(N__12101),
            .I(N__12098));
    LocalMux I__2771 (
            .O(N__12098),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_1 ));
    InMux I__2770 (
            .O(N__12095),
            .I(N__12092));
    LocalMux I__2769 (
            .O(N__12092),
            .I(N__12089));
    Odrv4 I__2768 (
            .O(N__12089),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_2 ));
    InMux I__2767 (
            .O(N__12086),
            .I(N__12083));
    LocalMux I__2766 (
            .O(N__12083),
            .I(N__12080));
    Odrv4 I__2765 (
            .O(N__12080),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_3 ));
    CascadeMux I__2764 (
            .O(N__12077),
            .I(\DUT.uart_inst0.g0_i_a3_0_cascade_ ));
    CascadeMux I__2763 (
            .O(N__12074),
            .I(N__12067));
    CascadeMux I__2762 (
            .O(N__12073),
            .I(N__12056));
    InMux I__2761 (
            .O(N__12072),
            .I(N__12053));
    InMux I__2760 (
            .O(N__12071),
            .I(N__12050));
    InMux I__2759 (
            .O(N__12070),
            .I(N__12047));
    InMux I__2758 (
            .O(N__12067),
            .I(N__12044));
    InMux I__2757 (
            .O(N__12066),
            .I(N__12041));
    InMux I__2756 (
            .O(N__12065),
            .I(N__12036));
    InMux I__2755 (
            .O(N__12064),
            .I(N__12036));
    InMux I__2754 (
            .O(N__12063),
            .I(N__12031));
    InMux I__2753 (
            .O(N__12062),
            .I(N__12031));
    InMux I__2752 (
            .O(N__12061),
            .I(N__12028));
    InMux I__2751 (
            .O(N__12060),
            .I(N__12025));
    InMux I__2750 (
            .O(N__12059),
            .I(N__12022));
    InMux I__2749 (
            .O(N__12056),
            .I(N__12019));
    LocalMux I__2748 (
            .O(N__12053),
            .I(N__12016));
    LocalMux I__2747 (
            .O(N__12050),
            .I(N__12013));
    LocalMux I__2746 (
            .O(N__12047),
            .I(N__12010));
    LocalMux I__2745 (
            .O(N__12044),
            .I(N__12007));
    LocalMux I__2744 (
            .O(N__12041),
            .I(N__12004));
    LocalMux I__2743 (
            .O(N__12036),
            .I(N__12001));
    LocalMux I__2742 (
            .O(N__12031),
            .I(N__11997));
    LocalMux I__2741 (
            .O(N__12028),
            .I(N__11994));
    LocalMux I__2740 (
            .O(N__12025),
            .I(N__11990));
    LocalMux I__2739 (
            .O(N__12022),
            .I(N__11986));
    LocalMux I__2738 (
            .O(N__12019),
            .I(N__11982));
    Glb2LocalMux I__2737 (
            .O(N__12016),
            .I(N__11930));
    Glb2LocalMux I__2736 (
            .O(N__12013),
            .I(N__11930));
    Glb2LocalMux I__2735 (
            .O(N__12010),
            .I(N__11930));
    Glb2LocalMux I__2734 (
            .O(N__12007),
            .I(N__11930));
    Glb2LocalMux I__2733 (
            .O(N__12004),
            .I(N__11930));
    Glb2LocalMux I__2732 (
            .O(N__12001),
            .I(N__11930));
    CEMux I__2731 (
            .O(N__12000),
            .I(N__11930));
    Glb2LocalMux I__2730 (
            .O(N__11997),
            .I(N__11930));
    Glb2LocalMux I__2729 (
            .O(N__11994),
            .I(N__11930));
    CEMux I__2728 (
            .O(N__11993),
            .I(N__11930));
    Glb2LocalMux I__2727 (
            .O(N__11990),
            .I(N__11930));
    CEMux I__2726 (
            .O(N__11989),
            .I(N__11930));
    Glb2LocalMux I__2725 (
            .O(N__11986),
            .I(N__11930));
    CEMux I__2724 (
            .O(N__11985),
            .I(N__11930));
    Glb2LocalMux I__2723 (
            .O(N__11982),
            .I(N__11930));
    CEMux I__2722 (
            .O(N__11981),
            .I(N__11930));
    CEMux I__2721 (
            .O(N__11980),
            .I(N__11930));
    CEMux I__2720 (
            .O(N__11979),
            .I(N__11930));
    CEMux I__2719 (
            .O(N__11978),
            .I(N__11930));
    CEMux I__2718 (
            .O(N__11977),
            .I(N__11930));
    CEMux I__2717 (
            .O(N__11976),
            .I(N__11930));
    CEMux I__2716 (
            .O(N__11975),
            .I(N__11930));
    GlobalMux I__2715 (
            .O(N__11930),
            .I(N__11927));
    gio2CtrlBuf I__2714 (
            .O(N__11927),
            .I(wPllLocked_g));
    InMux I__2713 (
            .O(N__11924),
            .I(N__11921));
    LocalMux I__2712 (
            .O(N__11921),
            .I(N__11915));
    CascadeMux I__2711 (
            .O(N__11920),
            .I(N__11912));
    InMux I__2710 (
            .O(N__11919),
            .I(N__11907));
    InMux I__2709 (
            .O(N__11918),
            .I(N__11904));
    Span4Mux_h I__2708 (
            .O(N__11915),
            .I(N__11901));
    InMux I__2707 (
            .O(N__11912),
            .I(N__11894));
    InMux I__2706 (
            .O(N__11911),
            .I(N__11894));
    InMux I__2705 (
            .O(N__11910),
            .I(N__11894));
    LocalMux I__2704 (
            .O(N__11907),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_4 ));
    LocalMux I__2703 (
            .O(N__11904),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_4 ));
    Odrv4 I__2702 (
            .O(N__11901),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_4 ));
    LocalMux I__2701 (
            .O(N__11894),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_4 ));
    InMux I__2700 (
            .O(N__11885),
            .I(N__11875));
    InMux I__2699 (
            .O(N__11884),
            .I(N__11872));
    CascadeMux I__2698 (
            .O(N__11883),
            .I(N__11869));
    InMux I__2697 (
            .O(N__11882),
            .I(N__11861));
    InMux I__2696 (
            .O(N__11881),
            .I(N__11861));
    InMux I__2695 (
            .O(N__11880),
            .I(N__11861));
    InMux I__2694 (
            .O(N__11879),
            .I(N__11856));
    InMux I__2693 (
            .O(N__11878),
            .I(N__11856));
    LocalMux I__2692 (
            .O(N__11875),
            .I(N__11853));
    LocalMux I__2691 (
            .O(N__11872),
            .I(N__11850));
    InMux I__2690 (
            .O(N__11869),
            .I(N__11845));
    InMux I__2689 (
            .O(N__11868),
            .I(N__11845));
    LocalMux I__2688 (
            .O(N__11861),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_3 ));
    LocalMux I__2687 (
            .O(N__11856),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_3 ));
    Odrv4 I__2686 (
            .O(N__11853),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_3 ));
    Odrv4 I__2685 (
            .O(N__11850),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_3 ));
    LocalMux I__2684 (
            .O(N__11845),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_3 ));
    InMux I__2683 (
            .O(N__11834),
            .I(N__11830));
    CascadeMux I__2682 (
            .O(N__11833),
            .I(N__11826));
    LocalMux I__2681 (
            .O(N__11830),
            .I(N__11823));
    CascadeMux I__2680 (
            .O(N__11829),
            .I(N__11818));
    InMux I__2679 (
            .O(N__11826),
            .I(N__11815));
    Span4Mux_h I__2678 (
            .O(N__11823),
            .I(N__11812));
    InMux I__2677 (
            .O(N__11822),
            .I(N__11809));
    InMux I__2676 (
            .O(N__11821),
            .I(N__11804));
    InMux I__2675 (
            .O(N__11818),
            .I(N__11804));
    LocalMux I__2674 (
            .O(N__11815),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_5 ));
    Odrv4 I__2673 (
            .O(N__11812),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_5 ));
    LocalMux I__2672 (
            .O(N__11809),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_5 ));
    LocalMux I__2671 (
            .O(N__11804),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_5 ));
    InMux I__2670 (
            .O(N__11795),
            .I(N__11792));
    LocalMux I__2669 (
            .O(N__11792),
            .I(\DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0 ));
    CascadeMux I__2668 (
            .O(N__11789),
            .I(\DUT.uart_inst0.g0_11_a3_2_cascade_ ));
    InMux I__2667 (
            .O(N__11786),
            .I(N__11783));
    LocalMux I__2666 (
            .O(N__11783),
            .I(N__11780));
    Odrv4 I__2665 (
            .O(N__11780),
            .I(\DUT.uart_inst0.N_7 ));
    InMux I__2664 (
            .O(N__11777),
            .I(N__11774));
    LocalMux I__2663 (
            .O(N__11774),
            .I(N__11769));
    InMux I__2662 (
            .O(N__11773),
            .I(N__11760));
    InMux I__2661 (
            .O(N__11772),
            .I(N__11757));
    Span4Mux_h I__2660 (
            .O(N__11769),
            .I(N__11754));
    InMux I__2659 (
            .O(N__11768),
            .I(N__11745));
    InMux I__2658 (
            .O(N__11767),
            .I(N__11745));
    InMux I__2657 (
            .O(N__11766),
            .I(N__11745));
    InMux I__2656 (
            .O(N__11765),
            .I(N__11745));
    InMux I__2655 (
            .O(N__11764),
            .I(N__11740));
    InMux I__2654 (
            .O(N__11763),
            .I(N__11740));
    LocalMux I__2653 (
            .O(N__11760),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_1 ));
    LocalMux I__2652 (
            .O(N__11757),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_1 ));
    Odrv4 I__2651 (
            .O(N__11754),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_1 ));
    LocalMux I__2650 (
            .O(N__11745),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_1 ));
    LocalMux I__2649 (
            .O(N__11740),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_1 ));
    CascadeMux I__2648 (
            .O(N__11729),
            .I(N__11725));
    CascadeMux I__2647 (
            .O(N__11728),
            .I(N__11720));
    InMux I__2646 (
            .O(N__11725),
            .I(N__11714));
    InMux I__2645 (
            .O(N__11724),
            .I(N__11705));
    InMux I__2644 (
            .O(N__11723),
            .I(N__11705));
    InMux I__2643 (
            .O(N__11720),
            .I(N__11705));
    InMux I__2642 (
            .O(N__11719),
            .I(N__11705));
    InMux I__2641 (
            .O(N__11718),
            .I(N__11700));
    InMux I__2640 (
            .O(N__11717),
            .I(N__11700));
    LocalMux I__2639 (
            .O(N__11714),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_2 ));
    LocalMux I__2638 (
            .O(N__11705),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_2 ));
    LocalMux I__2637 (
            .O(N__11700),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_2 ));
    InMux I__2636 (
            .O(N__11693),
            .I(N__11690));
    LocalMux I__2635 (
            .O(N__11690),
            .I(\DUT.uart_inst0.N_6_i ));
    InMux I__2634 (
            .O(N__11687),
            .I(N__11681));
    InMux I__2633 (
            .O(N__11686),
            .I(N__11677));
    InMux I__2632 (
            .O(N__11685),
            .I(N__11672));
    InMux I__2631 (
            .O(N__11684),
            .I(N__11672));
    LocalMux I__2630 (
            .O(N__11681),
            .I(N__11669));
    InMux I__2629 (
            .O(N__11680),
            .I(N__11666));
    LocalMux I__2628 (
            .O(N__11677),
            .I(N__11657));
    LocalMux I__2627 (
            .O(N__11672),
            .I(N__11652));
    Span4Mux_v I__2626 (
            .O(N__11669),
            .I(N__11652));
    LocalMux I__2625 (
            .O(N__11666),
            .I(N__11649));
    InMux I__2624 (
            .O(N__11665),
            .I(N__11638));
    InMux I__2623 (
            .O(N__11664),
            .I(N__11638));
    InMux I__2622 (
            .O(N__11663),
            .I(N__11638));
    InMux I__2621 (
            .O(N__11662),
            .I(N__11638));
    InMux I__2620 (
            .O(N__11661),
            .I(N__11638));
    InMux I__2619 (
            .O(N__11660),
            .I(N__11633));
    Span4Mux_h I__2618 (
            .O(N__11657),
            .I(N__11628));
    Span4Mux_v I__2617 (
            .O(N__11652),
            .I(N__11628));
    Span4Mux_v I__2616 (
            .O(N__11649),
            .I(N__11623));
    LocalMux I__2615 (
            .O(N__11638),
            .I(N__11623));
    InMux I__2614 (
            .O(N__11637),
            .I(N__11618));
    InMux I__2613 (
            .O(N__11636),
            .I(N__11618));
    LocalMux I__2612 (
            .O(N__11633),
            .I(\DUT.rTransmitZ0 ));
    Odrv4 I__2611 (
            .O(N__11628),
            .I(\DUT.rTransmitZ0 ));
    Odrv4 I__2610 (
            .O(N__11623),
            .I(\DUT.rTransmitZ0 ));
    LocalMux I__2609 (
            .O(N__11618),
            .I(\DUT.rTransmitZ0 ));
    InMux I__2608 (
            .O(N__11609),
            .I(N__11590));
    InMux I__2607 (
            .O(N__11608),
            .I(N__11585));
    InMux I__2606 (
            .O(N__11607),
            .I(N__11585));
    InMux I__2605 (
            .O(N__11606),
            .I(N__11582));
    InMux I__2604 (
            .O(N__11605),
            .I(N__11577));
    InMux I__2603 (
            .O(N__11604),
            .I(N__11577));
    CascadeMux I__2602 (
            .O(N__11603),
            .I(N__11573));
    CascadeMux I__2601 (
            .O(N__11602),
            .I(N__11570));
    CascadeMux I__2600 (
            .O(N__11601),
            .I(N__11567));
    CascadeMux I__2599 (
            .O(N__11600),
            .I(N__11561));
    CascadeMux I__2598 (
            .O(N__11599),
            .I(N__11558));
    CascadeMux I__2597 (
            .O(N__11598),
            .I(N__11555));
    CascadeMux I__2596 (
            .O(N__11597),
            .I(N__11552));
    CascadeMux I__2595 (
            .O(N__11596),
            .I(N__11549));
    CascadeMux I__2594 (
            .O(N__11595),
            .I(N__11542));
    CascadeMux I__2593 (
            .O(N__11594),
            .I(N__11538));
    CascadeMux I__2592 (
            .O(N__11593),
            .I(N__11533));
    LocalMux I__2591 (
            .O(N__11590),
            .I(N__11530));
    LocalMux I__2590 (
            .O(N__11585),
            .I(N__11527));
    LocalMux I__2589 (
            .O(N__11582),
            .I(N__11524));
    LocalMux I__2588 (
            .O(N__11577),
            .I(N__11521));
    InMux I__2587 (
            .O(N__11576),
            .I(N__11508));
    InMux I__2586 (
            .O(N__11573),
            .I(N__11508));
    InMux I__2585 (
            .O(N__11570),
            .I(N__11508));
    InMux I__2584 (
            .O(N__11567),
            .I(N__11508));
    InMux I__2583 (
            .O(N__11566),
            .I(N__11508));
    InMux I__2582 (
            .O(N__11565),
            .I(N__11508));
    InMux I__2581 (
            .O(N__11564),
            .I(N__11505));
    InMux I__2580 (
            .O(N__11561),
            .I(N__11500));
    InMux I__2579 (
            .O(N__11558),
            .I(N__11500));
    InMux I__2578 (
            .O(N__11555),
            .I(N__11483));
    InMux I__2577 (
            .O(N__11552),
            .I(N__11483));
    InMux I__2576 (
            .O(N__11549),
            .I(N__11483));
    InMux I__2575 (
            .O(N__11548),
            .I(N__11483));
    InMux I__2574 (
            .O(N__11547),
            .I(N__11483));
    InMux I__2573 (
            .O(N__11546),
            .I(N__11483));
    InMux I__2572 (
            .O(N__11545),
            .I(N__11483));
    InMux I__2571 (
            .O(N__11542),
            .I(N__11483));
    InMux I__2570 (
            .O(N__11541),
            .I(N__11480));
    InMux I__2569 (
            .O(N__11538),
            .I(N__11477));
    InMux I__2568 (
            .O(N__11537),
            .I(N__11472));
    InMux I__2567 (
            .O(N__11536),
            .I(N__11472));
    InMux I__2566 (
            .O(N__11533),
            .I(N__11469));
    Span4Mux_v I__2565 (
            .O(N__11530),
            .I(N__11462));
    Span4Mux_v I__2564 (
            .O(N__11527),
            .I(N__11462));
    Span4Mux_v I__2563 (
            .O(N__11524),
            .I(N__11462));
    Span4Mux_v I__2562 (
            .O(N__11521),
            .I(N__11457));
    LocalMux I__2561 (
            .O(N__11508),
            .I(N__11457));
    LocalMux I__2560 (
            .O(N__11505),
            .I(\DUT.tx_state_0 ));
    LocalMux I__2559 (
            .O(N__11500),
            .I(\DUT.tx_state_0 ));
    LocalMux I__2558 (
            .O(N__11483),
            .I(\DUT.tx_state_0 ));
    LocalMux I__2557 (
            .O(N__11480),
            .I(\DUT.tx_state_0 ));
    LocalMux I__2556 (
            .O(N__11477),
            .I(\DUT.tx_state_0 ));
    LocalMux I__2555 (
            .O(N__11472),
            .I(\DUT.tx_state_0 ));
    LocalMux I__2554 (
            .O(N__11469),
            .I(\DUT.tx_state_0 ));
    Odrv4 I__2553 (
            .O(N__11462),
            .I(\DUT.tx_state_0 ));
    Odrv4 I__2552 (
            .O(N__11457),
            .I(\DUT.tx_state_0 ));
    InMux I__2551 (
            .O(N__11438),
            .I(N__11434));
    InMux I__2550 (
            .O(N__11437),
            .I(N__11428));
    LocalMux I__2549 (
            .O(N__11434),
            .I(N__11425));
    InMux I__2548 (
            .O(N__11433),
            .I(N__11420));
    InMux I__2547 (
            .O(N__11432),
            .I(N__11420));
    InMux I__2546 (
            .O(N__11431),
            .I(N__11417));
    LocalMux I__2545 (
            .O(N__11428),
            .I(N__11403));
    Span4Mux_h I__2544 (
            .O(N__11425),
            .I(N__11398));
    LocalMux I__2543 (
            .O(N__11420),
            .I(N__11398));
    LocalMux I__2542 (
            .O(N__11417),
            .I(N__11395));
    InMux I__2541 (
            .O(N__11416),
            .I(N__11388));
    InMux I__2540 (
            .O(N__11415),
            .I(N__11388));
    InMux I__2539 (
            .O(N__11414),
            .I(N__11388));
    InMux I__2538 (
            .O(N__11413),
            .I(N__11377));
    InMux I__2537 (
            .O(N__11412),
            .I(N__11377));
    InMux I__2536 (
            .O(N__11411),
            .I(N__11377));
    InMux I__2535 (
            .O(N__11410),
            .I(N__11377));
    InMux I__2534 (
            .O(N__11409),
            .I(N__11377));
    InMux I__2533 (
            .O(N__11408),
            .I(N__11374));
    InMux I__2532 (
            .O(N__11407),
            .I(N__11371));
    InMux I__2531 (
            .O(N__11406),
            .I(N__11368));
    Span4Mux_v I__2530 (
            .O(N__11403),
            .I(N__11361));
    Span4Mux_v I__2529 (
            .O(N__11398),
            .I(N__11361));
    Span4Mux_v I__2528 (
            .O(N__11395),
            .I(N__11361));
    LocalMux I__2527 (
            .O(N__11388),
            .I(N__11358));
    LocalMux I__2526 (
            .O(N__11377),
            .I(N__11355));
    LocalMux I__2525 (
            .O(N__11374),
            .I(\DUT.uart_inst0.tx_stateZ0Z_1 ));
    LocalMux I__2524 (
            .O(N__11371),
            .I(\DUT.uart_inst0.tx_stateZ0Z_1 ));
    LocalMux I__2523 (
            .O(N__11368),
            .I(\DUT.uart_inst0.tx_stateZ0Z_1 ));
    Odrv4 I__2522 (
            .O(N__11361),
            .I(\DUT.uart_inst0.tx_stateZ0Z_1 ));
    Odrv4 I__2521 (
            .O(N__11358),
            .I(\DUT.uart_inst0.tx_stateZ0Z_1 ));
    Odrv4 I__2520 (
            .O(N__11355),
            .I(\DUT.uart_inst0.tx_stateZ0Z_1 ));
    InMux I__2519 (
            .O(N__11342),
            .I(N__11339));
    LocalMux I__2518 (
            .O(N__11339),
            .I(N__11336));
    Odrv4 I__2517 (
            .O(N__11336),
            .I(\DUT.uart_inst0.N_11_1 ));
    CascadeMux I__2516 (
            .O(N__11333),
            .I(N__11330));
    InMux I__2515 (
            .O(N__11330),
            .I(N__11326));
    InMux I__2514 (
            .O(N__11329),
            .I(N__11323));
    LocalMux I__2513 (
            .O(N__11326),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_9 ));
    LocalMux I__2512 (
            .O(N__11323),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_9 ));
    InMux I__2511 (
            .O(N__11318),
            .I(N__11314));
    InMux I__2510 (
            .O(N__11317),
            .I(N__11311));
    LocalMux I__2509 (
            .O(N__11314),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_10 ));
    LocalMux I__2508 (
            .O(N__11311),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_10 ));
    CascadeMux I__2507 (
            .O(N__11306),
            .I(N__11302));
    CascadeMux I__2506 (
            .O(N__11305),
            .I(N__11299));
    InMux I__2505 (
            .O(N__11302),
            .I(N__11296));
    InMux I__2504 (
            .O(N__11299),
            .I(N__11293));
    LocalMux I__2503 (
            .O(N__11296),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_11 ));
    LocalMux I__2502 (
            .O(N__11293),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_11 ));
    InMux I__2501 (
            .O(N__11288),
            .I(N__11284));
    InMux I__2500 (
            .O(N__11287),
            .I(N__11281));
    LocalMux I__2499 (
            .O(N__11284),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_8 ));
    LocalMux I__2498 (
            .O(N__11281),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_8 ));
    SRMux I__2497 (
            .O(N__11276),
            .I(N__11273));
    LocalMux I__2496 (
            .O(N__11273),
            .I(N__11269));
    SRMux I__2495 (
            .O(N__11272),
            .I(N__11265));
    Span4Mux_h I__2494 (
            .O(N__11269),
            .I(N__11262));
    SRMux I__2493 (
            .O(N__11268),
            .I(N__11259));
    LocalMux I__2492 (
            .O(N__11265),
            .I(\DUT.uart_inst0.N_20 ));
    Odrv4 I__2491 (
            .O(N__11262),
            .I(\DUT.uart_inst0.N_20 ));
    LocalMux I__2490 (
            .O(N__11259),
            .I(\DUT.uart_inst0.N_20 ));
    InMux I__2489 (
            .O(N__11252),
            .I(N__11248));
    InMux I__2488 (
            .O(N__11251),
            .I(N__11245));
    LocalMux I__2487 (
            .O(N__11248),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_1 ));
    LocalMux I__2486 (
            .O(N__11245),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_1 ));
    InMux I__2485 (
            .O(N__11240),
            .I(N__11235));
    InMux I__2484 (
            .O(N__11239),
            .I(N__11230));
    InMux I__2483 (
            .O(N__11238),
            .I(N__11230));
    LocalMux I__2482 (
            .O(N__11235),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_0 ));
    LocalMux I__2481 (
            .O(N__11230),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_0 ));
    CascadeMux I__2480 (
            .O(N__11225),
            .I(\DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0_cascade_ ));
    InMux I__2479 (
            .O(N__11222),
            .I(N__11218));
    InMux I__2478 (
            .O(N__11221),
            .I(N__11215));
    LocalMux I__2477 (
            .O(N__11218),
            .I(\DUT.uart_inst0.N_77 ));
    LocalMux I__2476 (
            .O(N__11215),
            .I(\DUT.uart_inst0.N_77 ));
    InMux I__2475 (
            .O(N__11210),
            .I(N__11207));
    LocalMux I__2474 (
            .O(N__11207),
            .I(\DUT.uart_inst0.g0_i_o2_2 ));
    InMux I__2473 (
            .O(N__11204),
            .I(N__11201));
    LocalMux I__2472 (
            .O(N__11201),
            .I(\DUT.uart_inst0.g0_i_o2_3 ));
    CascadeMux I__2471 (
            .O(N__11198),
            .I(N__11195));
    InMux I__2470 (
            .O(N__11195),
            .I(N__11192));
    LocalMux I__2469 (
            .O(N__11192),
            .I(N__11189));
    Span4Mux_h I__2468 (
            .O(N__11189),
            .I(N__11186));
    Odrv4 I__2467 (
            .O(N__11186),
            .I(\DUT.uart_inst0.N_11 ));
    InMux I__2466 (
            .O(N__11183),
            .I(N__11180));
    LocalMux I__2465 (
            .O(N__11180),
            .I(N__11177));
    Span4Mux_h I__2464 (
            .O(N__11177),
            .I(N__11174));
    Odrv4 I__2463 (
            .O(N__11174),
            .I(\DUT.uart_inst0.g0_11_a4_2 ));
    CascadeMux I__2462 (
            .O(N__11171),
            .I(N__11168));
    InMux I__2461 (
            .O(N__11168),
            .I(N__11165));
    LocalMux I__2460 (
            .O(N__11165),
            .I(N__11162));
    Span4Mux_v I__2459 (
            .O(N__11162),
            .I(N__11159));
    Span4Mux_h I__2458 (
            .O(N__11159),
            .I(N__11156));
    Odrv4 I__2457 (
            .O(N__11156),
            .I(\DUT.uart_inst0.N_9 ));
    CascadeMux I__2456 (
            .O(N__11153),
            .I(\DUT.uart_inst0.tx_state_ns_i_i_o2_a0_2_0_cascade_ ));
    InMux I__2455 (
            .O(N__11150),
            .I(N__11146));
    InMux I__2454 (
            .O(N__11149),
            .I(N__11143));
    LocalMux I__2453 (
            .O(N__11146),
            .I(\DUT.uart_inst0.N_71_i ));
    LocalMux I__2452 (
            .O(N__11143),
            .I(\DUT.uart_inst0.N_71_i ));
    CascadeMux I__2451 (
            .O(N__11138),
            .I(N__11135));
    InMux I__2450 (
            .O(N__11135),
            .I(N__11132));
    LocalMux I__2449 (
            .O(N__11132),
            .I(N__11129));
    Span4Mux_h I__2448 (
            .O(N__11129),
            .I(N__11126));
    Odrv4 I__2447 (
            .O(N__11126),
            .I(\DUT.uart_inst0.N_8_1 ));
    InMux I__2446 (
            .O(N__11123),
            .I(N__11117));
    InMux I__2445 (
            .O(N__11122),
            .I(N__11112));
    InMux I__2444 (
            .O(N__11121),
            .I(N__11112));
    InMux I__2443 (
            .O(N__11120),
            .I(N__11109));
    LocalMux I__2442 (
            .O(N__11117),
            .I(N__11105));
    LocalMux I__2441 (
            .O(N__11112),
            .I(N__11100));
    LocalMux I__2440 (
            .O(N__11109),
            .I(N__11100));
    InMux I__2439 (
            .O(N__11108),
            .I(N__11097));
    Span4Mux_v I__2438 (
            .O(N__11105),
            .I(N__11094));
    Span4Mux_v I__2437 (
            .O(N__11100),
            .I(N__11089));
    LocalMux I__2436 (
            .O(N__11097),
            .I(N__11089));
    Sp12to4 I__2435 (
            .O(N__11094),
            .I(N__11086));
    Span4Mux_v I__2434 (
            .O(N__11089),
            .I(N__11083));
    Span12Mux_h I__2433 (
            .O(N__11086),
            .I(N__11080));
    Sp12to4 I__2432 (
            .O(N__11083),
            .I(N__11077));
    Span12Mux_v I__2431 (
            .O(N__11080),
            .I(N__11074));
    Span12Mux_h I__2430 (
            .O(N__11077),
            .I(N__11071));
    Odrv12 I__2429 (
            .O(N__11074),
            .I(iRxF_n_c));
    Odrv12 I__2428 (
            .O(N__11071),
            .I(iRxF_n_c));
    InMux I__2427 (
            .O(N__11066),
            .I(N__11062));
    InMux I__2426 (
            .O(N__11065),
            .I(N__11058));
    LocalMux I__2425 (
            .O(N__11062),
            .I(N__11055));
    InMux I__2424 (
            .O(N__11061),
            .I(N__11052));
    LocalMux I__2423 (
            .O(N__11058),
            .I(N__11049));
    Span4Mux_v I__2422 (
            .O(N__11055),
            .I(N__11044));
    LocalMux I__2421 (
            .O(N__11052),
            .I(N__11044));
    Span4Mux_v I__2420 (
            .O(N__11049),
            .I(N__11041));
    Span4Mux_v I__2419 (
            .O(N__11044),
            .I(N__11038));
    Sp12to4 I__2418 (
            .O(N__11041),
            .I(N__11035));
    Sp12to4 I__2417 (
            .O(N__11038),
            .I(N__11032));
    Span12Mux_h I__2416 (
            .O(N__11035),
            .I(N__11029));
    Span12Mux_h I__2415 (
            .O(N__11032),
            .I(N__11026));
    Span12Mux_v I__2414 (
            .O(N__11029),
            .I(N__11023));
    Span12Mux_v I__2413 (
            .O(N__11026),
            .I(N__11020));
    Odrv12 I__2412 (
            .O(N__11023),
            .I(iTxE_n_c));
    Odrv12 I__2411 (
            .O(N__11020),
            .I(iTxE_n_c));
    InMux I__2410 (
            .O(N__11015),
            .I(N__11012));
    LocalMux I__2409 (
            .O(N__11012),
            .I(N__11006));
    InMux I__2408 (
            .O(N__11011),
            .I(N__11000));
    InMux I__2407 (
            .O(N__11010),
            .I(N__11000));
    InMux I__2406 (
            .O(N__11009),
            .I(N__10997));
    Span4Mux_v I__2405 (
            .O(N__11006),
            .I(N__10994));
    InMux I__2404 (
            .O(N__11005),
            .I(N__10991));
    LocalMux I__2403 (
            .O(N__11000),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_0 ));
    LocalMux I__2402 (
            .O(N__10997),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_0 ));
    Odrv4 I__2401 (
            .O(N__10994),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_0 ));
    LocalMux I__2400 (
            .O(N__10991),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_0 ));
    InMux I__2399 (
            .O(N__10982),
            .I(N__10979));
    LocalMux I__2398 (
            .O(N__10979),
            .I(\fifo_inst.ft2232h_inst.N_101 ));
    CascadeMux I__2397 (
            .O(N__10976),
            .I(\DUT.uart_inst0.N_13_cascade_ ));
    CascadeMux I__2396 (
            .O(N__10973),
            .I(\DUT.uart_inst0.g0_i_0_cascade_ ));
    InMux I__2395 (
            .O(N__10970),
            .I(N__10967));
    LocalMux I__2394 (
            .O(N__10967),
            .I(N__10964));
    Odrv4 I__2393 (
            .O(N__10964),
            .I(\DUT.uart_inst0.g0_i_a6_0 ));
    CascadeMux I__2392 (
            .O(N__10961),
            .I(\DUT.uart_inst0.g0_i_1_cascade_ ));
    InMux I__2391 (
            .O(N__10958),
            .I(N__10955));
    LocalMux I__2390 (
            .O(N__10955),
            .I(\DUT.uart_inst0.g0_i_a6_3_0 ));
    CascadeMux I__2389 (
            .O(N__10952),
            .I(\DUT.uart_inst0.g0_i_o2_1_cascade_ ));
    InMux I__2388 (
            .O(N__10949),
            .I(N__10946));
    LocalMux I__2387 (
            .O(N__10946),
            .I(N__10943));
    Span4Mux_v I__2386 (
            .O(N__10943),
            .I(N__10940));
    Odrv4 I__2385 (
            .O(N__10940),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_5 ));
    CascadeMux I__2384 (
            .O(N__10937),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ));
    InMux I__2383 (
            .O(N__10934),
            .I(N__10931));
    LocalMux I__2382 (
            .O(N__10931),
            .I(N__10928));
    Span4Mux_h I__2381 (
            .O(N__10928),
            .I(N__10925));
    Odrv4 I__2380 (
            .O(N__10925),
            .I(\DUT.rFifoDatarx_5 ));
    InMux I__2379 (
            .O(N__10922),
            .I(N__10919));
    LocalMux I__2378 (
            .O(N__10919),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_5 ));
    CascadeMux I__2377 (
            .O(N__10916),
            .I(N__10911));
    InMux I__2376 (
            .O(N__10915),
            .I(N__10896));
    InMux I__2375 (
            .O(N__10914),
            .I(N__10896));
    InMux I__2374 (
            .O(N__10911),
            .I(N__10893));
    InMux I__2373 (
            .O(N__10910),
            .I(N__10886));
    InMux I__2372 (
            .O(N__10909),
            .I(N__10886));
    InMux I__2371 (
            .O(N__10908),
            .I(N__10886));
    InMux I__2370 (
            .O(N__10907),
            .I(N__10879));
    InMux I__2369 (
            .O(N__10906),
            .I(N__10879));
    InMux I__2368 (
            .O(N__10905),
            .I(N__10879));
    InMux I__2367 (
            .O(N__10904),
            .I(N__10872));
    InMux I__2366 (
            .O(N__10903),
            .I(N__10872));
    InMux I__2365 (
            .O(N__10902),
            .I(N__10872));
    InMux I__2364 (
            .O(N__10901),
            .I(N__10869));
    LocalMux I__2363 (
            .O(N__10896),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__2362 (
            .O(N__10893),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__2361 (
            .O(N__10886),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__2360 (
            .O(N__10879),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__2359 (
            .O(N__10872),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__2358 (
            .O(N__10869),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    CascadeMux I__2357 (
            .O(N__10856),
            .I(N__10843));
    CascadeMux I__2356 (
            .O(N__10855),
            .I(N__10836));
    CascadeMux I__2355 (
            .O(N__10854),
            .I(N__10833));
    CascadeMux I__2354 (
            .O(N__10853),
            .I(N__10827));
    CascadeMux I__2353 (
            .O(N__10852),
            .I(N__10822));
    InMux I__2352 (
            .O(N__10851),
            .I(N__10819));
    InMux I__2351 (
            .O(N__10850),
            .I(N__10816));
    InMux I__2350 (
            .O(N__10849),
            .I(N__10803));
    InMux I__2349 (
            .O(N__10848),
            .I(N__10803));
    InMux I__2348 (
            .O(N__10847),
            .I(N__10803));
    InMux I__2347 (
            .O(N__10846),
            .I(N__10803));
    InMux I__2346 (
            .O(N__10843),
            .I(N__10803));
    InMux I__2345 (
            .O(N__10842),
            .I(N__10803));
    InMux I__2344 (
            .O(N__10841),
            .I(N__10790));
    InMux I__2343 (
            .O(N__10840),
            .I(N__10790));
    InMux I__2342 (
            .O(N__10839),
            .I(N__10790));
    InMux I__2341 (
            .O(N__10836),
            .I(N__10790));
    InMux I__2340 (
            .O(N__10833),
            .I(N__10790));
    InMux I__2339 (
            .O(N__10832),
            .I(N__10790));
    InMux I__2338 (
            .O(N__10831),
            .I(N__10779));
    InMux I__2337 (
            .O(N__10830),
            .I(N__10779));
    InMux I__2336 (
            .O(N__10827),
            .I(N__10779));
    InMux I__2335 (
            .O(N__10826),
            .I(N__10779));
    InMux I__2334 (
            .O(N__10825),
            .I(N__10779));
    InMux I__2333 (
            .O(N__10822),
            .I(N__10776));
    LocalMux I__2332 (
            .O(N__10819),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__2331 (
            .O(N__10816),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__2330 (
            .O(N__10803),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__2329 (
            .O(N__10790),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__2328 (
            .O(N__10779),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__2327 (
            .O(N__10776),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    CascadeMux I__2326 (
            .O(N__10763),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_ ));
    InMux I__2325 (
            .O(N__10760),
            .I(N__10757));
    LocalMux I__2324 (
            .O(N__10757),
            .I(N__10754));
    Span4Mux_h I__2323 (
            .O(N__10754),
            .I(N__10751));
    Odrv4 I__2322 (
            .O(N__10751),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_6 ));
    InMux I__2321 (
            .O(N__10748),
            .I(N__10745));
    LocalMux I__2320 (
            .O(N__10745),
            .I(N__10742));
    Span4Mux_v I__2319 (
            .O(N__10742),
            .I(N__10739));
    Odrv4 I__2318 (
            .O(N__10739),
            .I(\DUT.rFifoDatarx_6 ));
    CascadeMux I__2317 (
            .O(N__10736),
            .I(N__10731));
    CascadeMux I__2316 (
            .O(N__10735),
            .I(N__10726));
    CascadeMux I__2315 (
            .O(N__10734),
            .I(N__10723));
    InMux I__2314 (
            .O(N__10731),
            .I(N__10718));
    InMux I__2313 (
            .O(N__10730),
            .I(N__10718));
    InMux I__2312 (
            .O(N__10729),
            .I(N__10715));
    InMux I__2311 (
            .O(N__10726),
            .I(N__10710));
    InMux I__2310 (
            .O(N__10723),
            .I(N__10710));
    LocalMux I__2309 (
            .O(N__10718),
            .I(\DUT.rFifoCount_0 ));
    LocalMux I__2308 (
            .O(N__10715),
            .I(\DUT.rFifoCount_0 ));
    LocalMux I__2307 (
            .O(N__10710),
            .I(\DUT.rFifoCount_0 ));
    CascadeMux I__2306 (
            .O(N__10703),
            .I(N__10700));
    InMux I__2305 (
            .O(N__10700),
            .I(N__10697));
    LocalMux I__2304 (
            .O(N__10697),
            .I(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0 ));
    CascadeMux I__2303 (
            .O(N__10694),
            .I(N__10691));
    InMux I__2302 (
            .O(N__10691),
            .I(N__10688));
    LocalMux I__2301 (
            .O(N__10688),
            .I(\DUT.fifo_tx_inst.rFifoCount_RNIBPFMZ0Z_1 ));
    InMux I__2300 (
            .O(N__10685),
            .I(N__10679));
    InMux I__2299 (
            .O(N__10684),
            .I(N__10672));
    InMux I__2298 (
            .O(N__10683),
            .I(N__10672));
    InMux I__2297 (
            .O(N__10682),
            .I(N__10672));
    LocalMux I__2296 (
            .O(N__10679),
            .I(\DUT.rFifoCount_1 ));
    LocalMux I__2295 (
            .O(N__10672),
            .I(\DUT.rFifoCount_1 ));
    InMux I__2294 (
            .O(N__10667),
            .I(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0 ));
    InMux I__2293 (
            .O(N__10664),
            .I(N__10660));
    InMux I__2292 (
            .O(N__10663),
            .I(N__10649));
    LocalMux I__2291 (
            .O(N__10660),
            .I(N__10644));
    InMux I__2290 (
            .O(N__10659),
            .I(N__10633));
    InMux I__2289 (
            .O(N__10658),
            .I(N__10633));
    InMux I__2288 (
            .O(N__10657),
            .I(N__10633));
    InMux I__2287 (
            .O(N__10656),
            .I(N__10633));
    InMux I__2286 (
            .O(N__10655),
            .I(N__10633));
    InMux I__2285 (
            .O(N__10654),
            .I(N__10630));
    InMux I__2284 (
            .O(N__10653),
            .I(N__10627));
    InMux I__2283 (
            .O(N__10652),
            .I(N__10624));
    LocalMux I__2282 (
            .O(N__10649),
            .I(N__10621));
    InMux I__2281 (
            .O(N__10648),
            .I(N__10616));
    InMux I__2280 (
            .O(N__10647),
            .I(N__10616));
    Span4Mux_h I__2279 (
            .O(N__10644),
            .I(N__10611));
    LocalMux I__2278 (
            .O(N__10633),
            .I(N__10611));
    LocalMux I__2277 (
            .O(N__10630),
            .I(rRxReadZ0));
    LocalMux I__2276 (
            .O(N__10627),
            .I(rRxReadZ0));
    LocalMux I__2275 (
            .O(N__10624),
            .I(rRxReadZ0));
    Odrv4 I__2274 (
            .O(N__10621),
            .I(rRxReadZ0));
    LocalMux I__2273 (
            .O(N__10616),
            .I(rRxReadZ0));
    Odrv4 I__2272 (
            .O(N__10611),
            .I(rRxReadZ0));
    InMux I__2271 (
            .O(N__10598),
            .I(N__10589));
    InMux I__2270 (
            .O(N__10597),
            .I(N__10589));
    InMux I__2269 (
            .O(N__10596),
            .I(N__10586));
    InMux I__2268 (
            .O(N__10595),
            .I(N__10581));
    InMux I__2267 (
            .O(N__10594),
            .I(N__10581));
    LocalMux I__2266 (
            .O(N__10589),
            .I(\DUT.fifo_tx_inst.N_83 ));
    LocalMux I__2265 (
            .O(N__10586),
            .I(\DUT.fifo_tx_inst.N_83 ));
    LocalMux I__2264 (
            .O(N__10581),
            .I(\DUT.fifo_tx_inst.N_83 ));
    InMux I__2263 (
            .O(N__10574),
            .I(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1 ));
    InMux I__2262 (
            .O(N__10571),
            .I(N__10568));
    LocalMux I__2261 (
            .O(N__10568),
            .I(N__10564));
    CascadeMux I__2260 (
            .O(N__10567),
            .I(N__10561));
    Span4Mux_h I__2259 (
            .O(N__10564),
            .I(N__10558));
    InMux I__2258 (
            .O(N__10561),
            .I(N__10550));
    Span4Mux_v I__2257 (
            .O(N__10558),
            .I(N__10547));
    InMux I__2256 (
            .O(N__10557),
            .I(N__10536));
    InMux I__2255 (
            .O(N__10556),
            .I(N__10536));
    InMux I__2254 (
            .O(N__10555),
            .I(N__10536));
    InMux I__2253 (
            .O(N__10554),
            .I(N__10536));
    InMux I__2252 (
            .O(N__10553),
            .I(N__10536));
    LocalMux I__2251 (
            .O(N__10550),
            .I(\DUT.rFifoCount_2 ));
    Odrv4 I__2250 (
            .O(N__10547),
            .I(\DUT.rFifoCount_2 ));
    LocalMux I__2249 (
            .O(N__10536),
            .I(\DUT.rFifoCount_2 ));
    SRMux I__2248 (
            .O(N__10529),
            .I(N__10502));
    SRMux I__2247 (
            .O(N__10528),
            .I(N__10502));
    SRMux I__2246 (
            .O(N__10527),
            .I(N__10502));
    SRMux I__2245 (
            .O(N__10526),
            .I(N__10502));
    SRMux I__2244 (
            .O(N__10525),
            .I(N__10502));
    SRMux I__2243 (
            .O(N__10524),
            .I(N__10502));
    SRMux I__2242 (
            .O(N__10523),
            .I(N__10502));
    SRMux I__2241 (
            .O(N__10522),
            .I(N__10502));
    SRMux I__2240 (
            .O(N__10521),
            .I(N__10502));
    GlobalMux I__2239 (
            .O(N__10502),
            .I(N__10499));
    gio2CtrlBuf I__2238 (
            .O(N__10499),
            .I(wPllLocked_i_g));
    InMux I__2237 (
            .O(N__10496),
            .I(N__10493));
    LocalMux I__2236 (
            .O(N__10493),
            .I(N__10487));
    InMux I__2235 (
            .O(N__10492),
            .I(N__10484));
    InMux I__2234 (
            .O(N__10491),
            .I(N__10481));
    InMux I__2233 (
            .O(N__10490),
            .I(N__10478));
    Span4Mux_h I__2232 (
            .O(N__10487),
            .I(N__10473));
    LocalMux I__2231 (
            .O(N__10484),
            .I(N__10473));
    LocalMux I__2230 (
            .O(N__10481),
            .I(N__10470));
    LocalMux I__2229 (
            .O(N__10478),
            .I(N__10466));
    Span4Mux_v I__2228 (
            .O(N__10473),
            .I(N__10461));
    Span4Mux_h I__2227 (
            .O(N__10470),
            .I(N__10461));
    InMux I__2226 (
            .O(N__10469),
            .I(N__10458));
    Odrv12 I__2225 (
            .O(N__10466),
            .I(\DUT.wRxByte_7 ));
    Odrv4 I__2224 (
            .O(N__10461),
            .I(\DUT.wRxByte_7 ));
    LocalMux I__2223 (
            .O(N__10458),
            .I(\DUT.wRxByte_7 ));
    InMux I__2222 (
            .O(N__10451),
            .I(N__10448));
    LocalMux I__2221 (
            .O(N__10448),
            .I(N__10445));
    Odrv4 I__2220 (
            .O(N__10445),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_7 ));
    CEMux I__2219 (
            .O(N__10442),
            .I(N__10438));
    CEMux I__2218 (
            .O(N__10441),
            .I(N__10434));
    LocalMux I__2217 (
            .O(N__10438),
            .I(N__10431));
    CEMux I__2216 (
            .O(N__10437),
            .I(N__10428));
    LocalMux I__2215 (
            .O(N__10434),
            .I(N__10425));
    Span4Mux_v I__2214 (
            .O(N__10431),
            .I(N__10421));
    LocalMux I__2213 (
            .O(N__10428),
            .I(N__10418));
    Span4Mux_h I__2212 (
            .O(N__10425),
            .I(N__10415));
    InMux I__2211 (
            .O(N__10424),
            .I(N__10412));
    Odrv4 I__2210 (
            .O(N__10421),
            .I(\DUT.fifo_rx_inst.rFifoData_awe0 ));
    Odrv4 I__2209 (
            .O(N__10418),
            .I(\DUT.fifo_rx_inst.rFifoData_awe0 ));
    Odrv4 I__2208 (
            .O(N__10415),
            .I(\DUT.fifo_rx_inst.rFifoData_awe0 ));
    LocalMux I__2207 (
            .O(N__10412),
            .I(\DUT.fifo_rx_inst.rFifoData_awe0 ));
    CascadeMux I__2206 (
            .O(N__10403),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ));
    InMux I__2205 (
            .O(N__10400),
            .I(N__10397));
    LocalMux I__2204 (
            .O(N__10397),
            .I(N__10394));
    Span4Mux_h I__2203 (
            .O(N__10394),
            .I(N__10391));
    Odrv4 I__2202 (
            .O(N__10391),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_0 ));
    InMux I__2201 (
            .O(N__10388),
            .I(N__10385));
    LocalMux I__2200 (
            .O(N__10385),
            .I(N__10382));
    Span4Mux_v I__2199 (
            .O(N__10382),
            .I(N__10379));
    Odrv4 I__2198 (
            .O(N__10379),
            .I(\DUT.rFifoDatarxZ0Z_0 ));
    InMux I__2197 (
            .O(N__10376),
            .I(N__10373));
    LocalMux I__2196 (
            .O(N__10373),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_0 ));
    InMux I__2195 (
            .O(N__10370),
            .I(N__10367));
    LocalMux I__2194 (
            .O(N__10367),
            .I(N__10364));
    Span4Mux_h I__2193 (
            .O(N__10364),
            .I(N__10361));
    Odrv4 I__2192 (
            .O(N__10361),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_1 ));
    CascadeMux I__2191 (
            .O(N__10358),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1_cascade_ ));
    InMux I__2190 (
            .O(N__10355),
            .I(N__10352));
    LocalMux I__2189 (
            .O(N__10352),
            .I(N__10349));
    Span4Mux_v I__2188 (
            .O(N__10349),
            .I(N__10346));
    Odrv4 I__2187 (
            .O(N__10346),
            .I(\DUT.rFifoDatarx_1 ));
    CascadeMux I__2186 (
            .O(N__10343),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_ ));
    InMux I__2185 (
            .O(N__10340),
            .I(N__10337));
    LocalMux I__2184 (
            .O(N__10337),
            .I(N__10334));
    Span4Mux_v I__2183 (
            .O(N__10334),
            .I(N__10331));
    Odrv4 I__2182 (
            .O(N__10331),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_4 ));
    InMux I__2181 (
            .O(N__10328),
            .I(N__10325));
    LocalMux I__2180 (
            .O(N__10325),
            .I(N__10322));
    Span4Mux_h I__2179 (
            .O(N__10322),
            .I(N__10319));
    Odrv4 I__2178 (
            .O(N__10319),
            .I(\DUT.rFifoDatarx_4 ));
    InMux I__2177 (
            .O(N__10316),
            .I(N__10313));
    LocalMux I__2176 (
            .O(N__10313),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_4 ));
    InMux I__2175 (
            .O(N__10310),
            .I(bfn_11_19_0_));
    InMux I__2174 (
            .O(N__10307),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_8 ));
    InMux I__2173 (
            .O(N__10304),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_9 ));
    InMux I__2172 (
            .O(N__10301),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_10 ));
    InMux I__2171 (
            .O(N__10298),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_11 ));
    InMux I__2170 (
            .O(N__10295),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_12 ));
    InMux I__2169 (
            .O(N__10292),
            .I(N__10289));
    LocalMux I__2168 (
            .O(N__10289),
            .I(N__10286));
    Odrv12 I__2167 (
            .O(N__10286),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_7 ));
    CascadeMux I__2166 (
            .O(N__10283),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_ ));
    InMux I__2165 (
            .O(N__10280),
            .I(N__10277));
    LocalMux I__2164 (
            .O(N__10277),
            .I(N__10274));
    Odrv4 I__2163 (
            .O(N__10274),
            .I(\DUT.rFifoDatarx_7 ));
    InMux I__2162 (
            .O(N__10271),
            .I(N__10268));
    LocalMux I__2161 (
            .O(N__10268),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_7 ));
    SRMux I__2160 (
            .O(N__10265),
            .I(N__10262));
    LocalMux I__2159 (
            .O(N__10262),
            .I(N__10259));
    Span4Mux_h I__2158 (
            .O(N__10259),
            .I(N__10256));
    Span4Mux_h I__2157 (
            .O(N__10256),
            .I(N__10253));
    Odrv4 I__2156 (
            .O(N__10253),
            .I(\DUT.uart_inst0.N_65_i ));
    CascadeMux I__2155 (
            .O(N__10250),
            .I(N__10247));
    InMux I__2154 (
            .O(N__10247),
            .I(N__10243));
    InMux I__2153 (
            .O(N__10246),
            .I(N__10240));
    LocalMux I__2152 (
            .O(N__10243),
            .I(\DUT.uart_inst0.tx_dataZ0Z_0 ));
    LocalMux I__2151 (
            .O(N__10240),
            .I(\DUT.uart_inst0.tx_dataZ0Z_0 ));
    InMux I__2150 (
            .O(N__10235),
            .I(N__10229));
    InMux I__2149 (
            .O(N__10234),
            .I(N__10226));
    InMux I__2148 (
            .O(N__10233),
            .I(N__10223));
    InMux I__2147 (
            .O(N__10232),
            .I(N__10220));
    LocalMux I__2146 (
            .O(N__10229),
            .I(\DUT.uart_inst0.N_85 ));
    LocalMux I__2145 (
            .O(N__10226),
            .I(\DUT.uart_inst0.N_85 ));
    LocalMux I__2144 (
            .O(N__10223),
            .I(\DUT.uart_inst0.N_85 ));
    LocalMux I__2143 (
            .O(N__10220),
            .I(\DUT.uart_inst0.N_85 ));
    InMux I__2142 (
            .O(N__10211),
            .I(N__10208));
    LocalMux I__2141 (
            .O(N__10208),
            .I(\DUT.uart_inst0.N_89 ));
    InMux I__2140 (
            .O(N__10205),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_0 ));
    InMux I__2139 (
            .O(N__10202),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_1 ));
    InMux I__2138 (
            .O(N__10199),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_2 ));
    InMux I__2137 (
            .O(N__10196),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_3 ));
    InMux I__2136 (
            .O(N__10193),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_4 ));
    InMux I__2135 (
            .O(N__10190),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_5 ));
    InMux I__2134 (
            .O(N__10187),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_6 ));
    CascadeMux I__2133 (
            .O(N__10184),
            .I(N__10181));
    InMux I__2132 (
            .O(N__10181),
            .I(N__10175));
    InMux I__2131 (
            .O(N__10180),
            .I(N__10175));
    LocalMux I__2130 (
            .O(N__10175),
            .I(\DUT.uart_inst0.N_100 ));
    CascadeMux I__2129 (
            .O(N__10172),
            .I(N__10166));
    CascadeMux I__2128 (
            .O(N__10171),
            .I(N__10162));
    InMux I__2127 (
            .O(N__10170),
            .I(N__10158));
    InMux I__2126 (
            .O(N__10169),
            .I(N__10155));
    InMux I__2125 (
            .O(N__10166),
            .I(N__10150));
    InMux I__2124 (
            .O(N__10165),
            .I(N__10150));
    InMux I__2123 (
            .O(N__10162),
            .I(N__10147));
    CascadeMux I__2122 (
            .O(N__10161),
            .I(N__10142));
    LocalMux I__2121 (
            .O(N__10158),
            .I(N__10137));
    LocalMux I__2120 (
            .O(N__10155),
            .I(N__10134));
    LocalMux I__2119 (
            .O(N__10150),
            .I(N__10129));
    LocalMux I__2118 (
            .O(N__10147),
            .I(N__10129));
    InMux I__2117 (
            .O(N__10146),
            .I(N__10126));
    InMux I__2116 (
            .O(N__10145),
            .I(N__10123));
    InMux I__2115 (
            .O(N__10142),
            .I(N__10120));
    InMux I__2114 (
            .O(N__10141),
            .I(N__10117));
    CascadeMux I__2113 (
            .O(N__10140),
            .I(N__10112));
    Span4Mux_v I__2112 (
            .O(N__10137),
            .I(N__10108));
    Span4Mux_v I__2111 (
            .O(N__10134),
            .I(N__10105));
    Span4Mux_v I__2110 (
            .O(N__10129),
            .I(N__10102));
    LocalMux I__2109 (
            .O(N__10126),
            .I(N__10095));
    LocalMux I__2108 (
            .O(N__10123),
            .I(N__10095));
    LocalMux I__2107 (
            .O(N__10120),
            .I(N__10095));
    LocalMux I__2106 (
            .O(N__10117),
            .I(N__10092));
    InMux I__2105 (
            .O(N__10116),
            .I(N__10085));
    InMux I__2104 (
            .O(N__10115),
            .I(N__10085));
    InMux I__2103 (
            .O(N__10112),
            .I(N__10085));
    InMux I__2102 (
            .O(N__10111),
            .I(N__10082));
    Span4Mux_v I__2101 (
            .O(N__10108),
            .I(N__10075));
    Span4Mux_v I__2100 (
            .O(N__10105),
            .I(N__10075));
    Span4Mux_v I__2099 (
            .O(N__10102),
            .I(N__10075));
    Span4Mux_v I__2098 (
            .O(N__10095),
            .I(N__10072));
    Span4Mux_h I__2097 (
            .O(N__10092),
            .I(N__10067));
    LocalMux I__2096 (
            .O(N__10085),
            .I(N__10067));
    LocalMux I__2095 (
            .O(N__10082),
            .I(N__10064));
    Sp12to4 I__2094 (
            .O(N__10075),
            .I(N__10061));
    Span4Mux_v I__2093 (
            .O(N__10072),
            .I(N__10056));
    Span4Mux_v I__2092 (
            .O(N__10067),
            .I(N__10056));
    Span12Mux_v I__2091 (
            .O(N__10064),
            .I(N__10049));
    Span12Mux_h I__2090 (
            .O(N__10061),
            .I(N__10049));
    Sp12to4 I__2089 (
            .O(N__10056),
            .I(N__10049));
    Odrv12 I__2088 (
            .O(N__10049),
            .I(P1A1_c));
    CascadeMux I__2087 (
            .O(N__10046),
            .I(N__10042));
    CascadeMux I__2086 (
            .O(N__10045),
            .I(N__10036));
    InMux I__2085 (
            .O(N__10042),
            .I(N__10032));
    InMux I__2084 (
            .O(N__10041),
            .I(N__10029));
    InMux I__2083 (
            .O(N__10040),
            .I(N__10026));
    InMux I__2082 (
            .O(N__10039),
            .I(N__10023));
    InMux I__2081 (
            .O(N__10036),
            .I(N__10020));
    CascadeMux I__2080 (
            .O(N__10035),
            .I(N__10016));
    LocalMux I__2079 (
            .O(N__10032),
            .I(N__10013));
    LocalMux I__2078 (
            .O(N__10029),
            .I(N__10010));
    LocalMux I__2077 (
            .O(N__10026),
            .I(N__10007));
    LocalMux I__2076 (
            .O(N__10023),
            .I(N__10004));
    LocalMux I__2075 (
            .O(N__10020),
            .I(N__10001));
    InMux I__2074 (
            .O(N__10019),
            .I(N__9998));
    InMux I__2073 (
            .O(N__10016),
            .I(N__9995));
    Span4Mux_v I__2072 (
            .O(N__10013),
            .I(N__9988));
    Span4Mux_h I__2071 (
            .O(N__10010),
            .I(N__9988));
    Span4Mux_v I__2070 (
            .O(N__10007),
            .I(N__9988));
    Odrv12 I__2069 (
            .O(N__10004),
            .I(\DUT.uart_inst0.recv_stateZ0Z_5 ));
    Odrv12 I__2068 (
            .O(N__10001),
            .I(\DUT.uart_inst0.recv_stateZ0Z_5 ));
    LocalMux I__2067 (
            .O(N__9998),
            .I(\DUT.uart_inst0.recv_stateZ0Z_5 ));
    LocalMux I__2066 (
            .O(N__9995),
            .I(\DUT.uart_inst0.recv_stateZ0Z_5 ));
    Odrv4 I__2065 (
            .O(N__9988),
            .I(\DUT.uart_inst0.recv_stateZ0Z_5 ));
    InMux I__2064 (
            .O(N__9977),
            .I(N__9973));
    InMux I__2063 (
            .O(N__9976),
            .I(N__9970));
    LocalMux I__2062 (
            .O(N__9973),
            .I(N__9965));
    LocalMux I__2061 (
            .O(N__9970),
            .I(N__9962));
    InMux I__2060 (
            .O(N__9969),
            .I(N__9959));
    InMux I__2059 (
            .O(N__9968),
            .I(N__9956));
    Span4Mux_h I__2058 (
            .O(N__9965),
            .I(N__9953));
    Span4Mux_h I__2057 (
            .O(N__9962),
            .I(N__9950));
    LocalMux I__2056 (
            .O(N__9959),
            .I(N__9947));
    LocalMux I__2055 (
            .O(N__9956),
            .I(\DUT.uart_inst0.recv_stateZ0Z_0 ));
    Odrv4 I__2054 (
            .O(N__9953),
            .I(\DUT.uart_inst0.recv_stateZ0Z_0 ));
    Odrv4 I__2053 (
            .O(N__9950),
            .I(\DUT.uart_inst0.recv_stateZ0Z_0 ));
    Odrv4 I__2052 (
            .O(N__9947),
            .I(\DUT.uart_inst0.recv_stateZ0Z_0 ));
    InMux I__2051 (
            .O(N__9938),
            .I(N__9933));
    InMux I__2050 (
            .O(N__9937),
            .I(N__9928));
    InMux I__2049 (
            .O(N__9936),
            .I(N__9928));
    LocalMux I__2048 (
            .O(N__9933),
            .I(N__9925));
    LocalMux I__2047 (
            .O(N__9928),
            .I(N__9922));
    Span12Mux_v I__2046 (
            .O(N__9925),
            .I(N__9919));
    Span4Mux_h I__2045 (
            .O(N__9922),
            .I(N__9916));
    Odrv12 I__2044 (
            .O(N__9919),
            .I(\DUT.uart_inst0.N_49 ));
    Odrv4 I__2043 (
            .O(N__9916),
            .I(\DUT.uart_inst0.N_49 ));
    InMux I__2042 (
            .O(N__9911),
            .I(N__9908));
    LocalMux I__2041 (
            .O(N__9908),
            .I(N__9905));
    Odrv12 I__2040 (
            .O(N__9905),
            .I(\fifo_inst.ft2232h_inst.rFifoStatec_0 ));
    CascadeMux I__2039 (
            .O(N__9902),
            .I(N__9898));
    CascadeMux I__2038 (
            .O(N__9901),
            .I(N__9893));
    InMux I__2037 (
            .O(N__9898),
            .I(N__9890));
    InMux I__2036 (
            .O(N__9897),
            .I(N__9883));
    InMux I__2035 (
            .O(N__9896),
            .I(N__9883));
    InMux I__2034 (
            .O(N__9893),
            .I(N__9883));
    LocalMux I__2033 (
            .O(N__9890),
            .I(N__9880));
    LocalMux I__2032 (
            .O(N__9883),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_3 ));
    Odrv4 I__2031 (
            .O(N__9880),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_3 ));
    InMux I__2030 (
            .O(N__9875),
            .I(N__9865));
    InMux I__2029 (
            .O(N__9874),
            .I(N__9865));
    InMux I__2028 (
            .O(N__9873),
            .I(N__9865));
    InMux I__2027 (
            .O(N__9872),
            .I(N__9862));
    LocalMux I__2026 (
            .O(N__9865),
            .I(\DUT.uart_inst0.N_139 ));
    LocalMux I__2025 (
            .O(N__9862),
            .I(\DUT.uart_inst0.N_139 ));
    CascadeMux I__2024 (
            .O(N__9857),
            .I(N__9853));
    InMux I__2023 (
            .O(N__9856),
            .I(N__9845));
    InMux I__2022 (
            .O(N__9853),
            .I(N__9845));
    InMux I__2021 (
            .O(N__9852),
            .I(N__9845));
    LocalMux I__2020 (
            .O(N__9845),
            .I(N__9840));
    InMux I__2019 (
            .O(N__9844),
            .I(N__9835));
    InMux I__2018 (
            .O(N__9843),
            .I(N__9835));
    Odrv4 I__2017 (
            .O(N__9840),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_2 ));
    LocalMux I__2016 (
            .O(N__9835),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_2 ));
    InMux I__2015 (
            .O(N__9830),
            .I(N__9826));
    InMux I__2014 (
            .O(N__9829),
            .I(N__9822));
    LocalMux I__2013 (
            .O(N__9826),
            .I(N__9819));
    InMux I__2012 (
            .O(N__9825),
            .I(N__9816));
    LocalMux I__2011 (
            .O(N__9822),
            .I(\DUT.rTransmitc_0 ));
    Odrv4 I__2010 (
            .O(N__9819),
            .I(\DUT.rTransmitc_0 ));
    LocalMux I__2009 (
            .O(N__9816),
            .I(\DUT.rTransmitc_0 ));
    CascadeMux I__2008 (
            .O(N__9809),
            .I(\DUT.uart_inst0.N_85_cascade_ ));
    InMux I__2007 (
            .O(N__9806),
            .I(N__9803));
    LocalMux I__2006 (
            .O(N__9803),
            .I(N__9798));
    InMux I__2005 (
            .O(N__9802),
            .I(N__9795));
    InMux I__2004 (
            .O(N__9801),
            .I(N__9792));
    Odrv4 I__2003 (
            .O(N__9798),
            .I(\DUT.uart_inst0.N_66 ));
    LocalMux I__2002 (
            .O(N__9795),
            .I(\DUT.uart_inst0.N_66 ));
    LocalMux I__2001 (
            .O(N__9792),
            .I(\DUT.uart_inst0.N_66 ));
    CascadeMux I__2000 (
            .O(N__9785),
            .I(\DUT.uart_inst0.N_22_cascade_ ));
    InMux I__1999 (
            .O(N__9782),
            .I(N__9773));
    InMux I__1998 (
            .O(N__9781),
            .I(N__9773));
    InMux I__1997 (
            .O(N__9780),
            .I(N__9773));
    LocalMux I__1996 (
            .O(N__9773),
            .I(N__9766));
    InMux I__1995 (
            .O(N__9772),
            .I(N__9757));
    InMux I__1994 (
            .O(N__9771),
            .I(N__9757));
    InMux I__1993 (
            .O(N__9770),
            .I(N__9757));
    InMux I__1992 (
            .O(N__9769),
            .I(N__9757));
    Odrv4 I__1991 (
            .O(N__9766),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_0 ));
    LocalMux I__1990 (
            .O(N__9757),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_0 ));
    InMux I__1989 (
            .O(N__9752),
            .I(N__9749));
    LocalMux I__1988 (
            .O(N__9749),
            .I(N__9744));
    InMux I__1987 (
            .O(N__9748),
            .I(N__9739));
    InMux I__1986 (
            .O(N__9747),
            .I(N__9739));
    Odrv4 I__1985 (
            .O(N__9744),
            .I(\DUT.uart_inst0.N_22 ));
    LocalMux I__1984 (
            .O(N__9739),
            .I(\DUT.uart_inst0.N_22 ));
    InMux I__1983 (
            .O(N__9734),
            .I(N__9723));
    InMux I__1982 (
            .O(N__9733),
            .I(N__9723));
    InMux I__1981 (
            .O(N__9732),
            .I(N__9723));
    CascadeMux I__1980 (
            .O(N__9731),
            .I(N__9720));
    CascadeMux I__1979 (
            .O(N__9730),
            .I(N__9717));
    LocalMux I__1978 (
            .O(N__9723),
            .I(N__9713));
    InMux I__1977 (
            .O(N__9720),
            .I(N__9706));
    InMux I__1976 (
            .O(N__9717),
            .I(N__9706));
    InMux I__1975 (
            .O(N__9716),
            .I(N__9706));
    Odrv4 I__1974 (
            .O(N__9713),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_1 ));
    LocalMux I__1973 (
            .O(N__9706),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_1 ));
    InMux I__1972 (
            .O(N__9701),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_16 ));
    CascadeMux I__1971 (
            .O(N__9698),
            .I(N__9694));
    InMux I__1970 (
            .O(N__9697),
            .I(N__9691));
    InMux I__1969 (
            .O(N__9694),
            .I(N__9688));
    LocalMux I__1968 (
            .O(N__9691),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_17 ));
    LocalMux I__1967 (
            .O(N__9688),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_17 ));
    InMux I__1966 (
            .O(N__9683),
            .I(N__9680));
    LocalMux I__1965 (
            .O(N__9680),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO ));
    InMux I__1964 (
            .O(N__9677),
            .I(N__9672));
    InMux I__1963 (
            .O(N__9676),
            .I(N__9669));
    InMux I__1962 (
            .O(N__9675),
            .I(N__9666));
    LocalMux I__1961 (
            .O(N__9672),
            .I(N__9661));
    LocalMux I__1960 (
            .O(N__9669),
            .I(N__9661));
    LocalMux I__1959 (
            .O(N__9666),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_12 ));
    Odrv4 I__1958 (
            .O(N__9661),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_12 ));
    InMux I__1957 (
            .O(N__9656),
            .I(N__9653));
    LocalMux I__1956 (
            .O(N__9653),
            .I(N__9650));
    Odrv12 I__1955 (
            .O(N__9650),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO ));
    InMux I__1954 (
            .O(N__9647),
            .I(N__9642));
    InMux I__1953 (
            .O(N__9646),
            .I(N__9639));
    InMux I__1952 (
            .O(N__9645),
            .I(N__9636));
    LocalMux I__1951 (
            .O(N__9642),
            .I(N__9633));
    LocalMux I__1950 (
            .O(N__9639),
            .I(N__9630));
    LocalMux I__1949 (
            .O(N__9636),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_2 ));
    Odrv4 I__1948 (
            .O(N__9633),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_2 ));
    Odrv4 I__1947 (
            .O(N__9630),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_2 ));
    InMux I__1946 (
            .O(N__9623),
            .I(N__9620));
    LocalMux I__1945 (
            .O(N__9620),
            .I(N__9617));
    Odrv4 I__1944 (
            .O(N__9617),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO ));
    CascadeMux I__1943 (
            .O(N__9614),
            .I(N__9602));
    CascadeMux I__1942 (
            .O(N__9613),
            .I(N__9596));
    CascadeMux I__1941 (
            .O(N__9612),
            .I(N__9592));
    InMux I__1940 (
            .O(N__9611),
            .I(N__9581));
    InMux I__1939 (
            .O(N__9610),
            .I(N__9581));
    InMux I__1938 (
            .O(N__9609),
            .I(N__9581));
    InMux I__1937 (
            .O(N__9608),
            .I(N__9581));
    InMux I__1936 (
            .O(N__9607),
            .I(N__9567));
    InMux I__1935 (
            .O(N__9606),
            .I(N__9567));
    InMux I__1934 (
            .O(N__9605),
            .I(N__9567));
    InMux I__1933 (
            .O(N__9602),
            .I(N__9567));
    InMux I__1932 (
            .O(N__9601),
            .I(N__9567));
    InMux I__1931 (
            .O(N__9600),
            .I(N__9567));
    InMux I__1930 (
            .O(N__9599),
            .I(N__9551));
    InMux I__1929 (
            .O(N__9596),
            .I(N__9551));
    InMux I__1928 (
            .O(N__9595),
            .I(N__9551));
    InMux I__1927 (
            .O(N__9592),
            .I(N__9551));
    InMux I__1926 (
            .O(N__9591),
            .I(N__9551));
    InMux I__1925 (
            .O(N__9590),
            .I(N__9551));
    LocalMux I__1924 (
            .O(N__9581),
            .I(N__9548));
    InMux I__1923 (
            .O(N__9580),
            .I(N__9545));
    LocalMux I__1922 (
            .O(N__9567),
            .I(N__9542));
    InMux I__1921 (
            .O(N__9566),
            .I(N__9536));
    InMux I__1920 (
            .O(N__9565),
            .I(N__9533));
    InMux I__1919 (
            .O(N__9564),
            .I(N__9530));
    LocalMux I__1918 (
            .O(N__9551),
            .I(N__9527));
    Span4Mux_h I__1917 (
            .O(N__9548),
            .I(N__9524));
    LocalMux I__1916 (
            .O(N__9545),
            .I(N__9519));
    Span4Mux_h I__1915 (
            .O(N__9542),
            .I(N__9519));
    InMux I__1914 (
            .O(N__9541),
            .I(N__9516));
    InMux I__1913 (
            .O(N__9540),
            .I(N__9511));
    InMux I__1912 (
            .O(N__9539),
            .I(N__9511));
    LocalMux I__1911 (
            .O(N__9536),
            .I(N__9506));
    LocalMux I__1910 (
            .O(N__9533),
            .I(N__9506));
    LocalMux I__1909 (
            .O(N__9530),
            .I(\DUT.uart_inst0.N_50 ));
    Odrv4 I__1908 (
            .O(N__9527),
            .I(\DUT.uart_inst0.N_50 ));
    Odrv4 I__1907 (
            .O(N__9524),
            .I(\DUT.uart_inst0.N_50 ));
    Odrv4 I__1906 (
            .O(N__9519),
            .I(\DUT.uart_inst0.N_50 ));
    LocalMux I__1905 (
            .O(N__9516),
            .I(\DUT.uart_inst0.N_50 ));
    LocalMux I__1904 (
            .O(N__9511),
            .I(\DUT.uart_inst0.N_50 ));
    Odrv4 I__1903 (
            .O(N__9506),
            .I(\DUT.uart_inst0.N_50 ));
    CascadeMux I__1902 (
            .O(N__9491),
            .I(N__9487));
    InMux I__1901 (
            .O(N__9490),
            .I(N__9483));
    InMux I__1900 (
            .O(N__9487),
            .I(N__9480));
    InMux I__1899 (
            .O(N__9486),
            .I(N__9477));
    LocalMux I__1898 (
            .O(N__9483),
            .I(N__9474));
    LocalMux I__1897 (
            .O(N__9480),
            .I(N__9471));
    LocalMux I__1896 (
            .O(N__9477),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_4 ));
    Odrv4 I__1895 (
            .O(N__9474),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_4 ));
    Odrv4 I__1894 (
            .O(N__9471),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_4 ));
    CascadeMux I__1893 (
            .O(N__9464),
            .I(\DUT.uart_inst0.N_98_cascade_ ));
    IoInMux I__1892 (
            .O(N__9461),
            .I(N__9458));
    LocalMux I__1891 (
            .O(N__9458),
            .I(N__9455));
    Span4Mux_s3_v I__1890 (
            .O(N__9455),
            .I(N__9452));
    Span4Mux_v I__1889 (
            .O(N__9452),
            .I(N__9449));
    Span4Mux_v I__1888 (
            .O(N__9449),
            .I(N__9445));
    InMux I__1887 (
            .O(N__9448),
            .I(N__9442));
    Span4Mux_v I__1886 (
            .O(N__9445),
            .I(N__9439));
    LocalMux I__1885 (
            .O(N__9442),
            .I(N__9436));
    Odrv4 I__1884 (
            .O(N__9439),
            .I(P1A7_c));
    Odrv4 I__1883 (
            .O(N__9436),
            .I(P1A7_c));
    InMux I__1882 (
            .O(N__9431),
            .I(N__9428));
    LocalMux I__1881 (
            .O(N__9428),
            .I(\DUT.uart_inst0.N_82 ));
    InMux I__1880 (
            .O(N__9425),
            .I(N__9419));
    InMux I__1879 (
            .O(N__9424),
            .I(N__9419));
    LocalMux I__1878 (
            .O(N__9419),
            .I(\DUT.uart_inst0.N_99 ));
    CascadeMux I__1877 (
            .O(N__9416),
            .I(N__9411));
    InMux I__1876 (
            .O(N__9415),
            .I(N__9408));
    InMux I__1875 (
            .O(N__9414),
            .I(N__9403));
    InMux I__1874 (
            .O(N__9411),
            .I(N__9403));
    LocalMux I__1873 (
            .O(N__9408),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_9 ));
    LocalMux I__1872 (
            .O(N__9403),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_9 ));
    CascadeMux I__1871 (
            .O(N__9398),
            .I(N__9395));
    InMux I__1870 (
            .O(N__9395),
            .I(N__9392));
    LocalMux I__1869 (
            .O(N__9392),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO ));
    InMux I__1868 (
            .O(N__9389),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_8 ));
    InMux I__1867 (
            .O(N__9386),
            .I(N__9381));
    InMux I__1866 (
            .O(N__9385),
            .I(N__9378));
    InMux I__1865 (
            .O(N__9384),
            .I(N__9375));
    LocalMux I__1864 (
            .O(N__9381),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_10 ));
    LocalMux I__1863 (
            .O(N__9378),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_10 ));
    LocalMux I__1862 (
            .O(N__9375),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_10 ));
    InMux I__1861 (
            .O(N__9368),
            .I(N__9365));
    LocalMux I__1860 (
            .O(N__9365),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO ));
    InMux I__1859 (
            .O(N__9362),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_9 ));
    InMux I__1858 (
            .O(N__9359),
            .I(N__9354));
    InMux I__1857 (
            .O(N__9358),
            .I(N__9351));
    InMux I__1856 (
            .O(N__9357),
            .I(N__9348));
    LocalMux I__1855 (
            .O(N__9354),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_11 ));
    LocalMux I__1854 (
            .O(N__9351),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_11 ));
    LocalMux I__1853 (
            .O(N__9348),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_11 ));
    InMux I__1852 (
            .O(N__9341),
            .I(N__9338));
    LocalMux I__1851 (
            .O(N__9338),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO ));
    InMux I__1850 (
            .O(N__9335),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_10 ));
    InMux I__1849 (
            .O(N__9332),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_11 ));
    InMux I__1848 (
            .O(N__9329),
            .I(N__9324));
    InMux I__1847 (
            .O(N__9328),
            .I(N__9319));
    InMux I__1846 (
            .O(N__9327),
            .I(N__9319));
    LocalMux I__1845 (
            .O(N__9324),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_13 ));
    LocalMux I__1844 (
            .O(N__9319),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_13 ));
    InMux I__1843 (
            .O(N__9314),
            .I(N__9311));
    LocalMux I__1842 (
            .O(N__9311),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO ));
    InMux I__1841 (
            .O(N__9308),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_12 ));
    InMux I__1840 (
            .O(N__9305),
            .I(N__9300));
    InMux I__1839 (
            .O(N__9304),
            .I(N__9297));
    InMux I__1838 (
            .O(N__9303),
            .I(N__9294));
    LocalMux I__1837 (
            .O(N__9300),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_14 ));
    LocalMux I__1836 (
            .O(N__9297),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_14 ));
    LocalMux I__1835 (
            .O(N__9294),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_14 ));
    InMux I__1834 (
            .O(N__9287),
            .I(N__9284));
    LocalMux I__1833 (
            .O(N__9284),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO ));
    InMux I__1832 (
            .O(N__9281),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_13 ));
    InMux I__1831 (
            .O(N__9278),
            .I(N__9273));
    InMux I__1830 (
            .O(N__9277),
            .I(N__9268));
    InMux I__1829 (
            .O(N__9276),
            .I(N__9268));
    LocalMux I__1828 (
            .O(N__9273),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_15 ));
    LocalMux I__1827 (
            .O(N__9268),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_15 ));
    InMux I__1826 (
            .O(N__9263),
            .I(N__9260));
    LocalMux I__1825 (
            .O(N__9260),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO ));
    InMux I__1824 (
            .O(N__9257),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_14 ));
    InMux I__1823 (
            .O(N__9254),
            .I(N__9249));
    InMux I__1822 (
            .O(N__9253),
            .I(N__9246));
    InMux I__1821 (
            .O(N__9252),
            .I(N__9243));
    LocalMux I__1820 (
            .O(N__9249),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_16 ));
    LocalMux I__1819 (
            .O(N__9246),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_16 ));
    LocalMux I__1818 (
            .O(N__9243),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_16 ));
    InMux I__1817 (
            .O(N__9236),
            .I(N__9233));
    LocalMux I__1816 (
            .O(N__9233),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO ));
    InMux I__1815 (
            .O(N__9230),
            .I(bfn_11_15_0_));
    InMux I__1814 (
            .O(N__9227),
            .I(N__9224));
    LocalMux I__1813 (
            .O(N__9224),
            .I(N__9221));
    Span4Mux_h I__1812 (
            .O(N__9221),
            .I(N__9216));
    InMux I__1811 (
            .O(N__9220),
            .I(N__9211));
    InMux I__1810 (
            .O(N__9219),
            .I(N__9211));
    Odrv4 I__1809 (
            .O(N__9216),
            .I(\DUT.uart_inst0.rx_clk_dividerZ1Z_1 ));
    LocalMux I__1808 (
            .O(N__9211),
            .I(\DUT.uart_inst0.rx_clk_dividerZ1Z_1 ));
    InMux I__1807 (
            .O(N__9206),
            .I(N__9203));
    LocalMux I__1806 (
            .O(N__9203),
            .I(N__9200));
    Span4Mux_h I__1805 (
            .O(N__9200),
            .I(N__9197));
    Odrv4 I__1804 (
            .O(N__9197),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO ));
    InMux I__1803 (
            .O(N__9194),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_0 ));
    InMux I__1802 (
            .O(N__9191),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_1 ));
    InMux I__1801 (
            .O(N__9188),
            .I(N__9185));
    LocalMux I__1800 (
            .O(N__9185),
            .I(N__9182));
    Span4Mux_h I__1799 (
            .O(N__9182),
            .I(N__9177));
    InMux I__1798 (
            .O(N__9181),
            .I(N__9172));
    InMux I__1797 (
            .O(N__9180),
            .I(N__9172));
    Odrv4 I__1796 (
            .O(N__9177),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_3 ));
    LocalMux I__1795 (
            .O(N__9172),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_3 ));
    CascadeMux I__1794 (
            .O(N__9167),
            .I(N__9164));
    InMux I__1793 (
            .O(N__9164),
            .I(N__9161));
    LocalMux I__1792 (
            .O(N__9161),
            .I(N__9158));
    Span4Mux_v I__1791 (
            .O(N__9158),
            .I(N__9155));
    Span4Mux_h I__1790 (
            .O(N__9155),
            .I(N__9152));
    Odrv4 I__1789 (
            .O(N__9152),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_2_THRU_CO ));
    InMux I__1788 (
            .O(N__9149),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_2 ));
    InMux I__1787 (
            .O(N__9146),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_3 ));
    InMux I__1786 (
            .O(N__9143),
            .I(N__9138));
    InMux I__1785 (
            .O(N__9142),
            .I(N__9133));
    InMux I__1784 (
            .O(N__9141),
            .I(N__9133));
    LocalMux I__1783 (
            .O(N__9138),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_5 ));
    LocalMux I__1782 (
            .O(N__9133),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_5 ));
    InMux I__1781 (
            .O(N__9128),
            .I(N__9125));
    LocalMux I__1780 (
            .O(N__9125),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_4_THRU_CO ));
    InMux I__1779 (
            .O(N__9122),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_4 ));
    CascadeMux I__1778 (
            .O(N__9119),
            .I(N__9115));
    InMux I__1777 (
            .O(N__9118),
            .I(N__9111));
    InMux I__1776 (
            .O(N__9115),
            .I(N__9106));
    InMux I__1775 (
            .O(N__9114),
            .I(N__9106));
    LocalMux I__1774 (
            .O(N__9111),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_6 ));
    LocalMux I__1773 (
            .O(N__9106),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_6 ));
    InMux I__1772 (
            .O(N__9101),
            .I(N__9098));
    LocalMux I__1771 (
            .O(N__9098),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_5_THRU_CO ));
    InMux I__1770 (
            .O(N__9095),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_5 ));
    InMux I__1769 (
            .O(N__9092),
            .I(N__9087));
    InMux I__1768 (
            .O(N__9091),
            .I(N__9084));
    InMux I__1767 (
            .O(N__9090),
            .I(N__9081));
    LocalMux I__1766 (
            .O(N__9087),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_7 ));
    LocalMux I__1765 (
            .O(N__9084),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_7 ));
    LocalMux I__1764 (
            .O(N__9081),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_7 ));
    InMux I__1763 (
            .O(N__9074),
            .I(N__9071));
    LocalMux I__1762 (
            .O(N__9071),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO ));
    InMux I__1761 (
            .O(N__9068),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_6 ));
    CascadeMux I__1760 (
            .O(N__9065),
            .I(N__9060));
    InMux I__1759 (
            .O(N__9064),
            .I(N__9057));
    InMux I__1758 (
            .O(N__9063),
            .I(N__9052));
    InMux I__1757 (
            .O(N__9060),
            .I(N__9052));
    LocalMux I__1756 (
            .O(N__9057),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_8 ));
    LocalMux I__1755 (
            .O(N__9052),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_8 ));
    InMux I__1754 (
            .O(N__9047),
            .I(N__9044));
    LocalMux I__1753 (
            .O(N__9044),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO ));
    InMux I__1752 (
            .O(N__9041),
            .I(bfn_11_14_0_));
    CascadeMux I__1751 (
            .O(N__9038),
            .I(N__9035));
    InMux I__1750 (
            .O(N__9035),
            .I(N__9029));
    InMux I__1749 (
            .O(N__9034),
            .I(N__9029));
    LocalMux I__1748 (
            .O(N__9029),
            .I(\DUT.fifo_tx_inst.un1_i11_2_i ));
    CascadeMux I__1747 (
            .O(N__9026),
            .I(N__9021));
    CascadeMux I__1746 (
            .O(N__9025),
            .I(N__9012));
    CascadeMux I__1745 (
            .O(N__9024),
            .I(N__9006));
    InMux I__1744 (
            .O(N__9021),
            .I(N__9000));
    InMux I__1743 (
            .O(N__9020),
            .I(N__8995));
    InMux I__1742 (
            .O(N__9019),
            .I(N__8995));
    InMux I__1741 (
            .O(N__9018),
            .I(N__8978));
    InMux I__1740 (
            .O(N__9017),
            .I(N__8978));
    InMux I__1739 (
            .O(N__9016),
            .I(N__8978));
    InMux I__1738 (
            .O(N__9015),
            .I(N__8978));
    InMux I__1737 (
            .O(N__9012),
            .I(N__8978));
    InMux I__1736 (
            .O(N__9011),
            .I(N__8978));
    InMux I__1735 (
            .O(N__9010),
            .I(N__8978));
    InMux I__1734 (
            .O(N__9009),
            .I(N__8978));
    InMux I__1733 (
            .O(N__9006),
            .I(N__8969));
    InMux I__1732 (
            .O(N__9005),
            .I(N__8969));
    InMux I__1731 (
            .O(N__9004),
            .I(N__8969));
    CascadeMux I__1730 (
            .O(N__9003),
            .I(N__8965));
    LocalMux I__1729 (
            .O(N__9000),
            .I(N__8961));
    LocalMux I__1728 (
            .O(N__8995),
            .I(N__8956));
    LocalMux I__1727 (
            .O(N__8978),
            .I(N__8956));
    InMux I__1726 (
            .O(N__8977),
            .I(N__8953));
    InMux I__1725 (
            .O(N__8976),
            .I(N__8950));
    LocalMux I__1724 (
            .O(N__8969),
            .I(N__8947));
    CascadeMux I__1723 (
            .O(N__8968),
            .I(N__8943));
    InMux I__1722 (
            .O(N__8965),
            .I(N__8938));
    InMux I__1721 (
            .O(N__8964),
            .I(N__8938));
    Span4Mux_v I__1720 (
            .O(N__8961),
            .I(N__8935));
    Span4Mux_v I__1719 (
            .O(N__8956),
            .I(N__8930));
    LocalMux I__1718 (
            .O(N__8953),
            .I(N__8930));
    LocalMux I__1717 (
            .O(N__8950),
            .I(N__8925));
    Span4Mux_h I__1716 (
            .O(N__8947),
            .I(N__8925));
    InMux I__1715 (
            .O(N__8946),
            .I(N__8920));
    InMux I__1714 (
            .O(N__8943),
            .I(N__8920));
    LocalMux I__1713 (
            .O(N__8938),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    Odrv4 I__1712 (
            .O(N__8935),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    Odrv4 I__1711 (
            .O(N__8930),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    Odrv4 I__1710 (
            .O(N__8925),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__1709 (
            .O(N__8920),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    InMux I__1708 (
            .O(N__8909),
            .I(N__8906));
    LocalMux I__1707 (
            .O(N__8906),
            .I(N__8903));
    Span4Mux_v I__1706 (
            .O(N__8903),
            .I(N__8900));
    Odrv4 I__1705 (
            .O(N__8900),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_1 ));
    CascadeMux I__1704 (
            .O(N__8897),
            .I(N__8894));
    InMux I__1703 (
            .O(N__8894),
            .I(N__8891));
    LocalMux I__1702 (
            .O(N__8891),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_1 ));
    InMux I__1701 (
            .O(N__8888),
            .I(N__8885));
    LocalMux I__1700 (
            .O(N__8885),
            .I(N__8882));
    Odrv12 I__1699 (
            .O(N__8882),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1 ));
    CEMux I__1698 (
            .O(N__8879),
            .I(N__8874));
    CEMux I__1697 (
            .O(N__8878),
            .I(N__8871));
    CEMux I__1696 (
            .O(N__8877),
            .I(N__8868));
    LocalMux I__1695 (
            .O(N__8874),
            .I(N__8865));
    LocalMux I__1694 (
            .O(N__8871),
            .I(N__8862));
    LocalMux I__1693 (
            .O(N__8868),
            .I(N__8859));
    Odrv4 I__1692 (
            .O(N__8865),
            .I(N_92_i_0));
    Odrv4 I__1691 (
            .O(N__8862),
            .I(N_92_i_0));
    Odrv4 I__1690 (
            .O(N__8859),
            .I(N_92_i_0));
    SRMux I__1689 (
            .O(N__8852),
            .I(N__8848));
    SRMux I__1688 (
            .O(N__8851),
            .I(N__8845));
    LocalMux I__1687 (
            .O(N__8848),
            .I(N__8841));
    LocalMux I__1686 (
            .O(N__8845),
            .I(N__8838));
    SRMux I__1685 (
            .O(N__8844),
            .I(N__8835));
    Span4Mux_h I__1684 (
            .O(N__8841),
            .I(N__8832));
    Span4Mux_h I__1683 (
            .O(N__8838),
            .I(N__8829));
    LocalMux I__1682 (
            .O(N__8835),
            .I(N__8826));
    Odrv4 I__1681 (
            .O(N__8832),
            .I(rFifoDatarff_0_RNIHJV05));
    Odrv4 I__1680 (
            .O(N__8829),
            .I(rFifoDatarff_0_RNIHJV05));
    Odrv4 I__1679 (
            .O(N__8826),
            .I(rFifoDatarff_0_RNIHJV05));
    CascadeMux I__1678 (
            .O(N__8819),
            .I(N__8816));
    InMux I__1677 (
            .O(N__8816),
            .I(N__8812));
    InMux I__1676 (
            .O(N__8815),
            .I(N__8809));
    LocalMux I__1675 (
            .O(N__8812),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_2 ));
    LocalMux I__1674 (
            .O(N__8809),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_2 ));
    IoInMux I__1673 (
            .O(N__8804),
            .I(N__8801));
    LocalMux I__1672 (
            .O(N__8801),
            .I(N__8797));
    IoInMux I__1671 (
            .O(N__8800),
            .I(N__8794));
    IoSpan4Mux I__1670 (
            .O(N__8797),
            .I(N__8791));
    LocalMux I__1669 (
            .O(N__8794),
            .I(N__8788));
    Span4Mux_s2_v I__1668 (
            .O(N__8791),
            .I(N__8785));
    IoSpan4Mux I__1667 (
            .O(N__8788),
            .I(N__8782));
    Sp12to4 I__1666 (
            .O(N__8785),
            .I(N__8779));
    Sp12to4 I__1665 (
            .O(N__8782),
            .I(N__8776));
    Span12Mux_s8_v I__1664 (
            .O(N__8779),
            .I(N__8770));
    Span12Mux_s9_v I__1663 (
            .O(N__8776),
            .I(N__8770));
    InMux I__1662 (
            .O(N__8775),
            .I(N__8767));
    Odrv12 I__1661 (
            .O(N__8770),
            .I(P1A4_c));
    LocalMux I__1660 (
            .O(N__8767),
            .I(P1A4_c));
    InMux I__1659 (
            .O(N__8762),
            .I(N__8756));
    InMux I__1658 (
            .O(N__8761),
            .I(N__8756));
    LocalMux I__1657 (
            .O(N__8756),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_3 ));
    IoInMux I__1656 (
            .O(N__8753),
            .I(N__8747));
    IoInMux I__1655 (
            .O(N__8752),
            .I(N__8744));
    IoInMux I__1654 (
            .O(N__8751),
            .I(N__8740));
    IoInMux I__1653 (
            .O(N__8750),
            .I(N__8737));
    LocalMux I__1652 (
            .O(N__8747),
            .I(N__8732));
    LocalMux I__1651 (
            .O(N__8744),
            .I(N__8732));
    IoInMux I__1650 (
            .O(N__8743),
            .I(N__8729));
    LocalMux I__1649 (
            .O(N__8740),
            .I(N__8723));
    LocalMux I__1648 (
            .O(N__8737),
            .I(N__8723));
    IoSpan4Mux I__1647 (
            .O(N__8732),
            .I(N__8717));
    LocalMux I__1646 (
            .O(N__8729),
            .I(N__8717));
    IoInMux I__1645 (
            .O(N__8728),
            .I(N__8714));
    Span4Mux_s2_v I__1644 (
            .O(N__8723),
            .I(N__8711));
    IoInMux I__1643 (
            .O(N__8722),
            .I(N__8708));
    IoSpan4Mux I__1642 (
            .O(N__8717),
            .I(N__8705));
    LocalMux I__1641 (
            .O(N__8714),
            .I(N__8702));
    Span4Mux_h I__1640 (
            .O(N__8711),
            .I(N__8699));
    LocalMux I__1639 (
            .O(N__8708),
            .I(N__8695));
    Span4Mux_s3_v I__1638 (
            .O(N__8705),
            .I(N__8692));
    Span4Mux_s3_v I__1637 (
            .O(N__8702),
            .I(N__8689));
    Span4Mux_v I__1636 (
            .O(N__8699),
            .I(N__8686));
    IoInMux I__1635 (
            .O(N__8698),
            .I(N__8683));
    Span4Mux_s3_v I__1634 (
            .O(N__8695),
            .I(N__8680));
    Sp12to4 I__1633 (
            .O(N__8692),
            .I(N__8674));
    Sp12to4 I__1632 (
            .O(N__8689),
            .I(N__8674));
    Sp12to4 I__1631 (
            .O(N__8686),
            .I(N__8671));
    LocalMux I__1630 (
            .O(N__8683),
            .I(N__8668));
    Span4Mux_v I__1629 (
            .O(N__8680),
            .I(N__8665));
    CascadeMux I__1628 (
            .O(N__8679),
            .I(N__8662));
    Span12Mux_h I__1627 (
            .O(N__8674),
            .I(N__8659));
    Span12Mux_v I__1626 (
            .O(N__8671),
            .I(N__8654));
    Span12Mux_s11_v I__1625 (
            .O(N__8668),
            .I(N__8654));
    Span4Mux_v I__1624 (
            .O(N__8665),
            .I(N__8651));
    InMux I__1623 (
            .O(N__8662),
            .I(N__8648));
    Odrv12 I__1622 (
            .O(N__8659),
            .I(rTxBusReady));
    Odrv12 I__1621 (
            .O(N__8654),
            .I(rTxBusReady));
    Odrv4 I__1620 (
            .O(N__8651),
            .I(rTxBusReady));
    LocalMux I__1619 (
            .O(N__8648),
            .I(rTxBusReady));
    InMux I__1618 (
            .O(N__8639),
            .I(N__8632));
    InMux I__1617 (
            .O(N__8638),
            .I(N__8623));
    InMux I__1616 (
            .O(N__8637),
            .I(N__8623));
    InMux I__1615 (
            .O(N__8636),
            .I(N__8623));
    InMux I__1614 (
            .O(N__8635),
            .I(N__8623));
    LocalMux I__1613 (
            .O(N__8632),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_4 ));
    LocalMux I__1612 (
            .O(N__8623),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_4 ));
    CascadeMux I__1611 (
            .O(N__8618),
            .I(N__8614));
    CascadeMux I__1610 (
            .O(N__8617),
            .I(N__8609));
    InMux I__1609 (
            .O(N__8614),
            .I(N__8601));
    InMux I__1608 (
            .O(N__8613),
            .I(N__8601));
    InMux I__1607 (
            .O(N__8612),
            .I(N__8601));
    InMux I__1606 (
            .O(N__8609),
            .I(N__8596));
    InMux I__1605 (
            .O(N__8608),
            .I(N__8596));
    LocalMux I__1604 (
            .O(N__8601),
            .I(\fifo_inst.ft2232h_inst.rTxRdEnZ0 ));
    LocalMux I__1603 (
            .O(N__8596),
            .I(\fifo_inst.ft2232h_inst.rTxRdEnZ0 ));
    InMux I__1602 (
            .O(N__8591),
            .I(N__8586));
    InMux I__1601 (
            .O(N__8590),
            .I(N__8581));
    InMux I__1600 (
            .O(N__8589),
            .I(N__8581));
    LocalMux I__1599 (
            .O(N__8586),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_1 ));
    LocalMux I__1598 (
            .O(N__8581),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_1 ));
    InMux I__1597 (
            .O(N__8576),
            .I(N__8571));
    InMux I__1596 (
            .O(N__8575),
            .I(N__8563));
    InMux I__1595 (
            .O(N__8574),
            .I(N__8563));
    LocalMux I__1594 (
            .O(N__8571),
            .I(N__8560));
    CascadeMux I__1593 (
            .O(N__8570),
            .I(N__8557));
    InMux I__1592 (
            .O(N__8569),
            .I(N__8552));
    InMux I__1591 (
            .O(N__8568),
            .I(N__8552));
    LocalMux I__1590 (
            .O(N__8563),
            .I(N__8549));
    Span4Mux_v I__1589 (
            .O(N__8560),
            .I(N__8546));
    InMux I__1588 (
            .O(N__8557),
            .I(N__8543));
    LocalMux I__1587 (
            .O(N__8552),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_0 ));
    Odrv12 I__1586 (
            .O(N__8549),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_0 ));
    Odrv4 I__1585 (
            .O(N__8546),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_0 ));
    LocalMux I__1584 (
            .O(N__8543),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_0 ));
    InMux I__1583 (
            .O(N__8534),
            .I(N__8525));
    InMux I__1582 (
            .O(N__8533),
            .I(N__8525));
    InMux I__1581 (
            .O(N__8532),
            .I(N__8522));
    InMux I__1580 (
            .O(N__8531),
            .I(N__8519));
    InMux I__1579 (
            .O(N__8530),
            .I(N__8516));
    LocalMux I__1578 (
            .O(N__8525),
            .I(N__8511));
    LocalMux I__1577 (
            .O(N__8522),
            .I(N__8511));
    LocalMux I__1576 (
            .O(N__8519),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_1 ));
    LocalMux I__1575 (
            .O(N__8516),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_1 ));
    Odrv4 I__1574 (
            .O(N__8511),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_1 ));
    CascadeMux I__1573 (
            .O(N__8504),
            .I(\DUT.fifo_tx_inst.N_83_cascade_ ));
    InMux I__1572 (
            .O(N__8501),
            .I(N__8498));
    LocalMux I__1571 (
            .O(N__8498),
            .I(\DUT.fifo_tx_inst.N_88 ));
    CascadeMux I__1570 (
            .O(N__8495),
            .I(\DUT.fifo_tx_inst.N_88_cascade_ ));
    InMux I__1569 (
            .O(N__8492),
            .I(N__8489));
    LocalMux I__1568 (
            .O(N__8489),
            .I(\DUT.rTransmitc ));
    InMux I__1567 (
            .O(N__8486),
            .I(N__8480));
    InMux I__1566 (
            .O(N__8485),
            .I(N__8480));
    LocalMux I__1565 (
            .O(N__8480),
            .I(N__8477));
    Span4Mux_v I__1564 (
            .O(N__8477),
            .I(N__8471));
    InMux I__1563 (
            .O(N__8476),
            .I(N__8466));
    InMux I__1562 (
            .O(N__8475),
            .I(N__8466));
    InMux I__1561 (
            .O(N__8474),
            .I(N__8463));
    Odrv4 I__1560 (
            .O(N__8471),
            .I(\DUT.fifo_tx_inst.rWritePtr16 ));
    LocalMux I__1559 (
            .O(N__8466),
            .I(\DUT.fifo_tx_inst.rWritePtr16 ));
    LocalMux I__1558 (
            .O(N__8463),
            .I(\DUT.fifo_tx_inst.rWritePtr16 ));
    InMux I__1557 (
            .O(N__8456),
            .I(N__8453));
    LocalMux I__1556 (
            .O(N__8453),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_3 ));
    InMux I__1555 (
            .O(N__8450),
            .I(N__8446));
    InMux I__1554 (
            .O(N__8449),
            .I(N__8443));
    LocalMux I__1553 (
            .O(N__8446),
            .I(\DUT.fifo_tx_inst.rFifoDataro_0 ));
    LocalMux I__1552 (
            .O(N__8443),
            .I(\DUT.fifo_tx_inst.rFifoDataro_0 ));
    CascadeMux I__1551 (
            .O(N__8438),
            .I(N__8434));
    InMux I__1550 (
            .O(N__8437),
            .I(N__8431));
    InMux I__1549 (
            .O(N__8434),
            .I(N__8428));
    LocalMux I__1548 (
            .O(N__8431),
            .I(\DUT.fifo_tx_inst.rFifoDataro_1 ));
    LocalMux I__1547 (
            .O(N__8428),
            .I(\DUT.fifo_tx_inst.rFifoDataro_1 ));
    CascadeMux I__1546 (
            .O(N__8423),
            .I(N__8420));
    InMux I__1545 (
            .O(N__8420),
            .I(N__8417));
    LocalMux I__1544 (
            .O(N__8417),
            .I(\DUT.rFifoDataror_1 ));
    CascadeMux I__1543 (
            .O(N__8414),
            .I(\DUT.rFifoDataror_1_cascade_ ));
    InMux I__1542 (
            .O(N__8411),
            .I(N__8408));
    LocalMux I__1541 (
            .O(N__8408),
            .I(N__8404));
    InMux I__1540 (
            .O(N__8407),
            .I(N__8401));
    Odrv4 I__1539 (
            .O(N__8404),
            .I(\DUT.rFifoDataror_0_0 ));
    LocalMux I__1538 (
            .O(N__8401),
            .I(\DUT.rFifoDataror_0_0 ));
    CascadeMux I__1537 (
            .O(N__8396),
            .I(N__8392));
    InMux I__1536 (
            .O(N__8395),
            .I(N__8382));
    InMux I__1535 (
            .O(N__8392),
            .I(N__8382));
    InMux I__1534 (
            .O(N__8391),
            .I(N__8371));
    InMux I__1533 (
            .O(N__8390),
            .I(N__8371));
    InMux I__1532 (
            .O(N__8389),
            .I(N__8371));
    InMux I__1531 (
            .O(N__8388),
            .I(N__8371));
    InMux I__1530 (
            .O(N__8387),
            .I(N__8371));
    LocalMux I__1529 (
            .O(N__8382),
            .I(N__8366));
    LocalMux I__1528 (
            .O(N__8371),
            .I(N__8366));
    Odrv4 I__1527 (
            .O(N__8366),
            .I(\DUT.rFifoDataror_0 ));
    IoInMux I__1526 (
            .O(N__8363),
            .I(N__8359));
    CascadeMux I__1525 (
            .O(N__8362),
            .I(N__8354));
    LocalMux I__1524 (
            .O(N__8359),
            .I(N__8349));
    InMux I__1523 (
            .O(N__8358),
            .I(N__8343));
    InMux I__1522 (
            .O(N__8357),
            .I(N__8343));
    InMux I__1521 (
            .O(N__8354),
            .I(N__8340));
    InMux I__1520 (
            .O(N__8353),
            .I(N__8337));
    InMux I__1519 (
            .O(N__8352),
            .I(N__8333));
    Span4Mux_s1_v I__1518 (
            .O(N__8349),
            .I(N__8329));
    CascadeMux I__1517 (
            .O(N__8348),
            .I(N__8325));
    LocalMux I__1516 (
            .O(N__8343),
            .I(N__8320));
    LocalMux I__1515 (
            .O(N__8340),
            .I(N__8320));
    LocalMux I__1514 (
            .O(N__8337),
            .I(N__8317));
    InMux I__1513 (
            .O(N__8336),
            .I(N__8314));
    LocalMux I__1512 (
            .O(N__8333),
            .I(N__8311));
    InMux I__1511 (
            .O(N__8332),
            .I(N__8308));
    Sp12to4 I__1510 (
            .O(N__8329),
            .I(N__8305));
    InMux I__1509 (
            .O(N__8328),
            .I(N__8300));
    InMux I__1508 (
            .O(N__8325),
            .I(N__8300));
    Span4Mux_v I__1507 (
            .O(N__8320),
            .I(N__8293));
    Span4Mux_v I__1506 (
            .O(N__8317),
            .I(N__8293));
    LocalMux I__1505 (
            .O(N__8314),
            .I(N__8293));
    Span4Mux_h I__1504 (
            .O(N__8311),
            .I(N__8290));
    LocalMux I__1503 (
            .O(N__8308),
            .I(N__8287));
    Span12Mux_h I__1502 (
            .O(N__8305),
            .I(N__8284));
    LocalMux I__1501 (
            .O(N__8300),
            .I(N__8281));
    Span4Mux_v I__1500 (
            .O(N__8293),
            .I(N__8278));
    Span4Mux_v I__1499 (
            .O(N__8290),
            .I(N__8273));
    Span4Mux_h I__1498 (
            .O(N__8287),
            .I(N__8273));
    Span12Mux_v I__1497 (
            .O(N__8284),
            .I(N__8268));
    Span12Mux_h I__1496 (
            .O(N__8281),
            .I(N__8268));
    Sp12to4 I__1495 (
            .O(N__8278),
            .I(N__8265));
    Sp12to4 I__1494 (
            .O(N__8273),
            .I(N__8262));
    Span12Mux_v I__1493 (
            .O(N__8268),
            .I(N__8259));
    Span12Mux_h I__1492 (
            .O(N__8265),
            .I(N__8256));
    Span12Mux_v I__1491 (
            .O(N__8262),
            .I(N__8253));
    Odrv12 I__1490 (
            .O(N__8259),
            .I(wPllLocked));
    Odrv12 I__1489 (
            .O(N__8256),
            .I(wPllLocked));
    Odrv12 I__1488 (
            .O(N__8253),
            .I(wPllLocked));
    InMux I__1487 (
            .O(N__8246),
            .I(N__8240));
    InMux I__1486 (
            .O(N__8245),
            .I(N__8240));
    LocalMux I__1485 (
            .O(N__8240),
            .I(\DUT.fifo_rx_inst.CO0 ));
    InMux I__1484 (
            .O(N__8237),
            .I(N__8234));
    LocalMux I__1483 (
            .O(N__8234),
            .I(\DUT.fifo_rx_inst.un1_i11_2_i ));
    CascadeMux I__1482 (
            .O(N__8231),
            .I(\DUT.fifo_rx_inst.un1_i11_2_i_cascade_ ));
    InMux I__1481 (
            .O(N__8228),
            .I(N__8224));
    InMux I__1480 (
            .O(N__8227),
            .I(N__8218));
    LocalMux I__1479 (
            .O(N__8224),
            .I(N__8215));
    InMux I__1478 (
            .O(N__8223),
            .I(N__8210));
    InMux I__1477 (
            .O(N__8222),
            .I(N__8210));
    InMux I__1476 (
            .O(N__8221),
            .I(N__8207));
    LocalMux I__1475 (
            .O(N__8218),
            .I(\DUT.fifo_rx_inst.N_92 ));
    Odrv4 I__1474 (
            .O(N__8215),
            .I(\DUT.fifo_rx_inst.N_92 ));
    LocalMux I__1473 (
            .O(N__8210),
            .I(\DUT.fifo_rx_inst.N_92 ));
    LocalMux I__1472 (
            .O(N__8207),
            .I(\DUT.fifo_rx_inst.N_92 ));
    InMux I__1471 (
            .O(N__8198),
            .I(N__8183));
    InMux I__1470 (
            .O(N__8197),
            .I(N__8183));
    InMux I__1469 (
            .O(N__8196),
            .I(N__8183));
    InMux I__1468 (
            .O(N__8195),
            .I(N__8183));
    InMux I__1467 (
            .O(N__8194),
            .I(N__8177));
    InMux I__1466 (
            .O(N__8193),
            .I(N__8177));
    InMux I__1465 (
            .O(N__8192),
            .I(N__8173));
    LocalMux I__1464 (
            .O(N__8183),
            .I(N__8170));
    InMux I__1463 (
            .O(N__8182),
            .I(N__8167));
    LocalMux I__1462 (
            .O(N__8177),
            .I(N__8164));
    InMux I__1461 (
            .O(N__8176),
            .I(N__8158));
    LocalMux I__1460 (
            .O(N__8173),
            .I(N__8155));
    Span4Mux_v I__1459 (
            .O(N__8170),
            .I(N__8150));
    LocalMux I__1458 (
            .O(N__8167),
            .I(N__8150));
    Span4Mux_h I__1457 (
            .O(N__8164),
            .I(N__8147));
    InMux I__1456 (
            .O(N__8163),
            .I(N__8144));
    InMux I__1455 (
            .O(N__8162),
            .I(N__8139));
    InMux I__1454 (
            .O(N__8161),
            .I(N__8139));
    LocalMux I__1453 (
            .O(N__8158),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    Odrv4 I__1452 (
            .O(N__8155),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    Odrv4 I__1451 (
            .O(N__8150),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    Odrv4 I__1450 (
            .O(N__8147),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__1449 (
            .O(N__8144),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__1448 (
            .O(N__8139),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    CascadeMux I__1447 (
            .O(N__8126),
            .I(\DUT.uart_inst0.N_79_cascade_ ));
    InMux I__1446 (
            .O(N__8123),
            .I(N__8120));
    LocalMux I__1445 (
            .O(N__8120),
            .I(N__8117));
    Odrv12 I__1444 (
            .O(N__8117),
            .I(\DUT.uart_inst0.tx_state_ns_i_i_0_0 ));
    CascadeMux I__1443 (
            .O(N__8114),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_ ));
    InMux I__1442 (
            .O(N__8111),
            .I(N__8108));
    LocalMux I__1441 (
            .O(N__8108),
            .I(N__8105));
    Span4Mux_h I__1440 (
            .O(N__8105),
            .I(N__8102));
    Odrv4 I__1439 (
            .O(N__8102),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_2 ));
    InMux I__1438 (
            .O(N__8099),
            .I(N__8096));
    LocalMux I__1437 (
            .O(N__8096),
            .I(N__8093));
    Odrv4 I__1436 (
            .O(N__8093),
            .I(\DUT.rFifoDatarx_2 ));
    InMux I__1435 (
            .O(N__8090),
            .I(N__8087));
    LocalMux I__1434 (
            .O(N__8087),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_2 ));
    InMux I__1433 (
            .O(N__8084),
            .I(N__8081));
    LocalMux I__1432 (
            .O(N__8081),
            .I(N__8078));
    Span4Mux_h I__1431 (
            .O(N__8078),
            .I(N__8075));
    Odrv4 I__1430 (
            .O(N__8075),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_3 ));
    CascadeMux I__1429 (
            .O(N__8072),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ));
    InMux I__1428 (
            .O(N__8069),
            .I(N__8066));
    LocalMux I__1427 (
            .O(N__8066),
            .I(N__8063));
    Odrv4 I__1426 (
            .O(N__8063),
            .I(\DUT.rFifoDatarx_3 ));
    CascadeMux I__1425 (
            .O(N__8060),
            .I(N__8057));
    InMux I__1424 (
            .O(N__8057),
            .I(N__8054));
    LocalMux I__1423 (
            .O(N__8054),
            .I(\DUT.uart_inst0.tx_dataZ0Z_1 ));
    InMux I__1422 (
            .O(N__8051),
            .I(N__8048));
    LocalMux I__1421 (
            .O(N__8048),
            .I(\DUT.uart_inst0.tx_dataZ0Z_2 ));
    InMux I__1420 (
            .O(N__8045),
            .I(N__8042));
    LocalMux I__1419 (
            .O(N__8042),
            .I(\DUT.uart_inst0.tx_dataZ0Z_3 ));
    CascadeMux I__1418 (
            .O(N__8039),
            .I(N__8036));
    InMux I__1417 (
            .O(N__8036),
            .I(N__8033));
    LocalMux I__1416 (
            .O(N__8033),
            .I(\DUT.uart_inst0.tx_dataZ0Z_4 ));
    InMux I__1415 (
            .O(N__8030),
            .I(N__8027));
    LocalMux I__1414 (
            .O(N__8027),
            .I(N__8024));
    Odrv4 I__1413 (
            .O(N__8024),
            .I(\DUT.uart_inst0.tx_dataZ0Z_5 ));
    CascadeMux I__1412 (
            .O(N__8021),
            .I(N__8018));
    InMux I__1411 (
            .O(N__8018),
            .I(N__8015));
    LocalMux I__1410 (
            .O(N__8015),
            .I(\DUT.uart_inst0.tx_dataZ0Z_6 ));
    InMux I__1409 (
            .O(N__8012),
            .I(N__8009));
    LocalMux I__1408 (
            .O(N__8009),
            .I(N__8006));
    Odrv4 I__1407 (
            .O(N__8006),
            .I(\DUT.uart_inst0.tx_dataZ0Z_7 ));
    CEMux I__1406 (
            .O(N__8003),
            .I(N__7999));
    CEMux I__1405 (
            .O(N__8002),
            .I(N__7996));
    LocalMux I__1404 (
            .O(N__7999),
            .I(N__7993));
    LocalMux I__1403 (
            .O(N__7996),
            .I(N__7990));
    Span4Mux_h I__1402 (
            .O(N__7993),
            .I(N__7987));
    Odrv4 I__1401 (
            .O(N__7990),
            .I(\DUT.uart_inst0.N_22_i ));
    Odrv4 I__1400 (
            .O(N__7987),
            .I(\DUT.uart_inst0.N_22_i ));
    CascadeMux I__1399 (
            .O(N__7982),
            .I(\DUT.uart_inst0.g0_i_o6_0_4_cascade_ ));
    InMux I__1398 (
            .O(N__7979),
            .I(N__7976));
    LocalMux I__1397 (
            .O(N__7976),
            .I(\DUT.uart_inst0.g0_i_o6_0_5 ));
    CascadeMux I__1396 (
            .O(N__7973),
            .I(\DUT.uart_inst0.N_139_0_cascade_ ));
    InMux I__1395 (
            .O(N__7970),
            .I(N__7967));
    LocalMux I__1394 (
            .O(N__7967),
            .I(\DUT.uart_inst0.tx_bits_remaining_RNO_1Z0Z_3 ));
    InMux I__1393 (
            .O(N__7964),
            .I(N__7961));
    LocalMux I__1392 (
            .O(N__7961),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_9 ));
    InMux I__1391 (
            .O(N__7958),
            .I(N__7955));
    LocalMux I__1390 (
            .O(N__7955),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_13 ));
    CascadeMux I__1389 (
            .O(N__7952),
            .I(\DUT.uart_inst0.un1_N_5_mux_cascade_ ));
    InMux I__1388 (
            .O(N__7949),
            .I(N__7946));
    LocalMux I__1387 (
            .O(N__7946),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_1 ));
    InMux I__1386 (
            .O(N__7943),
            .I(N__7940));
    LocalMux I__1385 (
            .O(N__7940),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_10 ));
    InMux I__1384 (
            .O(N__7937),
            .I(N__7930));
    InMux I__1383 (
            .O(N__7936),
            .I(N__7930));
    InMux I__1382 (
            .O(N__7935),
            .I(N__7927));
    LocalMux I__1381 (
            .O(N__7930),
            .I(N__7914));
    LocalMux I__1380 (
            .O(N__7927),
            .I(N__7910));
    InMux I__1379 (
            .O(N__7926),
            .I(N__7907));
    InMux I__1378 (
            .O(N__7925),
            .I(N__7904));
    InMux I__1377 (
            .O(N__7924),
            .I(N__7901));
    CascadeMux I__1376 (
            .O(N__7923),
            .I(N__7896));
    InMux I__1375 (
            .O(N__7922),
            .I(N__7888));
    InMux I__1374 (
            .O(N__7921),
            .I(N__7888));
    InMux I__1373 (
            .O(N__7920),
            .I(N__7881));
    InMux I__1372 (
            .O(N__7919),
            .I(N__7881));
    InMux I__1371 (
            .O(N__7918),
            .I(N__7881));
    InMux I__1370 (
            .O(N__7917),
            .I(N__7878));
    Span4Mux_h I__1369 (
            .O(N__7914),
            .I(N__7875));
    InMux I__1368 (
            .O(N__7913),
            .I(N__7872));
    Span4Mux_h I__1367 (
            .O(N__7910),
            .I(N__7863));
    LocalMux I__1366 (
            .O(N__7907),
            .I(N__7863));
    LocalMux I__1365 (
            .O(N__7904),
            .I(N__7863));
    LocalMux I__1364 (
            .O(N__7901),
            .I(N__7863));
    InMux I__1363 (
            .O(N__7900),
            .I(N__7858));
    InMux I__1362 (
            .O(N__7899),
            .I(N__7858));
    InMux I__1361 (
            .O(N__7896),
            .I(N__7851));
    InMux I__1360 (
            .O(N__7895),
            .I(N__7851));
    InMux I__1359 (
            .O(N__7894),
            .I(N__7851));
    InMux I__1358 (
            .O(N__7893),
            .I(N__7848));
    LocalMux I__1357 (
            .O(N__7888),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    LocalMux I__1356 (
            .O(N__7881),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    LocalMux I__1355 (
            .O(N__7878),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    Odrv4 I__1354 (
            .O(N__7875),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    LocalMux I__1353 (
            .O(N__7872),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    Odrv4 I__1352 (
            .O(N__7863),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    LocalMux I__1351 (
            .O(N__7858),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    LocalMux I__1350 (
            .O(N__7851),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    LocalMux I__1349 (
            .O(N__7848),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    InMux I__1348 (
            .O(N__7829),
            .I(N__7826));
    LocalMux I__1347 (
            .O(N__7826),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_11 ));
    CascadeMux I__1346 (
            .O(N__7823),
            .I(N__7820));
    InMux I__1345 (
            .O(N__7820),
            .I(N__7817));
    LocalMux I__1344 (
            .O(N__7817),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_12 ));
    InMux I__1343 (
            .O(N__7814),
            .I(N__7811));
    LocalMux I__1342 (
            .O(N__7811),
            .I(N__7806));
    InMux I__1341 (
            .O(N__7810),
            .I(N__7803));
    InMux I__1340 (
            .O(N__7809),
            .I(N__7799));
    Span4Mux_v I__1339 (
            .O(N__7806),
            .I(N__7794));
    LocalMux I__1338 (
            .O(N__7803),
            .I(N__7794));
    InMux I__1337 (
            .O(N__7802),
            .I(N__7791));
    LocalMux I__1336 (
            .O(N__7799),
            .I(N__7788));
    Span4Mux_v I__1335 (
            .O(N__7794),
            .I(N__7784));
    LocalMux I__1334 (
            .O(N__7791),
            .I(N__7781));
    Span4Mux_h I__1333 (
            .O(N__7788),
            .I(N__7778));
    InMux I__1332 (
            .O(N__7787),
            .I(N__7775));
    Odrv4 I__1331 (
            .O(N__7784),
            .I(\DUT.wRxByte_3 ));
    Odrv12 I__1330 (
            .O(N__7781),
            .I(\DUT.wRxByte_3 ));
    Odrv4 I__1329 (
            .O(N__7778),
            .I(\DUT.wRxByte_3 ));
    LocalMux I__1328 (
            .O(N__7775),
            .I(\DUT.wRxByte_3 ));
    InMux I__1327 (
            .O(N__7766),
            .I(N__7763));
    LocalMux I__1326 (
            .O(N__7763),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_3 ));
    InMux I__1325 (
            .O(N__7760),
            .I(N__7755));
    InMux I__1324 (
            .O(N__7759),
            .I(N__7751));
    InMux I__1323 (
            .O(N__7758),
            .I(N__7748));
    LocalMux I__1322 (
            .O(N__7755),
            .I(N__7745));
    InMux I__1321 (
            .O(N__7754),
            .I(N__7742));
    LocalMux I__1320 (
            .O(N__7751),
            .I(N__7739));
    LocalMux I__1319 (
            .O(N__7748),
            .I(N__7732));
    Span4Mux_h I__1318 (
            .O(N__7745),
            .I(N__7732));
    LocalMux I__1317 (
            .O(N__7742),
            .I(N__7732));
    Span4Mux_v I__1316 (
            .O(N__7739),
            .I(N__7728));
    Span4Mux_v I__1315 (
            .O(N__7732),
            .I(N__7725));
    InMux I__1314 (
            .O(N__7731),
            .I(N__7722));
    Odrv4 I__1313 (
            .O(N__7728),
            .I(\DUT.wRxByte_4 ));
    Odrv4 I__1312 (
            .O(N__7725),
            .I(\DUT.wRxByte_4 ));
    LocalMux I__1311 (
            .O(N__7722),
            .I(\DUT.wRxByte_4 ));
    InMux I__1310 (
            .O(N__7715),
            .I(N__7712));
    LocalMux I__1309 (
            .O(N__7712),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_4 ));
    InMux I__1308 (
            .O(N__7709),
            .I(N__7704));
    InMux I__1307 (
            .O(N__7708),
            .I(N__7700));
    InMux I__1306 (
            .O(N__7707),
            .I(N__7697));
    LocalMux I__1305 (
            .O(N__7704),
            .I(N__7694));
    InMux I__1304 (
            .O(N__7703),
            .I(N__7691));
    LocalMux I__1303 (
            .O(N__7700),
            .I(N__7688));
    LocalMux I__1302 (
            .O(N__7697),
            .I(N__7681));
    Span4Mux_h I__1301 (
            .O(N__7694),
            .I(N__7681));
    LocalMux I__1300 (
            .O(N__7691),
            .I(N__7681));
    Span4Mux_v I__1299 (
            .O(N__7688),
            .I(N__7677));
    Span4Mux_v I__1298 (
            .O(N__7681),
            .I(N__7674));
    InMux I__1297 (
            .O(N__7680),
            .I(N__7671));
    Odrv4 I__1296 (
            .O(N__7677),
            .I(\DUT.wRxByte_5 ));
    Odrv4 I__1295 (
            .O(N__7674),
            .I(\DUT.wRxByte_5 ));
    LocalMux I__1294 (
            .O(N__7671),
            .I(\DUT.wRxByte_5 ));
    InMux I__1293 (
            .O(N__7664),
            .I(N__7661));
    LocalMux I__1292 (
            .O(N__7661),
            .I(N__7658));
    Odrv4 I__1291 (
            .O(N__7658),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_5 ));
    InMux I__1290 (
            .O(N__7655),
            .I(N__7649));
    InMux I__1289 (
            .O(N__7654),
            .I(N__7646));
    InMux I__1288 (
            .O(N__7653),
            .I(N__7643));
    InMux I__1287 (
            .O(N__7652),
            .I(N__7640));
    LocalMux I__1286 (
            .O(N__7649),
            .I(N__7637));
    LocalMux I__1285 (
            .O(N__7646),
            .I(N__7632));
    LocalMux I__1284 (
            .O(N__7643),
            .I(N__7632));
    LocalMux I__1283 (
            .O(N__7640),
            .I(N__7629));
    Span4Mux_h I__1282 (
            .O(N__7637),
            .I(N__7625));
    Span4Mux_v I__1281 (
            .O(N__7632),
            .I(N__7620));
    Span4Mux_h I__1280 (
            .O(N__7629),
            .I(N__7620));
    InMux I__1279 (
            .O(N__7628),
            .I(N__7617));
    Odrv4 I__1278 (
            .O(N__7625),
            .I(\DUT.wRxByte_6 ));
    Odrv4 I__1277 (
            .O(N__7620),
            .I(\DUT.wRxByte_6 ));
    LocalMux I__1276 (
            .O(N__7617),
            .I(\DUT.wRxByte_6 ));
    InMux I__1275 (
            .O(N__7610),
            .I(N__7607));
    LocalMux I__1274 (
            .O(N__7607),
            .I(N__7604));
    Span4Mux_v I__1273 (
            .O(N__7604),
            .I(N__7601));
    Odrv4 I__1272 (
            .O(N__7601),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_6 ));
    CascadeMux I__1271 (
            .O(N__7598),
            .I(N__7595));
    InMux I__1270 (
            .O(N__7595),
            .I(N__7592));
    LocalMux I__1269 (
            .O(N__7592),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_7 ));
    CEMux I__1268 (
            .O(N__7589),
            .I(N__7586));
    LocalMux I__1267 (
            .O(N__7586),
            .I(N__7582));
    InMux I__1266 (
            .O(N__7585),
            .I(N__7579));
    Span4Mux_v I__1265 (
            .O(N__7582),
            .I(N__7576));
    LocalMux I__1264 (
            .O(N__7579),
            .I(N__7573));
    Span4Mux_h I__1263 (
            .O(N__7576),
            .I(N__7570));
    Span4Mux_h I__1262 (
            .O(N__7573),
            .I(N__7567));
    Odrv4 I__1261 (
            .O(N__7570),
            .I(\DUT.fifo_rx_inst.rFifoData_awe3 ));
    Odrv4 I__1260 (
            .O(N__7567),
            .I(\DUT.fifo_rx_inst.rFifoData_awe3 ));
    InMux I__1259 (
            .O(N__7562),
            .I(N__7559));
    LocalMux I__1258 (
            .O(N__7559),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_7 ));
    InMux I__1257 (
            .O(N__7556),
            .I(N__7553));
    LocalMux I__1256 (
            .O(N__7553),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7 ));
    IoInMux I__1255 (
            .O(N__7550),
            .I(N__7547));
    LocalMux I__1254 (
            .O(N__7547),
            .I(N__7543));
    IoInMux I__1253 (
            .O(N__7546),
            .I(N__7540));
    IoSpan4Mux I__1252 (
            .O(N__7543),
            .I(N__7537));
    LocalMux I__1251 (
            .O(N__7540),
            .I(N__7534));
    IoSpan4Mux I__1250 (
            .O(N__7537),
            .I(N__7531));
    Span4Mux_s3_v I__1249 (
            .O(N__7534),
            .I(N__7528));
    Span4Mux_s3_v I__1248 (
            .O(N__7531),
            .I(N__7523));
    Span4Mux_h I__1247 (
            .O(N__7528),
            .I(N__7523));
    Sp12to4 I__1246 (
            .O(N__7523),
            .I(N__7519));
    InMux I__1245 (
            .O(N__7522),
            .I(N__7516));
    Odrv12 I__1244 (
            .O(N__7519),
            .I(P1A3_c));
    LocalMux I__1243 (
            .O(N__7516),
            .I(P1A3_c));
    CEMux I__1242 (
            .O(N__7511),
            .I(N__7508));
    LocalMux I__1241 (
            .O(N__7508),
            .I(N__7504));
    InMux I__1240 (
            .O(N__7507),
            .I(N__7501));
    Odrv12 I__1239 (
            .O(N__7504),
            .I(\DUT.fifo_rx_inst.rFifoData_awe1 ));
    LocalMux I__1238 (
            .O(N__7501),
            .I(\DUT.fifo_rx_inst.rFifoData_awe1 ));
    InMux I__1237 (
            .O(N__7496),
            .I(N__7490));
    InMux I__1236 (
            .O(N__7495),
            .I(N__7490));
    LocalMux I__1235 (
            .O(N__7490),
            .I(\DUT.fifo_rx_inst.rFifoDataro_1 ));
    CEMux I__1234 (
            .O(N__7487),
            .I(N__7484));
    LocalMux I__1233 (
            .O(N__7484),
            .I(N__7481));
    Span4Mux_h I__1232 (
            .O(N__7481),
            .I(N__7477));
    InMux I__1231 (
            .O(N__7480),
            .I(N__7474));
    Odrv4 I__1230 (
            .O(N__7477),
            .I(\DUT.fifo_rx_inst.rFifoData_awe2 ));
    LocalMux I__1229 (
            .O(N__7474),
            .I(\DUT.fifo_rx_inst.rFifoData_awe2 ));
    InMux I__1228 (
            .O(N__7469),
            .I(N__7463));
    InMux I__1227 (
            .O(N__7468),
            .I(N__7463));
    LocalMux I__1226 (
            .O(N__7463),
            .I(\DUT.fifo_rx_inst.rFifoDataro_3 ));
    CascadeMux I__1225 (
            .O(N__7460),
            .I(N__7456));
    InMux I__1224 (
            .O(N__7459),
            .I(N__7451));
    InMux I__1223 (
            .O(N__7456),
            .I(N__7451));
    LocalMux I__1222 (
            .O(N__7451),
            .I(\DUT.fifo_rx_inst.rFifoDataro_2 ));
    InMux I__1221 (
            .O(N__7448),
            .I(N__7445));
    LocalMux I__1220 (
            .O(N__7445),
            .I(\DUT.fifo_rx_inst.rTxByte_42_1 ));
    CascadeMux I__1219 (
            .O(N__7442),
            .I(\DUT.fifo_rx_inst.rTxByte_42_0_cascade_ ));
    InMux I__1218 (
            .O(N__7439),
            .I(N__7436));
    LocalMux I__1217 (
            .O(N__7436),
            .I(N__7433));
    Odrv4 I__1216 (
            .O(N__7433),
            .I(N_92_i));
    CascadeMux I__1215 (
            .O(N__7430),
            .I(rFifoDatarff_0_RNIHJV05_cascade_));
    InMux I__1214 (
            .O(N__7427),
            .I(N__7423));
    InMux I__1213 (
            .O(N__7426),
            .I(N__7419));
    LocalMux I__1212 (
            .O(N__7423),
            .I(N__7415));
    InMux I__1211 (
            .O(N__7422),
            .I(N__7412));
    LocalMux I__1210 (
            .O(N__7419),
            .I(N__7409));
    InMux I__1209 (
            .O(N__7418),
            .I(N__7406));
    Span4Mux_v I__1208 (
            .O(N__7415),
            .I(N__7401));
    LocalMux I__1207 (
            .O(N__7412),
            .I(N__7401));
    Span4Mux_v I__1206 (
            .O(N__7409),
            .I(N__7396));
    LocalMux I__1205 (
            .O(N__7406),
            .I(N__7396));
    Span4Mux_v I__1204 (
            .O(N__7401),
            .I(N__7393));
    Span4Mux_h I__1203 (
            .O(N__7396),
            .I(N__7390));
    Odrv4 I__1202 (
            .O(N__7393),
            .I(\DUT.wRxByte_0 ));
    Odrv4 I__1201 (
            .O(N__7390),
            .I(\DUT.wRxByte_0 ));
    InMux I__1200 (
            .O(N__7385),
            .I(N__7382));
    LocalMux I__1199 (
            .O(N__7382),
            .I(N__7379));
    Odrv4 I__1198 (
            .O(N__7379),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_0 ));
    InMux I__1197 (
            .O(N__7376),
            .I(N__7371));
    InMux I__1196 (
            .O(N__7375),
            .I(N__7367));
    InMux I__1195 (
            .O(N__7374),
            .I(N__7364));
    LocalMux I__1194 (
            .O(N__7371),
            .I(N__7361));
    InMux I__1193 (
            .O(N__7370),
            .I(N__7358));
    LocalMux I__1192 (
            .O(N__7367),
            .I(N__7355));
    LocalMux I__1191 (
            .O(N__7364),
            .I(N__7352));
    Span4Mux_v I__1190 (
            .O(N__7361),
            .I(N__7348));
    LocalMux I__1189 (
            .O(N__7358),
            .I(N__7345));
    Span4Mux_v I__1188 (
            .O(N__7355),
            .I(N__7340));
    Span4Mux_h I__1187 (
            .O(N__7352),
            .I(N__7340));
    InMux I__1186 (
            .O(N__7351),
            .I(N__7337));
    Odrv4 I__1185 (
            .O(N__7348),
            .I(\DUT.wRxByte_1 ));
    Odrv12 I__1184 (
            .O(N__7345),
            .I(\DUT.wRxByte_1 ));
    Odrv4 I__1183 (
            .O(N__7340),
            .I(\DUT.wRxByte_1 ));
    LocalMux I__1182 (
            .O(N__7337),
            .I(\DUT.wRxByte_1 ));
    InMux I__1181 (
            .O(N__7328),
            .I(N__7323));
    InMux I__1180 (
            .O(N__7327),
            .I(N__7320));
    InMux I__1179 (
            .O(N__7326),
            .I(N__7316));
    LocalMux I__1178 (
            .O(N__7323),
            .I(N__7313));
    LocalMux I__1177 (
            .O(N__7320),
            .I(N__7310));
    InMux I__1176 (
            .O(N__7319),
            .I(N__7307));
    LocalMux I__1175 (
            .O(N__7316),
            .I(N__7304));
    Span4Mux_v I__1174 (
            .O(N__7313),
            .I(N__7298));
    Span4Mux_h I__1173 (
            .O(N__7310),
            .I(N__7298));
    LocalMux I__1172 (
            .O(N__7307),
            .I(N__7295));
    Span4Mux_h I__1171 (
            .O(N__7304),
            .I(N__7292));
    InMux I__1170 (
            .O(N__7303),
            .I(N__7289));
    Odrv4 I__1169 (
            .O(N__7298),
            .I(\DUT.wRxByte_2 ));
    Odrv12 I__1168 (
            .O(N__7295),
            .I(\DUT.wRxByte_2 ));
    Odrv4 I__1167 (
            .O(N__7292),
            .I(\DUT.wRxByte_2 ));
    LocalMux I__1166 (
            .O(N__7289),
            .I(\DUT.wRxByte_2 ));
    InMux I__1165 (
            .O(N__7280),
            .I(N__7277));
    LocalMux I__1164 (
            .O(N__7277),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_2 ));
    InMux I__1163 (
            .O(N__7274),
            .I(N__7268));
    InMux I__1162 (
            .O(N__7273),
            .I(N__7259));
    InMux I__1161 (
            .O(N__7272),
            .I(N__7259));
    InMux I__1160 (
            .O(N__7271),
            .I(N__7256));
    LocalMux I__1159 (
            .O(N__7268),
            .I(N__7253));
    InMux I__1158 (
            .O(N__7267),
            .I(N__7244));
    InMux I__1157 (
            .O(N__7266),
            .I(N__7244));
    InMux I__1156 (
            .O(N__7265),
            .I(N__7244));
    InMux I__1155 (
            .O(N__7264),
            .I(N__7244));
    LocalMux I__1154 (
            .O(N__7259),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ));
    LocalMux I__1153 (
            .O(N__7256),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ));
    Odrv4 I__1152 (
            .O(N__7253),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ));
    LocalMux I__1151 (
            .O(N__7244),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ));
    CascadeMux I__1150 (
            .O(N__7235),
            .I(N__7230));
    InMux I__1149 (
            .O(N__7234),
            .I(N__7225));
    InMux I__1148 (
            .O(N__7233),
            .I(N__7222));
    InMux I__1147 (
            .O(N__7230),
            .I(N__7217));
    InMux I__1146 (
            .O(N__7229),
            .I(N__7217));
    InMux I__1145 (
            .O(N__7228),
            .I(N__7214));
    LocalMux I__1144 (
            .O(N__7225),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_1 ));
    LocalMux I__1143 (
            .O(N__7222),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_1 ));
    LocalMux I__1142 (
            .O(N__7217),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_1 ));
    LocalMux I__1141 (
            .O(N__7214),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_1 ));
    CEMux I__1140 (
            .O(N__7205),
            .I(N__7202));
    LocalMux I__1139 (
            .O(N__7202),
            .I(N__7199));
    Span4Mux_h I__1138 (
            .O(N__7199),
            .I(N__7196));
    Odrv4 I__1137 (
            .O(N__7196),
            .I(\DUT.fifo_tx_inst.rFifoData_awe2 ));
    CascadeMux I__1136 (
            .O(N__7193),
            .I(\DUT.fifo_tx_inst.rFifoData_awe2_cascade_ ));
    InMux I__1135 (
            .O(N__7190),
            .I(N__7184));
    InMux I__1134 (
            .O(N__7189),
            .I(N__7184));
    LocalMux I__1133 (
            .O(N__7184),
            .I(\DUT.fifo_tx_inst.rFifoDataro_3 ));
    InMux I__1132 (
            .O(N__7181),
            .I(N__7175));
    InMux I__1131 (
            .O(N__7180),
            .I(N__7175));
    LocalMux I__1130 (
            .O(N__7175),
            .I(\DUT.fifo_tx_inst.rFifoDataro_2 ));
    CascadeMux I__1129 (
            .O(N__7172),
            .I(\DUT.fifo_tx_inst.rFifoData_awe0_cascade_ ));
    InMux I__1128 (
            .O(N__7169),
            .I(N__7163));
    InMux I__1127 (
            .O(N__7168),
            .I(N__7163));
    LocalMux I__1126 (
            .O(N__7163),
            .I(\DUT.fifo_rx_inst.rFifoDataro_0 ));
    CEMux I__1125 (
            .O(N__7160),
            .I(N__7157));
    LocalMux I__1124 (
            .O(N__7157),
            .I(N__7154));
    Odrv12 I__1123 (
            .O(N__7154),
            .I(\DUT.uart_inst0.rx_bits_remaining_2_sqmuxa ));
    CascadeMux I__1122 (
            .O(N__7151),
            .I(\DUT.fifo_rx_inst.N_87_cascade_ ));
    InMux I__1121 (
            .O(N__7148),
            .I(N__7145));
    LocalMux I__1120 (
            .O(N__7145),
            .I(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0 ));
    InMux I__1119 (
            .O(N__7142),
            .I(N__7135));
    CascadeMux I__1118 (
            .O(N__7141),
            .I(N__7132));
    InMux I__1117 (
            .O(N__7140),
            .I(N__7127));
    InMux I__1116 (
            .O(N__7139),
            .I(N__7122));
    InMux I__1115 (
            .O(N__7138),
            .I(N__7122));
    LocalMux I__1114 (
            .O(N__7135),
            .I(N__7119));
    InMux I__1113 (
            .O(N__7132),
            .I(N__7112));
    InMux I__1112 (
            .O(N__7131),
            .I(N__7112));
    InMux I__1111 (
            .O(N__7130),
            .I(N__7112));
    LocalMux I__1110 (
            .O(N__7127),
            .I(N__7107));
    LocalMux I__1109 (
            .O(N__7122),
            .I(N__7107));
    Span4Mux_v I__1108 (
            .O(N__7119),
            .I(N__7099));
    LocalMux I__1107 (
            .O(N__7112),
            .I(N__7099));
    Span4Mux_h I__1106 (
            .O(N__7107),
            .I(N__7099));
    InMux I__1105 (
            .O(N__7106),
            .I(N__7096));
    Sp12to4 I__1104 (
            .O(N__7099),
            .I(N__7091));
    LocalMux I__1103 (
            .O(N__7096),
            .I(N__7091));
    Odrv12 I__1102 (
            .O(N__7091),
            .I(\DUT.wRcvd ));
    CascadeMux I__1101 (
            .O(N__7088),
            .I(N__7085));
    InMux I__1100 (
            .O(N__7085),
            .I(N__7082));
    LocalMux I__1099 (
            .O(N__7082),
            .I(\DUT.fifo_rx_inst.N_87 ));
    CascadeMux I__1098 (
            .O(N__7079),
            .I(\DUT.fifo_rx_inst.N_92_cascade_ ));
    CascadeMux I__1097 (
            .O(N__7076),
            .I(N__7073));
    InMux I__1096 (
            .O(N__7073),
            .I(N__7065));
    InMux I__1095 (
            .O(N__7072),
            .I(N__7062));
    InMux I__1094 (
            .O(N__7071),
            .I(N__7053));
    InMux I__1093 (
            .O(N__7070),
            .I(N__7053));
    InMux I__1092 (
            .O(N__7069),
            .I(N__7053));
    InMux I__1091 (
            .O(N__7068),
            .I(N__7053));
    LocalMux I__1090 (
            .O(N__7065),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_0 ));
    LocalMux I__1089 (
            .O(N__7062),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_0 ));
    LocalMux I__1088 (
            .O(N__7053),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_0 ));
    CascadeMux I__1087 (
            .O(N__7046),
            .I(\DUT.fifo_tx_inst.rFifoData_awe3_cascade_ ));
    InMux I__1086 (
            .O(N__7043),
            .I(N__7040));
    LocalMux I__1085 (
            .O(N__7040),
            .I(\DUT.fifo_tx_inst.un1_i11_i ));
    CascadeMux I__1084 (
            .O(N__7037),
            .I(\DUT.fifo_tx_inst.un1_i11_i_cascade_ ));
    CascadeMux I__1083 (
            .O(N__7034),
            .I(N__7026));
    CascadeMux I__1082 (
            .O(N__7033),
            .I(N__7023));
    CascadeMux I__1081 (
            .O(N__7032),
            .I(N__7020));
    InMux I__1080 (
            .O(N__7031),
            .I(N__7013));
    InMux I__1079 (
            .O(N__7030),
            .I(N__7013));
    InMux I__1078 (
            .O(N__7029),
            .I(N__7010));
    InMux I__1077 (
            .O(N__7026),
            .I(N__7003));
    InMux I__1076 (
            .O(N__7023),
            .I(N__7003));
    InMux I__1075 (
            .O(N__7020),
            .I(N__7003));
    CascadeMux I__1074 (
            .O(N__7019),
            .I(N__6999));
    CascadeMux I__1073 (
            .O(N__7018),
            .I(N__6995));
    LocalMux I__1072 (
            .O(N__7013),
            .I(N__6986));
    LocalMux I__1071 (
            .O(N__7010),
            .I(N__6986));
    LocalMux I__1070 (
            .O(N__7003),
            .I(N__6986));
    InMux I__1069 (
            .O(N__7002),
            .I(N__6981));
    InMux I__1068 (
            .O(N__6999),
            .I(N__6981));
    InMux I__1067 (
            .O(N__6998),
            .I(N__6974));
    InMux I__1066 (
            .O(N__6995),
            .I(N__6974));
    InMux I__1065 (
            .O(N__6994),
            .I(N__6974));
    InMux I__1064 (
            .O(N__6993),
            .I(N__6971));
    Span4Mux_v I__1063 (
            .O(N__6986),
            .I(N__6966));
    LocalMux I__1062 (
            .O(N__6981),
            .I(N__6966));
    LocalMux I__1061 (
            .O(N__6974),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_4 ));
    LocalMux I__1060 (
            .O(N__6971),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_4 ));
    Odrv4 I__1059 (
            .O(N__6966),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_4 ));
    CascadeMux I__1058 (
            .O(N__6959),
            .I(N__6956));
    InMux I__1057 (
            .O(N__6956),
            .I(N__6948));
    InMux I__1056 (
            .O(N__6955),
            .I(N__6948));
    InMux I__1055 (
            .O(N__6954),
            .I(N__6942));
    InMux I__1054 (
            .O(N__6953),
            .I(N__6942));
    LocalMux I__1053 (
            .O(N__6948),
            .I(N__6932));
    CascadeMux I__1052 (
            .O(N__6947),
            .I(N__6929));
    LocalMux I__1051 (
            .O(N__6942),
            .I(N__6926));
    InMux I__1050 (
            .O(N__6941),
            .I(N__6923));
    InMux I__1049 (
            .O(N__6940),
            .I(N__6918));
    InMux I__1048 (
            .O(N__6939),
            .I(N__6918));
    InMux I__1047 (
            .O(N__6938),
            .I(N__6909));
    InMux I__1046 (
            .O(N__6937),
            .I(N__6909));
    InMux I__1045 (
            .O(N__6936),
            .I(N__6909));
    InMux I__1044 (
            .O(N__6935),
            .I(N__6909));
    Span4Mux_h I__1043 (
            .O(N__6932),
            .I(N__6906));
    InMux I__1042 (
            .O(N__6929),
            .I(N__6903));
    Odrv4 I__1041 (
            .O(N__6926),
            .I(\DUT.uart_inst0.rx_countdownZ1Z_3 ));
    LocalMux I__1040 (
            .O(N__6923),
            .I(\DUT.uart_inst0.rx_countdownZ1Z_3 ));
    LocalMux I__1039 (
            .O(N__6918),
            .I(\DUT.uart_inst0.rx_countdownZ1Z_3 ));
    LocalMux I__1038 (
            .O(N__6909),
            .I(\DUT.uart_inst0.rx_countdownZ1Z_3 ));
    Odrv4 I__1037 (
            .O(N__6906),
            .I(\DUT.uart_inst0.rx_countdownZ1Z_3 ));
    LocalMux I__1036 (
            .O(N__6903),
            .I(\DUT.uart_inst0.rx_countdownZ1Z_3 ));
    CascadeMux I__1035 (
            .O(N__6890),
            .I(N__6886));
    CascadeMux I__1034 (
            .O(N__6889),
            .I(N__6883));
    InMux I__1033 (
            .O(N__6886),
            .I(N__6880));
    InMux I__1032 (
            .O(N__6883),
            .I(N__6877));
    LocalMux I__1031 (
            .O(N__6880),
            .I(\DUT.uart_inst0.N_13_mux ));
    LocalMux I__1030 (
            .O(N__6877),
            .I(\DUT.uart_inst0.N_13_mux ));
    InMux I__1029 (
            .O(N__6872),
            .I(N__6864));
    InMux I__1028 (
            .O(N__6871),
            .I(N__6864));
    InMux I__1027 (
            .O(N__6870),
            .I(N__6859));
    CascadeMux I__1026 (
            .O(N__6869),
            .I(N__6855));
    LocalMux I__1025 (
            .O(N__6864),
            .I(N__6848));
    InMux I__1024 (
            .O(N__6863),
            .I(N__6843));
    InMux I__1023 (
            .O(N__6862),
            .I(N__6843));
    LocalMux I__1022 (
            .O(N__6859),
            .I(N__6840));
    InMux I__1021 (
            .O(N__6858),
            .I(N__6837));
    InMux I__1020 (
            .O(N__6855),
            .I(N__6834));
    InMux I__1019 (
            .O(N__6854),
            .I(N__6831));
    InMux I__1018 (
            .O(N__6853),
            .I(N__6828));
    InMux I__1017 (
            .O(N__6852),
            .I(N__6823));
    InMux I__1016 (
            .O(N__6851),
            .I(N__6823));
    Span4Mux_h I__1015 (
            .O(N__6848),
            .I(N__6818));
    LocalMux I__1014 (
            .O(N__6843),
            .I(N__6818));
    Span4Mux_v I__1013 (
            .O(N__6840),
            .I(N__6813));
    LocalMux I__1012 (
            .O(N__6837),
            .I(N__6813));
    LocalMux I__1011 (
            .O(N__6834),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_2 ));
    LocalMux I__1010 (
            .O(N__6831),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_2 ));
    LocalMux I__1009 (
            .O(N__6828),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_2 ));
    LocalMux I__1008 (
            .O(N__6823),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_2 ));
    Odrv4 I__1007 (
            .O(N__6818),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_2 ));
    Odrv4 I__1006 (
            .O(N__6813),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_2 ));
    InMux I__1005 (
            .O(N__6800),
            .I(N__6797));
    LocalMux I__1004 (
            .O(N__6797),
            .I(N__6785));
    CascadeMux I__1003 (
            .O(N__6796),
            .I(N__6782));
    InMux I__1002 (
            .O(N__6795),
            .I(N__6777));
    InMux I__1001 (
            .O(N__6794),
            .I(N__6768));
    InMux I__1000 (
            .O(N__6793),
            .I(N__6768));
    InMux I__999 (
            .O(N__6792),
            .I(N__6768));
    InMux I__998 (
            .O(N__6791),
            .I(N__6768));
    InMux I__997 (
            .O(N__6790),
            .I(N__6765));
    InMux I__996 (
            .O(N__6789),
            .I(N__6760));
    InMux I__995 (
            .O(N__6788),
            .I(N__6760));
    Span4Mux_h I__994 (
            .O(N__6785),
            .I(N__6757));
    InMux I__993 (
            .O(N__6782),
            .I(N__6754));
    InMux I__992 (
            .O(N__6781),
            .I(N__6749));
    InMux I__991 (
            .O(N__6780),
            .I(N__6749));
    LocalMux I__990 (
            .O(N__6777),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_5 ));
    LocalMux I__989 (
            .O(N__6768),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_5 ));
    LocalMux I__988 (
            .O(N__6765),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_5 ));
    LocalMux I__987 (
            .O(N__6760),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_5 ));
    Odrv4 I__986 (
            .O(N__6757),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_5 ));
    LocalMux I__985 (
            .O(N__6754),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_5 ));
    LocalMux I__984 (
            .O(N__6749),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_5 ));
    InMux I__983 (
            .O(N__6734),
            .I(N__6726));
    CascadeMux I__982 (
            .O(N__6733),
            .I(N__6723));
    CascadeMux I__981 (
            .O(N__6732),
            .I(N__6720));
    InMux I__980 (
            .O(N__6731),
            .I(N__6714));
    InMux I__979 (
            .O(N__6730),
            .I(N__6714));
    CascadeMux I__978 (
            .O(N__6729),
            .I(N__6708));
    LocalMux I__977 (
            .O(N__6726),
            .I(N__6705));
    InMux I__976 (
            .O(N__6723),
            .I(N__6700));
    InMux I__975 (
            .O(N__6720),
            .I(N__6700));
    InMux I__974 (
            .O(N__6719),
            .I(N__6692));
    LocalMux I__973 (
            .O(N__6714),
            .I(N__6689));
    InMux I__972 (
            .O(N__6713),
            .I(N__6680));
    InMux I__971 (
            .O(N__6712),
            .I(N__6680));
    CascadeMux I__970 (
            .O(N__6711),
            .I(N__6675));
    InMux I__969 (
            .O(N__6708),
            .I(N__6672));
    Span4Mux_h I__968 (
            .O(N__6705),
            .I(N__6669));
    LocalMux I__967 (
            .O(N__6700),
            .I(N__6666));
    InMux I__966 (
            .O(N__6699),
            .I(N__6659));
    InMux I__965 (
            .O(N__6698),
            .I(N__6659));
    InMux I__964 (
            .O(N__6697),
            .I(N__6659));
    InMux I__963 (
            .O(N__6696),
            .I(N__6654));
    InMux I__962 (
            .O(N__6695),
            .I(N__6654));
    LocalMux I__961 (
            .O(N__6692),
            .I(N__6649));
    Span4Mux_h I__960 (
            .O(N__6689),
            .I(N__6649));
    InMux I__959 (
            .O(N__6688),
            .I(N__6644));
    InMux I__958 (
            .O(N__6687),
            .I(N__6644));
    InMux I__957 (
            .O(N__6686),
            .I(N__6639));
    InMux I__956 (
            .O(N__6685),
            .I(N__6639));
    LocalMux I__955 (
            .O(N__6680),
            .I(N__6636));
    InMux I__954 (
            .O(N__6679),
            .I(N__6631));
    InMux I__953 (
            .O(N__6678),
            .I(N__6631));
    InMux I__952 (
            .O(N__6675),
            .I(N__6628));
    LocalMux I__951 (
            .O(N__6672),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    Odrv4 I__950 (
            .O(N__6669),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    Odrv4 I__949 (
            .O(N__6666),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    LocalMux I__948 (
            .O(N__6659),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    LocalMux I__947 (
            .O(N__6654),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    Odrv4 I__946 (
            .O(N__6649),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    LocalMux I__945 (
            .O(N__6644),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    LocalMux I__944 (
            .O(N__6639),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    Odrv4 I__943 (
            .O(N__6636),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    LocalMux I__942 (
            .O(N__6631),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    LocalMux I__941 (
            .O(N__6628),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    CascadeMux I__940 (
            .O(N__6605),
            .I(\DUT.uart_inst0.N_8_0_cascade_ ));
    InMux I__939 (
            .O(N__6602),
            .I(N__6599));
    LocalMux I__938 (
            .O(N__6599),
            .I(\DUT.uart_inst0.m10_0_1 ));
    InMux I__937 (
            .O(N__6596),
            .I(N__6593));
    LocalMux I__936 (
            .O(N__6593),
            .I(N__6590));
    Odrv4 I__935 (
            .O(N__6590),
            .I(\DUT.uart_inst0.m11_0 ));
    InMux I__934 (
            .O(N__6587),
            .I(N__6584));
    LocalMux I__933 (
            .O(N__6584),
            .I(N__6581));
    Odrv4 I__932 (
            .O(N__6581),
            .I(\DUT.uart_inst0.N_15_mux ));
    CascadeMux I__931 (
            .O(N__6578),
            .I(\DUT.uart_inst0.N_11_0_cascade_ ));
    CascadeMux I__930 (
            .O(N__6575),
            .I(N__6572));
    InMux I__929 (
            .O(N__6572),
            .I(N__6569));
    LocalMux I__928 (
            .O(N__6569),
            .I(\DUT.uart_inst0.N_81_mux_i_i_a5_1_3 ));
    CascadeMux I__927 (
            .O(N__6566),
            .I(N__6555));
    InMux I__926 (
            .O(N__6565),
            .I(N__6550));
    InMux I__925 (
            .O(N__6564),
            .I(N__6547));
    InMux I__924 (
            .O(N__6563),
            .I(N__6542));
    InMux I__923 (
            .O(N__6562),
            .I(N__6542));
    InMux I__922 (
            .O(N__6561),
            .I(N__6537));
    InMux I__921 (
            .O(N__6560),
            .I(N__6537));
    InMux I__920 (
            .O(N__6559),
            .I(N__6532));
    InMux I__919 (
            .O(N__6558),
            .I(N__6532));
    InMux I__918 (
            .O(N__6555),
            .I(N__6525));
    InMux I__917 (
            .O(N__6554),
            .I(N__6525));
    InMux I__916 (
            .O(N__6553),
            .I(N__6525));
    LocalMux I__915 (
            .O(N__6550),
            .I(N__6522));
    LocalMux I__914 (
            .O(N__6547),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_3 ));
    LocalMux I__913 (
            .O(N__6542),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_3 ));
    LocalMux I__912 (
            .O(N__6537),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_3 ));
    LocalMux I__911 (
            .O(N__6532),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_3 ));
    LocalMux I__910 (
            .O(N__6525),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_3 ));
    Odrv4 I__909 (
            .O(N__6522),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_3 ));
    CascadeMux I__908 (
            .O(N__6509),
            .I(\DUT.uart_inst0.N_300_cascade_ ));
    CascadeMux I__907 (
            .O(N__6506),
            .I(\DUT.uart_inst0.G_16_i_a3_3_cascade_ ));
    InMux I__906 (
            .O(N__6503),
            .I(N__6500));
    LocalMux I__905 (
            .O(N__6500),
            .I(N__6497));
    Odrv12 I__904 (
            .O(N__6497),
            .I(\DUT.uart_inst0.G_16_i_a3_4 ));
    InMux I__903 (
            .O(N__6494),
            .I(N__6488));
    InMux I__902 (
            .O(N__6493),
            .I(N__6484));
    CascadeMux I__901 (
            .O(N__6492),
            .I(N__6474));
    InMux I__900 (
            .O(N__6491),
            .I(N__6471));
    LocalMux I__899 (
            .O(N__6488),
            .I(N__6468));
    InMux I__898 (
            .O(N__6487),
            .I(N__6465));
    LocalMux I__897 (
            .O(N__6484),
            .I(N__6462));
    InMux I__896 (
            .O(N__6483),
            .I(N__6455));
    InMux I__895 (
            .O(N__6482),
            .I(N__6455));
    InMux I__894 (
            .O(N__6481),
            .I(N__6455));
    InMux I__893 (
            .O(N__6480),
            .I(N__6446));
    InMux I__892 (
            .O(N__6479),
            .I(N__6446));
    InMux I__891 (
            .O(N__6478),
            .I(N__6446));
    InMux I__890 (
            .O(N__6477),
            .I(N__6446));
    InMux I__889 (
            .O(N__6474),
            .I(N__6443));
    LocalMux I__888 (
            .O(N__6471),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_1 ));
    Odrv4 I__887 (
            .O(N__6468),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_1 ));
    LocalMux I__886 (
            .O(N__6465),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_1 ));
    Odrv4 I__885 (
            .O(N__6462),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_1 ));
    LocalMux I__884 (
            .O(N__6455),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_1 ));
    LocalMux I__883 (
            .O(N__6446),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_1 ));
    LocalMux I__882 (
            .O(N__6443),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_1 ));
    InMux I__881 (
            .O(N__6428),
            .I(N__6421));
    InMux I__880 (
            .O(N__6427),
            .I(N__6416));
    CascadeMux I__879 (
            .O(N__6426),
            .I(N__6413));
    InMux I__878 (
            .O(N__6425),
            .I(N__6409));
    CascadeMux I__877 (
            .O(N__6424),
            .I(N__6406));
    LocalMux I__876 (
            .O(N__6421),
            .I(N__6401));
    CascadeMux I__875 (
            .O(N__6420),
            .I(N__6397));
    InMux I__874 (
            .O(N__6419),
            .I(N__6393));
    LocalMux I__873 (
            .O(N__6416),
            .I(N__6390));
    InMux I__872 (
            .O(N__6413),
            .I(N__6385));
    InMux I__871 (
            .O(N__6412),
            .I(N__6385));
    LocalMux I__870 (
            .O(N__6409),
            .I(N__6382));
    InMux I__869 (
            .O(N__6406),
            .I(N__6379));
    InMux I__868 (
            .O(N__6405),
            .I(N__6374));
    InMux I__867 (
            .O(N__6404),
            .I(N__6374));
    Span4Mux_h I__866 (
            .O(N__6401),
            .I(N__6371));
    InMux I__865 (
            .O(N__6400),
            .I(N__6368));
    InMux I__864 (
            .O(N__6397),
            .I(N__6363));
    InMux I__863 (
            .O(N__6396),
            .I(N__6363));
    LocalMux I__862 (
            .O(N__6393),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_5 ));
    Odrv4 I__861 (
            .O(N__6390),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_5 ));
    LocalMux I__860 (
            .O(N__6385),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_5 ));
    Odrv4 I__859 (
            .O(N__6382),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_5 ));
    LocalMux I__858 (
            .O(N__6379),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_5 ));
    LocalMux I__857 (
            .O(N__6374),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_5 ));
    Odrv4 I__856 (
            .O(N__6371),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_5 ));
    LocalMux I__855 (
            .O(N__6368),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_5 ));
    LocalMux I__854 (
            .O(N__6363),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_5 ));
    InMux I__853 (
            .O(N__6344),
            .I(N__6341));
    LocalMux I__852 (
            .O(N__6341),
            .I(N__6338));
    Odrv12 I__851 (
            .O(N__6338),
            .I(\DUT.uart_inst0.N_11_2 ));
    CascadeMux I__850 (
            .O(N__6335),
            .I(N__6329));
    InMux I__849 (
            .O(N__6334),
            .I(N__6326));
    CascadeMux I__848 (
            .O(N__6333),
            .I(N__6322));
    CascadeMux I__847 (
            .O(N__6332),
            .I(N__6317));
    InMux I__846 (
            .O(N__6329),
            .I(N__6311));
    LocalMux I__845 (
            .O(N__6326),
            .I(N__6308));
    InMux I__844 (
            .O(N__6325),
            .I(N__6305));
    InMux I__843 (
            .O(N__6322),
            .I(N__6302));
    InMux I__842 (
            .O(N__6321),
            .I(N__6297));
    InMux I__841 (
            .O(N__6320),
            .I(N__6297));
    InMux I__840 (
            .O(N__6317),
            .I(N__6294));
    InMux I__839 (
            .O(N__6316),
            .I(N__6287));
    InMux I__838 (
            .O(N__6315),
            .I(N__6287));
    InMux I__837 (
            .O(N__6314),
            .I(N__6287));
    LocalMux I__836 (
            .O(N__6311),
            .I(N__6284));
    Odrv4 I__835 (
            .O(N__6308),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_2 ));
    LocalMux I__834 (
            .O(N__6305),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_2 ));
    LocalMux I__833 (
            .O(N__6302),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_2 ));
    LocalMux I__832 (
            .O(N__6297),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_2 ));
    LocalMux I__831 (
            .O(N__6294),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_2 ));
    LocalMux I__830 (
            .O(N__6287),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_2 ));
    Odrv4 I__829 (
            .O(N__6284),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_2 ));
    InMux I__828 (
            .O(N__6269),
            .I(N__6266));
    LocalMux I__827 (
            .O(N__6266),
            .I(\DUT.uart_inst0.G_16_i_a3_0_3 ));
    CascadeMux I__826 (
            .O(N__6263),
            .I(N__6260));
    InMux I__825 (
            .O(N__6260),
            .I(N__6257));
    LocalMux I__824 (
            .O(N__6257),
            .I(\DUT.uart_inst0.g1_1 ));
    CascadeMux I__823 (
            .O(N__6254),
            .I(N__6245));
    CascadeMux I__822 (
            .O(N__6253),
            .I(N__6239));
    CascadeMux I__821 (
            .O(N__6252),
            .I(N__6235));
    InMux I__820 (
            .O(N__6251),
            .I(N__6231));
    InMux I__819 (
            .O(N__6250),
            .I(N__6228));
    InMux I__818 (
            .O(N__6249),
            .I(N__6225));
    InMux I__817 (
            .O(N__6248),
            .I(N__6220));
    InMux I__816 (
            .O(N__6245),
            .I(N__6220));
    InMux I__815 (
            .O(N__6244),
            .I(N__6213));
    InMux I__814 (
            .O(N__6243),
            .I(N__6213));
    InMux I__813 (
            .O(N__6242),
            .I(N__6213));
    InMux I__812 (
            .O(N__6239),
            .I(N__6208));
    InMux I__811 (
            .O(N__6238),
            .I(N__6208));
    InMux I__810 (
            .O(N__6235),
            .I(N__6205));
    InMux I__809 (
            .O(N__6234),
            .I(N__6202));
    LocalMux I__808 (
            .O(N__6231),
            .I(N__6197));
    LocalMux I__807 (
            .O(N__6228),
            .I(N__6197));
    LocalMux I__806 (
            .O(N__6225),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_1 ));
    LocalMux I__805 (
            .O(N__6220),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_1 ));
    LocalMux I__804 (
            .O(N__6213),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_1 ));
    LocalMux I__803 (
            .O(N__6208),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_1 ));
    LocalMux I__802 (
            .O(N__6205),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_1 ));
    LocalMux I__801 (
            .O(N__6202),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_1 ));
    Odrv4 I__800 (
            .O(N__6197),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_1 ));
    InMux I__799 (
            .O(N__6182),
            .I(N__6179));
    LocalMux I__798 (
            .O(N__6179),
            .I(\DUT.uart_inst0.N_81_mux_i_i_a5_1_5_0 ));
    InMux I__797 (
            .O(N__6176),
            .I(N__6173));
    LocalMux I__796 (
            .O(N__6173),
            .I(\DUT.uart_inst0.rx_countdown_RNO_2Z0Z_2 ));
    CascadeMux I__795 (
            .O(N__6170),
            .I(\DUT.uart_inst0.G_21_0_1_0_cascade_ ));
    InMux I__794 (
            .O(N__6167),
            .I(N__6164));
    LocalMux I__793 (
            .O(N__6164),
            .I(\DUT.uart_inst0.G_9_i_o4_0 ));
    InMux I__792 (
            .O(N__6161),
            .I(N__6158));
    LocalMux I__791 (
            .O(N__6158),
            .I(\DUT.uart_inst0.g0_0_3 ));
    CascadeMux I__790 (
            .O(N__6155),
            .I(\DUT.uart_inst0.G_16_i_a3_0_2_cascade_ ));
    CascadeMux I__789 (
            .O(N__6152),
            .I(\DUT.uart_inst0.N_45_cascade_ ));
    InMux I__788 (
            .O(N__6149),
            .I(N__6146));
    LocalMux I__787 (
            .O(N__6146),
            .I(\DUT.uart_inst0.N_55 ));
    InMux I__786 (
            .O(N__6143),
            .I(N__6137));
    CascadeMux I__785 (
            .O(N__6142),
            .I(N__6133));
    CascadeMux I__784 (
            .O(N__6141),
            .I(N__6127));
    InMux I__783 (
            .O(N__6140),
            .I(N__6121));
    LocalMux I__782 (
            .O(N__6137),
            .I(N__6118));
    InMux I__781 (
            .O(N__6136),
            .I(N__6113));
    InMux I__780 (
            .O(N__6133),
            .I(N__6113));
    InMux I__779 (
            .O(N__6132),
            .I(N__6108));
    InMux I__778 (
            .O(N__6131),
            .I(N__6108));
    InMux I__777 (
            .O(N__6130),
            .I(N__6103));
    InMux I__776 (
            .O(N__6127),
            .I(N__6103));
    InMux I__775 (
            .O(N__6126),
            .I(N__6100));
    InMux I__774 (
            .O(N__6125),
            .I(N__6095));
    InMux I__773 (
            .O(N__6124),
            .I(N__6095));
    LocalMux I__772 (
            .O(N__6121),
            .I(N__6092));
    Odrv4 I__771 (
            .O(N__6118),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_4 ));
    LocalMux I__770 (
            .O(N__6113),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_4 ));
    LocalMux I__769 (
            .O(N__6108),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_4 ));
    LocalMux I__768 (
            .O(N__6103),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_4 ));
    LocalMux I__767 (
            .O(N__6100),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_4 ));
    LocalMux I__766 (
            .O(N__6095),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_4 ));
    Odrv4 I__765 (
            .O(N__6092),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_4 ));
    InMux I__764 (
            .O(N__6077),
            .I(N__6074));
    LocalMux I__763 (
            .O(N__6074),
            .I(\DUT.uart_inst0.N_10 ));
    CascadeMux I__762 (
            .O(N__6071),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0_cascade_ ));
    InMux I__761 (
            .O(N__6068),
            .I(N__6065));
    LocalMux I__760 (
            .O(N__6065),
            .I(\DUT.uart_inst0.G_21_0_1 ));
    InMux I__759 (
            .O(N__6062),
            .I(N__6059));
    LocalMux I__758 (
            .O(N__6059),
            .I(N__6055));
    InMux I__757 (
            .O(N__6058),
            .I(N__6052));
    Odrv4 I__756 (
            .O(N__6055),
            .I(\DUT.uart_inst0.recv_stateZ0Z_4 ));
    LocalMux I__755 (
            .O(N__6052),
            .I(\DUT.uart_inst0.recv_stateZ0Z_4 ));
    CascadeMux I__754 (
            .O(N__6047),
            .I(N__6043));
    InMux I__753 (
            .O(N__6046),
            .I(N__6039));
    InMux I__752 (
            .O(N__6043),
            .I(N__6034));
    InMux I__751 (
            .O(N__6042),
            .I(N__6034));
    LocalMux I__750 (
            .O(N__6039),
            .I(\DUT.uart_inst0.N_45 ));
    LocalMux I__749 (
            .O(N__6034),
            .I(\DUT.uart_inst0.N_45 ));
    InMux I__748 (
            .O(N__6029),
            .I(N__6026));
    LocalMux I__747 (
            .O(N__6026),
            .I(N__6023));
    Span4Mux_h I__746 (
            .O(N__6023),
            .I(N__6020));
    Odrv4 I__745 (
            .O(N__6020),
            .I(\DUT.uart_inst0.recv_state_ns_0_0_0 ));
    CascadeMux I__744 (
            .O(N__6017),
            .I(N__6014));
    InMux I__743 (
            .O(N__6014),
            .I(N__6011));
    LocalMux I__742 (
            .O(N__6011),
            .I(N__6008));
    Odrv4 I__741 (
            .O(N__6008),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_2 ));
    InMux I__740 (
            .O(N__6005),
            .I(N__6002));
    LocalMux I__739 (
            .O(N__6002),
            .I(N__5999));
    Odrv4 I__738 (
            .O(N__5999),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_3 ));
    CascadeMux I__737 (
            .O(N__5996),
            .I(N__5993));
    InMux I__736 (
            .O(N__5993),
            .I(N__5990));
    LocalMux I__735 (
            .O(N__5990),
            .I(N__5987));
    Odrv4 I__734 (
            .O(N__5987),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_4 ));
    CascadeMux I__733 (
            .O(N__5984),
            .I(N__5981));
    InMux I__732 (
            .O(N__5981),
            .I(N__5978));
    LocalMux I__731 (
            .O(N__5978),
            .I(N__5975));
    Odrv4 I__730 (
            .O(N__5975),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_5 ));
    CascadeMux I__729 (
            .O(N__5972),
            .I(N__5969));
    InMux I__728 (
            .O(N__5969),
            .I(N__5966));
    LocalMux I__727 (
            .O(N__5966),
            .I(N__5963));
    Odrv4 I__726 (
            .O(N__5963),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_6 ));
    InMux I__725 (
            .O(N__5960),
            .I(N__5957));
    LocalMux I__724 (
            .O(N__5957),
            .I(\DUT.uart_inst0.N_81_mux_i_i_a5_1_4 ));
    InMux I__723 (
            .O(N__5954),
            .I(N__5951));
    LocalMux I__722 (
            .O(N__5951),
            .I(\DUT.uart_inst0.N_13_0 ));
    InMux I__721 (
            .O(N__5948),
            .I(N__5945));
    LocalMux I__720 (
            .O(N__5945),
            .I(N__5942));
    Odrv4 I__719 (
            .O(N__5942),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_3 ));
    CascadeMux I__718 (
            .O(N__5939),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ));
    CascadeMux I__717 (
            .O(N__5936),
            .I(N__5933));
    InMux I__716 (
            .O(N__5933),
            .I(N__5930));
    LocalMux I__715 (
            .O(N__5930),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_0 ));
    InMux I__714 (
            .O(N__5927),
            .I(N__5924));
    LocalMux I__713 (
            .O(N__5924),
            .I(N__5921));
    Span4Mux_v I__712 (
            .O(N__5921),
            .I(N__5918));
    Odrv4 I__711 (
            .O(N__5918),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_0 ));
    CascadeMux I__710 (
            .O(N__5915),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ));
    InMux I__709 (
            .O(N__5912),
            .I(N__5909));
    LocalMux I__708 (
            .O(N__5909),
            .I(N__5906));
    Span4Mux_h I__707 (
            .O(N__5906),
            .I(N__5903));
    Odrv4 I__706 (
            .O(N__5903),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_7 ));
    InMux I__705 (
            .O(N__5900),
            .I(N__5897));
    LocalMux I__704 (
            .O(N__5897),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_1 ));
    InMux I__703 (
            .O(N__5894),
            .I(N__5891));
    LocalMux I__702 (
            .O(N__5891),
            .I(N__5888));
    Span4Mux_h I__701 (
            .O(N__5888),
            .I(N__5885));
    Odrv4 I__700 (
            .O(N__5885),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_2 ));
    InMux I__699 (
            .O(N__5882),
            .I(N__5879));
    LocalMux I__698 (
            .O(N__5879),
            .I(N__5876));
    Odrv4 I__697 (
            .O(N__5876),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2 ));
    InMux I__696 (
            .O(N__5873),
            .I(N__5870));
    LocalMux I__695 (
            .O(N__5870),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_0 ));
    CascadeMux I__694 (
            .O(N__5867),
            .I(N__5864));
    InMux I__693 (
            .O(N__5864),
            .I(N__5861));
    LocalMux I__692 (
            .O(N__5861),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_1 ));
    InMux I__691 (
            .O(N__5858),
            .I(N__5850));
    InMux I__690 (
            .O(N__5857),
            .I(N__5850));
    InMux I__689 (
            .O(N__5856),
            .I(N__5845));
    InMux I__688 (
            .O(N__5855),
            .I(N__5845));
    LocalMux I__687 (
            .O(N__5850),
            .I(\DUT.fifo_rx_inst.rWritePtr16 ));
    LocalMux I__686 (
            .O(N__5845),
            .I(\DUT.fifo_rx_inst.rWritePtr16 ));
    CascadeMux I__685 (
            .O(N__5840),
            .I(N__5836));
    InMux I__684 (
            .O(N__5839),
            .I(N__5826));
    InMux I__683 (
            .O(N__5836),
            .I(N__5826));
    InMux I__682 (
            .O(N__5835),
            .I(N__5826));
    CascadeMux I__681 (
            .O(N__5834),
            .I(N__5823));
    CascadeMux I__680 (
            .O(N__5833),
            .I(N__5819));
    LocalMux I__679 (
            .O(N__5826),
            .I(N__5816));
    InMux I__678 (
            .O(N__5823),
            .I(N__5809));
    InMux I__677 (
            .O(N__5822),
            .I(N__5809));
    InMux I__676 (
            .O(N__5819),
            .I(N__5809));
    Odrv4 I__675 (
            .O(N__5816),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_0 ));
    LocalMux I__674 (
            .O(N__5809),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_0 ));
    InMux I__673 (
            .O(N__5804),
            .I(N__5793));
    InMux I__672 (
            .O(N__5803),
            .I(N__5793));
    InMux I__671 (
            .O(N__5802),
            .I(N__5793));
    InMux I__670 (
            .O(N__5801),
            .I(N__5788));
    InMux I__669 (
            .O(N__5800),
            .I(N__5788));
    LocalMux I__668 (
            .O(N__5793),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_1 ));
    LocalMux I__667 (
            .O(N__5788),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_1 ));
    InMux I__666 (
            .O(N__5783),
            .I(N__5780));
    LocalMux I__665 (
            .O(N__5780),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_2 ));
    CascadeMux I__664 (
            .O(N__5777),
            .I(N__5774));
    InMux I__663 (
            .O(N__5774),
            .I(N__5771));
    LocalMux I__662 (
            .O(N__5771),
            .I(N__5768));
    Odrv4 I__661 (
            .O(N__5768),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_6 ));
    InMux I__660 (
            .O(N__5765),
            .I(N__5762));
    LocalMux I__659 (
            .O(N__5762),
            .I(N__5759));
    Odrv4 I__658 (
            .O(N__5759),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_4 ));
    InMux I__657 (
            .O(N__5756),
            .I(N__5753));
    LocalMux I__656 (
            .O(N__5753),
            .I(N__5750));
    Odrv4 I__655 (
            .O(N__5750),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_4 ));
    CascadeMux I__654 (
            .O(N__5747),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4_cascade_ ));
    InMux I__653 (
            .O(N__5744),
            .I(N__5741));
    LocalMux I__652 (
            .O(N__5741),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_5 ));
    CascadeMux I__651 (
            .O(N__5738),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ));
    InMux I__650 (
            .O(N__5735),
            .I(N__5732));
    LocalMux I__649 (
            .O(N__5732),
            .I(N__5729));
    Odrv4 I__648 (
            .O(N__5729),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_5 ));
    InMux I__647 (
            .O(N__5726),
            .I(N__5723));
    LocalMux I__646 (
            .O(N__5723),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_6 ));
    InMux I__645 (
            .O(N__5720),
            .I(N__5717));
    LocalMux I__644 (
            .O(N__5717),
            .I(N__5714));
    Odrv4 I__643 (
            .O(N__5714),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6 ));
    InMux I__642 (
            .O(N__5711),
            .I(N__5708));
    LocalMux I__641 (
            .O(N__5708),
            .I(N__5705));
    Odrv4 I__640 (
            .O(N__5705),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_3 ));
    CascadeMux I__639 (
            .O(N__5702),
            .I(\DUT.fifo_rx_inst.rFifoData_awe3_cascade_ ));
    CascadeMux I__638 (
            .O(N__5699),
            .I(\DUT.fifo_rx_inst.un1_i11_i_cascade_ ));
    InMux I__637 (
            .O(N__5696),
            .I(N__5693));
    LocalMux I__636 (
            .O(N__5693),
            .I(\DUT.fifo_rx_inst.un1_rFifoCount_1_axb_2 ));
    InMux I__635 (
            .O(N__5690),
            .I(N__5687));
    LocalMux I__634 (
            .O(N__5687),
            .I(\DUT.fifo_rx_inst.un1_i11_i ));
    CascadeMux I__633 (
            .O(N__5684),
            .I(N__5681));
    InMux I__632 (
            .O(N__5681),
            .I(N__5678));
    LocalMux I__631 (
            .O(N__5678),
            .I(\DUT.fifo_rx_inst.rFifoCount_RNIK3G92Z0Z_1 ));
    CascadeMux I__630 (
            .O(N__5675),
            .I(\DUT.fifo_rx_inst.rWritePtr16_cascade_ ));
    CascadeMux I__629 (
            .O(N__5672),
            .I(\DUT.uart_inst0.g0_0_i_a3_3_cascade_ ));
    InMux I__628 (
            .O(N__5669),
            .I(N__5666));
    LocalMux I__627 (
            .O(N__5666),
            .I(\DUT.uart_inst0.g0_0_i_a3_4 ));
    InMux I__626 (
            .O(N__5663),
            .I(N__5660));
    LocalMux I__625 (
            .O(N__5660),
            .I(N__5654));
    InMux I__624 (
            .O(N__5659),
            .I(N__5651));
    InMux I__623 (
            .O(N__5658),
            .I(N__5646));
    InMux I__622 (
            .O(N__5657),
            .I(N__5646));
    Span4Mux_h I__621 (
            .O(N__5654),
            .I(N__5639));
    LocalMux I__620 (
            .O(N__5651),
            .I(N__5634));
    LocalMux I__619 (
            .O(N__5646),
            .I(N__5634));
    InMux I__618 (
            .O(N__5645),
            .I(N__5629));
    InMux I__617 (
            .O(N__5644),
            .I(N__5629));
    InMux I__616 (
            .O(N__5643),
            .I(N__5626));
    InMux I__615 (
            .O(N__5642),
            .I(N__5623));
    Odrv4 I__614 (
            .O(N__5639),
            .I(\DUT.uart_inst0.recv_stateZ0Z_2 ));
    Odrv12 I__613 (
            .O(N__5634),
            .I(\DUT.uart_inst0.recv_stateZ0Z_2 ));
    LocalMux I__612 (
            .O(N__5629),
            .I(\DUT.uart_inst0.recv_stateZ0Z_2 ));
    LocalMux I__611 (
            .O(N__5626),
            .I(\DUT.uart_inst0.recv_stateZ0Z_2 ));
    LocalMux I__610 (
            .O(N__5623),
            .I(\DUT.uart_inst0.recv_stateZ0Z_2 ));
    IoInMux I__609 (
            .O(N__5612),
            .I(N__5609));
    LocalMux I__608 (
            .O(N__5609),
            .I(N__5606));
    Span4Mux_s2_v I__607 (
            .O(N__5606),
            .I(N__5603));
    Span4Mux_h I__606 (
            .O(N__5603),
            .I(N__5600));
    Span4Mux_v I__605 (
            .O(N__5600),
            .I(N__5597));
    Span4Mux_v I__604 (
            .O(N__5597),
            .I(N__5594));
    Odrv4 I__603 (
            .O(N__5594),
            .I(wPllLocked_i));
    InMux I__602 (
            .O(N__5591),
            .I(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0 ));
    InMux I__601 (
            .O(N__5588),
            .I(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1 ));
    InMux I__600 (
            .O(N__5585),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_4_s1 ));
    InMux I__599 (
            .O(N__5582),
            .I(N__5579));
    LocalMux I__598 (
            .O(N__5579),
            .I(\DUT.uart_inst0.m9_3 ));
    InMux I__597 (
            .O(N__5576),
            .I(N__5573));
    LocalMux I__596 (
            .O(N__5573),
            .I(\DUT.uart_inst0.m9_4 ));
    InMux I__595 (
            .O(N__5570),
            .I(N__5567));
    LocalMux I__594 (
            .O(N__5567),
            .I(\DUT.uart_inst0.N_8 ));
    CascadeMux I__593 (
            .O(N__5564),
            .I(N__5561));
    InMux I__592 (
            .O(N__5561),
            .I(N__5558));
    LocalMux I__591 (
            .O(N__5558),
            .I(\DUT.uart_inst0.N_81_mux_i_i_0_0 ));
    InMux I__590 (
            .O(N__5555),
            .I(N__5552));
    LocalMux I__589 (
            .O(N__5552),
            .I(\DUT.uart_inst0.N_81_mux_i_i_a5_0_5_0 ));
    CascadeMux I__588 (
            .O(N__5549),
            .I(\DUT.uart_inst0.m4_3_cascade_ ));
    CascadeMux I__587 (
            .O(N__5546),
            .I(N__5543));
    InMux I__586 (
            .O(N__5543),
            .I(N__5540));
    LocalMux I__585 (
            .O(N__5540),
            .I(\DUT.uart_inst0.N_18_mux ));
    CascadeMux I__584 (
            .O(N__5537),
            .I(\DUT.uart_inst0.N_297_cascade_ ));
    InMux I__583 (
            .O(N__5534),
            .I(N__5523));
    InMux I__582 (
            .O(N__5533),
            .I(N__5523));
    InMux I__581 (
            .O(N__5532),
            .I(N__5517));
    InMux I__580 (
            .O(N__5531),
            .I(N__5517));
    InMux I__579 (
            .O(N__5530),
            .I(N__5512));
    InMux I__578 (
            .O(N__5529),
            .I(N__5512));
    CascadeMux I__577 (
            .O(N__5528),
            .I(N__5508));
    LocalMux I__576 (
            .O(N__5523),
            .I(N__5503));
    InMux I__575 (
            .O(N__5522),
            .I(N__5500));
    LocalMux I__574 (
            .O(N__5517),
            .I(N__5495));
    LocalMux I__573 (
            .O(N__5512),
            .I(N__5495));
    InMux I__572 (
            .O(N__5511),
            .I(N__5492));
    InMux I__571 (
            .O(N__5508),
            .I(N__5489));
    InMux I__570 (
            .O(N__5507),
            .I(N__5486));
    InMux I__569 (
            .O(N__5506),
            .I(N__5483));
    Odrv4 I__568 (
            .O(N__5503),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    LocalMux I__567 (
            .O(N__5500),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    Odrv4 I__566 (
            .O(N__5495),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    LocalMux I__565 (
            .O(N__5492),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    LocalMux I__564 (
            .O(N__5489),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    LocalMux I__563 (
            .O(N__5486),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    LocalMux I__562 (
            .O(N__5483),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    InMux I__561 (
            .O(N__5468),
            .I(N__5465));
    LocalMux I__560 (
            .O(N__5465),
            .I(\DUT.uart_inst0.N_15_3 ));
    InMux I__559 (
            .O(N__5462),
            .I(N__5459));
    LocalMux I__558 (
            .O(N__5459),
            .I(N__5456));
    Odrv4 I__557 (
            .O(N__5456),
            .I(\DUT.uart_inst0.N_81_mux_i_i_a5_0_4 ));
    InMux I__556 (
            .O(N__5453),
            .I(N__5450));
    LocalMux I__555 (
            .O(N__5450),
            .I(\DUT.uart_inst0.N_81_mux_i_i_0 ));
    CascadeMux I__554 (
            .O(N__5447),
            .I(\DUT.uart_inst0.N_81_mux_i_i_a5_0_5_cascade_ ));
    InMux I__553 (
            .O(N__5444),
            .I(N__5441));
    LocalMux I__552 (
            .O(N__5441),
            .I(\DUT.uart_inst0.N_81_mux_i_i_a5_1_5 ));
    InMux I__551 (
            .O(N__5438),
            .I(N__5435));
    LocalMux I__550 (
            .O(N__5435),
            .I(N__5432));
    Odrv4 I__549 (
            .O(N__5432),
            .I(\DUT.uart_inst0.m8_e_2 ));
    InMux I__548 (
            .O(N__5429),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_0_s1 ));
    InMux I__547 (
            .O(N__5426),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_1_s1 ));
    InMux I__546 (
            .O(N__5423),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_2_s1 ));
    InMux I__545 (
            .O(N__5420),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_3_s1 ));
    InMux I__544 (
            .O(N__5417),
            .I(N__5414));
    LocalMux I__543 (
            .O(N__5414),
            .I(N__5411));
    Odrv4 I__542 (
            .O(N__5411),
            .I(\DUT.uart_inst0.m8_e_3 ));
    InMux I__541 (
            .O(N__5408),
            .I(N__5398));
    CascadeMux I__540 (
            .O(N__5407),
            .I(N__5395));
    InMux I__539 (
            .O(N__5406),
            .I(N__5384));
    InMux I__538 (
            .O(N__5405),
            .I(N__5384));
    InMux I__537 (
            .O(N__5404),
            .I(N__5384));
    InMux I__536 (
            .O(N__5403),
            .I(N__5384));
    InMux I__535 (
            .O(N__5402),
            .I(N__5384));
    InMux I__534 (
            .O(N__5401),
            .I(N__5381));
    LocalMux I__533 (
            .O(N__5398),
            .I(N__5378));
    InMux I__532 (
            .O(N__5395),
            .I(N__5375));
    LocalMux I__531 (
            .O(N__5384),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_1 ));
    LocalMux I__530 (
            .O(N__5381),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_1 ));
    Odrv12 I__529 (
            .O(N__5378),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_1 ));
    LocalMux I__528 (
            .O(N__5375),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_1 ));
    InMux I__527 (
            .O(N__5366),
            .I(N__5363));
    LocalMux I__526 (
            .O(N__5363),
            .I(N__5360));
    Odrv4 I__525 (
            .O(N__5360),
            .I(\DUT.uart_inst0.g0_i_a3_6 ));
    InMux I__524 (
            .O(N__5357),
            .I(N__5354));
    LocalMux I__523 (
            .O(N__5354),
            .I(N__5351));
    Odrv4 I__522 (
            .O(N__5351),
            .I(\DUT.uart_inst0.recv_state_ns_0_i_a2_0_0_3 ));
    InMux I__521 (
            .O(N__5348),
            .I(N__5339));
    InMux I__520 (
            .O(N__5347),
            .I(N__5339));
    InMux I__519 (
            .O(N__5346),
            .I(N__5339));
    LocalMux I__518 (
            .O(N__5339),
            .I(\DUT.uart_inst0.recv_stateZ0Z_3 ));
    InMux I__517 (
            .O(N__5336),
            .I(N__5333));
    LocalMux I__516 (
            .O(N__5333),
            .I(\DUT.uart_inst0.g0_0_0 ));
    InMux I__515 (
            .O(N__5330),
            .I(N__5327));
    LocalMux I__514 (
            .O(N__5327),
            .I(\DUT.uart_inst0.g0_0_1 ));
    CascadeMux I__513 (
            .O(N__5324),
            .I(\DUT.uart_inst0.N_81_mux_i_i_a5_0_4_0_cascade_ ));
    InMux I__512 (
            .O(N__5321),
            .I(N__5318));
    LocalMux I__511 (
            .O(N__5318),
            .I(\DUT.uart_inst0.N_35_0 ));
    CascadeMux I__510 (
            .O(N__5315),
            .I(\DUT.uart_inst0.g0_0_2_cascade_ ));
    InMux I__509 (
            .O(N__5312),
            .I(N__5307));
    InMux I__508 (
            .O(N__5311),
            .I(N__5303));
    InMux I__507 (
            .O(N__5310),
            .I(N__5300));
    LocalMux I__506 (
            .O(N__5307),
            .I(N__5296));
    InMux I__505 (
            .O(N__5306),
            .I(N__5292));
    LocalMux I__504 (
            .O(N__5303),
            .I(N__5287));
    LocalMux I__503 (
            .O(N__5300),
            .I(N__5287));
    InMux I__502 (
            .O(N__5299),
            .I(N__5284));
    Span4Mux_h I__501 (
            .O(N__5296),
            .I(N__5281));
    InMux I__500 (
            .O(N__5295),
            .I(N__5278));
    LocalMux I__499 (
            .O(N__5292),
            .I(N__5273));
    Span4Mux_v I__498 (
            .O(N__5287),
            .I(N__5273));
    LocalMux I__497 (
            .O(N__5284),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_2 ));
    Odrv4 I__496 (
            .O(N__5281),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_2 ));
    LocalMux I__495 (
            .O(N__5278),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_2 ));
    Odrv4 I__494 (
            .O(N__5273),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_2 ));
    InMux I__493 (
            .O(N__5264),
            .I(N__5261));
    LocalMux I__492 (
            .O(N__5261),
            .I(\DUT.uart_inst0.g0_i_a3_0_6 ));
    CascadeMux I__491 (
            .O(N__5258),
            .I(\DUT.uart_inst0.g0_i_a3_0_7_cascade_ ));
    CascadeMux I__490 (
            .O(N__5255),
            .I(\DUT.uart_inst0.N_6_0_cascade_ ));
    CascadeMux I__489 (
            .O(N__5252),
            .I(N__5249));
    InMux I__488 (
            .O(N__5249),
            .I(N__5246));
    LocalMux I__487 (
            .O(N__5246),
            .I(N__5243));
    Odrv12 I__486 (
            .O(N__5243),
            .I(\DUT.uart_inst0.N_40 ));
    CascadeMux I__485 (
            .O(N__5240),
            .I(N__5237));
    InMux I__484 (
            .O(N__5237),
            .I(N__5231));
    InMux I__483 (
            .O(N__5236),
            .I(N__5226));
    InMux I__482 (
            .O(N__5235),
            .I(N__5226));
    InMux I__481 (
            .O(N__5234),
            .I(N__5223));
    LocalMux I__480 (
            .O(N__5231),
            .I(N__5220));
    LocalMux I__479 (
            .O(N__5226),
            .I(N__5217));
    LocalMux I__478 (
            .O(N__5223),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_3 ));
    Odrv4 I__477 (
            .O(N__5220),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_3 ));
    Odrv4 I__476 (
            .O(N__5217),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_3 ));
    CascadeMux I__475 (
            .O(N__5210),
            .I(N__5205));
    InMux I__474 (
            .O(N__5209),
            .I(N__5200));
    InMux I__473 (
            .O(N__5208),
            .I(N__5197));
    InMux I__472 (
            .O(N__5205),
            .I(N__5192));
    InMux I__471 (
            .O(N__5204),
            .I(N__5192));
    CascadeMux I__470 (
            .O(N__5203),
            .I(N__5189));
    LocalMux I__469 (
            .O(N__5200),
            .I(N__5180));
    LocalMux I__468 (
            .O(N__5197),
            .I(N__5180));
    LocalMux I__467 (
            .O(N__5192),
            .I(N__5180));
    InMux I__466 (
            .O(N__5189),
            .I(N__5177));
    InMux I__465 (
            .O(N__5188),
            .I(N__5174));
    InMux I__464 (
            .O(N__5187),
            .I(N__5171));
    Span4Mux_v I__463 (
            .O(N__5180),
            .I(N__5166));
    LocalMux I__462 (
            .O(N__5177),
            .I(N__5166));
    LocalMux I__461 (
            .O(N__5174),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_0 ));
    LocalMux I__460 (
            .O(N__5171),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_0 ));
    Odrv4 I__459 (
            .O(N__5166),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_0 ));
    CEMux I__458 (
            .O(N__5159),
            .I(N__5156));
    LocalMux I__457 (
            .O(N__5156),
            .I(N__5153));
    Span4Mux_h I__456 (
            .O(N__5153),
            .I(N__5150));
    Odrv4 I__455 (
            .O(N__5150),
            .I(\DUT.uart_inst0.recv_state_RNIL139CZ0Z_2 ));
    InMux I__454 (
            .O(N__5147),
            .I(N__5144));
    LocalMux I__453 (
            .O(N__5144),
            .I(\DUT.uart_inst0.g0_0_i_a3_0_3 ));
    CascadeMux I__452 (
            .O(N__5141),
            .I(\DUT.uart_inst0.g0_0_i_a3_0_4_cascade_ ));
    InMux I__451 (
            .O(N__5138),
            .I(N__5135));
    LocalMux I__450 (
            .O(N__5135),
            .I(\DUT.uart_inst0.g0_0 ));
    CascadeMux I__449 (
            .O(N__5132),
            .I(\DUT.uart_inst0.g0_i_a3_0_5_cascade_ ));
    InMux I__448 (
            .O(N__5129),
            .I(N__5126));
    LocalMux I__447 (
            .O(N__5126),
            .I(\DUT.uart_inst0.g0_i_a3_8 ));
    CascadeMux I__446 (
            .O(N__5123),
            .I(\DUT.uart_inst0.recv_state_ns_0_i_a2_0_2_3_cascade_ ));
    CascadeMux I__445 (
            .O(N__5120),
            .I(\DUT.uart_inst0.m16_N_3L3_1_cascade_ ));
    InMux I__444 (
            .O(N__5117),
            .I(N__5114));
    LocalMux I__443 (
            .O(N__5114),
            .I(\DUT.uart_inst0.rx_bits_remaining_RNO_4Z0Z_1 ));
    CascadeMux I__442 (
            .O(N__5111),
            .I(\DUT.uart_inst0.g0_i_a3_5_cascade_ ));
    InMux I__441 (
            .O(N__5108),
            .I(N__5105));
    LocalMux I__440 (
            .O(N__5105),
            .I(\PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO ));
    CascadeMux I__439 (
            .O(N__5102),
            .I(\DUT.uart_inst0.rx_bits_remaining_RNO_1Z0Z_1_cascade_ ));
    CascadeMux I__438 (
            .O(N__5099),
            .I(\DUT.uart_inst0.m5_1_1_cascade_ ));
    InMux I__437 (
            .O(N__5096),
            .I(N__5093));
    LocalMux I__436 (
            .O(N__5093),
            .I(\DUT.uart_inst0.N_6_0_0 ));
    CascadeMux I__435 (
            .O(N__5090),
            .I(\DUT.uart_inst0.N_6_0_0_cascade_ ));
    InMux I__434 (
            .O(N__5087),
            .I(N__5084));
    LocalMux I__433 (
            .O(N__5084),
            .I(\DUT.uart_inst0.N_15_mux_0 ));
    IoInMux I__432 (
            .O(N__5081),
            .I(N__5078));
    LocalMux I__431 (
            .O(N__5078),
            .I(N__5075));
    Span12Mux_s9_v I__430 (
            .O(N__5075),
            .I(N__5072));
    Span12Mux_v I__429 (
            .O(N__5072),
            .I(N__5069));
    Odrv12 I__428 (
            .O(N__5069),
            .I(BTN_N_c));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_11_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_19_0_ (
            .carryinitin(\DUT.uart_inst0.tx_clk_divider_cry_7 ),
            .carryinitout(bfn_11_19_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(\DUT.uart_inst0.rx_clk_divider_1_cry_7 ),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(\DUT.uart_inst0.rx_clk_divider_1_cry_15 ),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_11_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_22_0_));
    defparam IN_MUX_bfv_8_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_18_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_15_0_));
    ICE_GB wPllLocked_i_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__5612),
            .GLOBALBUFFEROUTPUT(wPllLocked_i_g));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB \top_pll_inst.top_pll_inst_RNISDA2  (
            .USERSIGNALTOGLOBALBUFFER(N__8363),
            .GLOBALBUFFEROUTPUT(wPllLocked_g));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0 .C_ON=1'b0;
    defparam \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0 .SEQ_MODE=4'b0000;
    defparam \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5108),
            .lcout(wPllLocked),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_1_LC_7_13_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_1_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_1_LC_7_13_0 .LUT_INIT=16'b0011010101010101;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_1_1_LC_7_13_0  (
            .in0(N__5406),
            .in1(N__5096),
            .in2(N__8362),
            .in3(N__5117),
            .lcout(),
            .ltout(\DUT.uart_inst0.rx_bits_remaining_RNO_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_1_LC_7_13_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_1_LC_7_13_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_bits_remaining_1_LC_7_13_1 .LUT_INIT=16'b0000111100100111;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_1_LC_7_13_1  (
            .in0(N__8353),
            .in1(N__5087),
            .in2(N__5102),
            .in3(N__7935),
            .lcout(\DUT.uart_inst0.rx_bits_remainingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13055),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_3_LC_7_13_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_3_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_3_LC_7_13_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_0_3_LC_7_13_2  (
            .in0(N__5404),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5204),
            .lcout(\DUT.uart_inst0.N_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNIFF651_2_LC_7_13_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNIFF651_2_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNIFF651_2_LC_7_13_4 .LUT_INIT=16'b0101010100100010;
    LogicCell40 \DUT.uart_inst0.recv_state_RNIFF651_2_LC_7_13_4  (
            .in0(N__5529),
            .in1(N__10141),
            .in2(_gnd_net_),
            .in3(N__5657),
            .lcout(),
            .ltout(\DUT.uart_inst0.m5_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIO2V22_0_LC_7_13_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIO2V22_0_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIO2V22_0_LC_7_13_5 .LUT_INIT=16'b1000010100100000;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNIO2V22_0_LC_7_13_5  (
            .in0(N__5658),
            .in1(N__5208),
            .in2(N__5099),
            .in3(N__5402),
            .lcout(\DUT.uart_inst0.N_6_0_0 ),
            .ltout(\DUT.uart_inst0.N_6_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_1_LC_7_13_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_1_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_1_LC_7_13_6 .LUT_INIT=16'b0001110101010101;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_0_1_LC_7_13_6  (
            .in0(N__5403),
            .in1(N__5417),
            .in2(N__5090),
            .in3(N__5438),
            .lcout(\DUT.uart_inst0.N_15_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_2_2_LC_7_13_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_2_2_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_2_2_LC_7_13_7 .LUT_INIT=16'b1111111101010110;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_2_2_LC_7_13_7  (
            .in0(N__5299),
            .in1(N__5405),
            .in2(N__5210),
            .in3(N__5530),
            .lcout(\DUT.uart_inst0.N_35_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_1_3_LC_7_14_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_1_3_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_1_3_LC_7_14_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_1_3_LC_7_14_0  (
            .in0(N__5295),
            .in1(N__5401),
            .in2(N__5240),
            .in3(N__5209),
            .lcout(),
            .ltout(\DUT.uart_inst0.recv_state_ns_0_i_a2_0_2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_3_LC_7_14_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_3_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_3_LC_7_14_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_3_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5123),
            .in3(N__5659),
            .lcout(\DUT.uart_inst0.recv_state_ns_0_i_a2_0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_5_1_LC_7_14_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_5_1_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_5_1_LC_7_14_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_5_1_LC_7_14_2  (
            .in0(N__6320),
            .in1(N__6731),
            .in2(_gnd_net_),
            .in3(N__6243),
            .lcout(),
            .ltout(\DUT.uart_inst0.m16_N_3L3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_4_1_LC_7_14_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_4_1_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_4_1_LC_7_14_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_4_1_LC_7_14_3  (
            .in0(N__6136),
            .in1(N__6562),
            .in2(N__5120),
            .in3(N__6795),
            .lcout(\DUT.uart_inst0.rx_bits_remaining_RNO_4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_6_2_LC_7_14_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_6_2_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_6_2_LC_7_14_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_6_2_LC_7_14_4  (
            .in0(N__5511),
            .in1(N__6242),
            .in2(N__10171),
            .in3(N__6730),
            .lcout(\DUT.uart_inst0.m9_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_3_4_LC_7_14_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_3_4_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_3_4_LC_7_14_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_3_4_LC_7_14_5  (
            .in0(N__6244),
            .in1(N__6321),
            .in2(N__6142),
            .in3(N__6563),
            .lcout(\DUT.uart_inst0.N_81_mux_i_i_a5_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_4_LC_7_14_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_4_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_4_LC_7_14_6 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_4_LC_7_14_6  (
            .in0(N__12060),
            .in1(N__6058),
            .in2(_gnd_net_),
            .in3(N__10041),
            .lcout(\DUT.uart_inst0.N_81_mux_i_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_6_2_LC_7_15_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_6_2_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_6_2_LC_7_15_1 .LUT_INIT=16'b1000101010001000;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_6_2_LC_7_15_1  (
            .in0(N__8336),
            .in1(N__5642),
            .in2(N__10172),
            .in3(N__5507),
            .lcout(\DUT.uart_inst0.g0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_9_2_LC_7_15_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_9_2_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_9_2_LC_7_15_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_9_2_LC_7_15_2  (
            .in0(N__6427),
            .in1(N__6491),
            .in2(N__5203),
            .in3(N__6713),
            .lcout(),
            .ltout(\DUT.uart_inst0.g0_i_a3_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_4_2_LC_7_15_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_4_2_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_4_2_LC_7_15_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_4_2_LC_7_15_3  (
            .in0(N__5366),
            .in1(N__5236),
            .in2(N__5111),
            .in3(N__5312),
            .lcout(\DUT.uart_inst0.g0_i_a3_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNI69LM2_0_0_LC_7_15_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNI69LM2_0_0_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNI69LM2_0_0_LC_7_15_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNI69LM2_0_0_LC_7_15_4  (
            .in0(N__6553),
            .in1(N__6712),
            .in2(N__6252),
            .in3(N__6314),
            .lcout(\DUT.uart_inst0.g0_0_i_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_0_LC_7_15_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_0_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_0_LC_7_15_5 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_0_LC_7_15_5  (
            .in0(N__10165),
            .in1(N__9976),
            .in2(_gnd_net_),
            .in3(N__7142),
            .lcout(\DUT.uart_inst0.recv_state_ns_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_2_2_LC_7_15_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_2_2_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_2_2_LC_7_15_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_2_2_LC_7_15_6  (
            .in0(N__5235),
            .in1(N__6316),
            .in2(N__6566),
            .in3(N__6249),
            .lcout(\DUT.uart_inst0.g0_i_a3_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_7_2_LC_7_15_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_7_2_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_7_2_LC_7_15_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_7_2_LC_7_15_7  (
            .in0(N__6315),
            .in1(N__6126),
            .in2(N__6796),
            .in3(N__6554),
            .lcout(\DUT.uart_inst0.m9_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNIS6O94_0_LC_7_16_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNIS6O94_0_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNIS6O94_0_LC_7_16_0 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNIS6O94_0_LC_7_16_0  (
            .in0(N__6788),
            .in1(_gnd_net_),
            .in2(N__6141),
            .in3(N__5147),
            .lcout(),
            .ltout(\DUT.uart_inst0.g0_0_i_a3_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNIL139C_2_LC_7_16_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNIL139C_2_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNIL139C_2_LC_7_16_1 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNIL139C_2_LC_7_16_1  (
            .in0(N__5138),
            .in1(N__5669),
            .in2(N__5141),
            .in3(N__7937),
            .lcout(\DUT.uart_inst0.recv_state_RNIL139CZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNIBTG71_2_LC_7_16_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNIBTG71_2_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNIBTG71_2_LC_7_16_2 .LUT_INIT=16'b1101110000000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNIBTG71_2_LC_7_16_2  (
            .in0(N__10169),
            .in1(N__5644),
            .in2(N__5528),
            .in3(N__12066),
            .lcout(\DUT.uart_inst0.g0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_8_2_LC_7_16_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_8_2_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_8_2_LC_7_16_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_8_2_LC_7_16_3  (
            .in0(N__5310),
            .in1(N__5408),
            .in2(_gnd_net_),
            .in3(N__6789),
            .lcout(),
            .ltout(\DUT.uart_inst0.g0_i_a3_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_3_2_LC_7_16_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_3_2_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_3_2_LC_7_16_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_3_2_LC_7_16_4  (
            .in0(N__6130),
            .in1(N__5187),
            .in2(N__5132),
            .in3(N__6734),
            .lcout(),
            .ltout(\DUT.uart_inst0.g0_i_a3_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_2_LC_7_16_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_2_LC_7_16_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_2_LC_7_16_5 .LUT_INIT=16'b0011111101010101;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_2_LC_7_16_5  (
            .in0(N__5129),
            .in1(N__5264),
            .in2(N__5258),
            .in3(N__7936),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_2_LC_7_16_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_2_LC_7_16_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_2_LC_7_16_6 .LUT_INIT=16'b1010101010000000;
    LogicCell40 \DUT.uart_inst0.recv_state_2_LC_7_16_6  (
            .in0(N__8352),
            .in1(N__5645),
            .in2(N__5255),
            .in3(N__5570),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13048),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_3_LC_7_17_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_3_LC_7_17_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_bits_remaining_3_LC_7_17_0 .LUT_INIT=16'b1111111110101001;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_3_LC_7_17_0  (
            .in0(N__5234),
            .in1(N__5311),
            .in2(N__5252),
            .in3(N__5534),
            .lcout(\DUT.uart_inst0.rx_bits_remainingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13043),
            .ce(N__5159),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_0_LC_7_17_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_0_LC_7_17_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_bits_remaining_0_LC_7_17_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_0_LC_7_17_1  (
            .in0(N__5533),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5188),
            .lcout(\DUT.uart_inst0.rx_bits_remainingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13043),
            .ce(N__5159),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_7_19_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_7_19_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_7_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7418),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13037),
            .ce(N__7487),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_7_19_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_7_19_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_7_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7374),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13037),
            .ce(N__7487),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_7_19_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_7_19_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_7_19_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_7_19_2  (
            .in0(N__7326),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13037),
            .ce(N__7487),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_7_19_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_7_19_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_7_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7809),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13037),
            .ce(N__7487),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_7_19_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_7_19_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_7_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7754),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13037),
            .ce(N__7487),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_7_19_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_7_19_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_7_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7703),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13037),
            .ce(N__7487),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_7_19_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_7_19_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_7_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7652),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13037),
            .ce(N__7487),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_7_19_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_7_19_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_7_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_7_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10491),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13037),
            .ce(N__7487),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_7_20_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_7_20_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_7_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_7_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13088),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13032),
            .ce(N__7205),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_7_20_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_7_20_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_7_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_7_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13277),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13032),
            .ce(N__7205),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_7_20_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_7_20_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_7_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_7_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12497),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13032),
            .ce(N__7205),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_7_20_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_7_20_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_7_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_7_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12421),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13032),
            .ce(N__7205),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_7_20_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_7_20_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_7_20_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_7_20_4  (
            .in0(N__12381),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13032),
            .ce(N__7205),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_7_20_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_7_20_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_7_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_7_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13130),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13032),
            .ce(N__7205),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_7_20_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_7_20_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_7_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_7_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13209),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13032),
            .ce(N__7205),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_7_20_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_7_20_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_7_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_7_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13319),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13032),
            .ce(N__7205),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_7_21_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_7_21_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_7_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_7_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7422),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13027),
            .ce(N__10441),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_7_21_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_7_21_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_7_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_7_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7376),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13027),
            .ce(N__10441),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_7_21_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_7_21_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_7_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_7_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7327),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13027),
            .ce(N__10441),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_7_21_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_7_21_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_7_21_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_7_21_4  (
            .in0(N__7758),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13027),
            .ce(N__10441),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_7_21_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_7_21_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_7_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_7_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7707),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13027),
            .ce(N__10441),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_7_21_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_7_21_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_7_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_7_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7655),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13027),
            .ce(N__10441),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_7_22_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_7_22_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_7_22_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_7_22_4  (
            .in0(N__7810),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13021),
            .ce(N__10437),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_2_LC_8_13_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_2_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_2_LC_8_13_0 .LUT_INIT=16'b0010011100000000;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_0_2_LC_8_13_0  (
            .in0(N__7913),
            .in1(N__6334),
            .in2(N__6869),
            .in3(N__5330),
            .lcout(),
            .ltout(\DUT.uart_inst0.g0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_2_LC_8_13_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_2_LC_8_13_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_bits_remaining_2_LC_8_13_1 .LUT_INIT=16'b0101110011001100;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_2_LC_8_13_1  (
            .in0(N__5321),
            .in1(N__5306),
            .in2(N__5315),
            .in3(N__6161),
            .lcout(\DUT.uart_inst0.rx_bits_remainingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13054),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_6_LC_8_13_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_6_LC_8_13_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_6_LC_8_13_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \DUT.uart_inst0.recv_state_6_LC_8_13_2  (
            .in0(N__8358),
            .in1(N__5348),
            .in2(N__10140),
            .in3(N__6042),
            .lcout(\DUT.wRcvd ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13054),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_3_1_LC_8_13_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_3_1_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_3_1_LC_8_13_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_3_1_LC_8_13_3  (
            .in0(N__6852),
            .in1(N__6428),
            .in2(N__6959),
            .in3(N__6493),
            .lcout(\DUT.uart_inst0.m8_e_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_10_2_LC_8_13_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_10_2_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_10_2_LC_8_13_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_10_2_LC_8_13_4  (
            .in0(N__6993),
            .in1(N__6955),
            .in2(N__5407),
            .in3(N__6851),
            .lcout(\DUT.uart_inst0.g0_i_a3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_2_2_LC_8_13_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_2_2_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_2_2_LC_8_13_5 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_2_2_LC_8_13_5  (
            .in0(N__5531),
            .in1(N__10116),
            .in2(_gnd_net_),
            .in3(N__5663),
            .lcout(\DUT.uart_inst0.rx_countdown_RNO_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_5_LC_8_13_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_5_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_5_LC_8_13_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_5_LC_8_13_6  (
            .in0(N__10115),
            .in1(N__5346),
            .in2(_gnd_net_),
            .in3(N__5532),
            .lcout(\DUT.uart_inst0.N_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_3_LC_8_13_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_3_LC_8_13_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_3_LC_8_13_7 .LUT_INIT=16'b1000110010000000;
    LogicCell40 \DUT.uart_inst0.recv_state_3_LC_8_13_7  (
            .in0(N__5347),
            .in1(N__8357),
            .in2(N__6047),
            .in3(N__5357),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13054),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_3_2_LC_8_14_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_3_2_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_3_2_LC_8_14_0 .LUT_INIT=16'b0010000010101000;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_3_2_LC_8_14_0  (
            .in0(N__5336),
            .in1(N__6697),
            .in2(N__6263),
            .in3(N__6793),
            .lcout(\DUT.uart_inst0.g0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_1_LC_8_14_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_1_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_1_LC_8_14_1 .LUT_INIT=16'b0101010111110111;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_1_LC_8_14_1  (
            .in0(N__12059),
            .in1(N__9968),
            .in2(N__10161),
            .in3(N__5522),
            .lcout(\DUT.uart_inst0.N_81_mux_i_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_3_1_LC_8_14_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_3_1_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_3_1_LC_8_14_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_3_1_LC_8_14_2  (
            .in0(N__6132),
            .in1(N__6792),
            .in2(N__6333),
            .in3(N__6561),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_81_mux_i_i_a5_0_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_1_1_LC_8_14_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_1_1_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_1_1_LC_8_14_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_1_1_LC_8_14_3  (
            .in0(N__6699),
            .in1(N__9565),
            .in2(N__5324),
            .in3(N__6248),
            .lcout(\DUT.uart_inst0.N_81_mux_i_i_a5_0_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_1_4_LC_8_14_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_1_4_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_1_4_LC_8_14_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_1_4_LC_8_14_4  (
            .in0(N__10039),
            .in1(N__5462),
            .in2(N__6729),
            .in3(N__6794),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_81_mux_i_i_a5_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_4_LC_8_14_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_4_LC_8_14_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_4_LC_8_14_5 .LUT_INIT=16'b0000010100010001;
    LogicCell40 \DUT.uart_inst0.recv_state_4_LC_8_14_5  (
            .in0(N__5453),
            .in1(N__5444),
            .in2(N__5447),
            .in3(N__7917),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13052),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_4_2_LC_8_14_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_4_2_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_4_2_LC_8_14_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_4_2_LC_8_14_6  (
            .in0(N__6131),
            .in1(N__6560),
            .in2(N__6254),
            .in3(N__6791),
            .lcout(\DUT.uart_inst0.N_13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_2_4_LC_8_14_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_2_4_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_2_4_LC_8_14_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_2_4_LC_8_14_7  (
            .in0(N__6698),
            .in1(N__5960),
            .in2(N__10035),
            .in3(N__6853),
            .lcout(\DUT.uart_inst0.N_81_mux_i_i_a5_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_2_1_LC_8_15_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_2_1_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_2_1_LC_8_15_0 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_2_1_LC_8_15_0  (
            .in0(N__7002),
            .in1(_gnd_net_),
            .in2(N__6711),
            .in3(_gnd_net_),
            .lcout(\DUT.uart_inst0.m8_e_2 ),
            .ltout(),
            .carryin(bfn_8_15_0_),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_s1_c_RNIKPDT_LC_8_15_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_s1_c_RNIKPDT_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_s1_c_RNIKPDT_LC_8_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_0_s1_c_RNIKPDT_LC_8_15_1  (
            .in0(_gnd_net_),
            .in1(N__12747),
            .in2(N__6492),
            .in3(N__5429),
            .lcout(\DUT.uart_inst0.rx_countdown_3_s1_1 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_countdown_3_cry_0_s1 ),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNIMVNN_LC_8_15_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNIMVNN_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNIMVNN_LC_8_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNIMVNN_LC_8_15_2  (
            .in0(_gnd_net_),
            .in1(N__6858),
            .in2(N__12807),
            .in3(N__5426),
            .lcout(\DUT.uart_inst0.rx_countdown_3_s1_2 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_countdown_3_cry_1_s1 ),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_2_s1_c_RNIO52I_LC_8_15_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_2_s1_c_RNIO52I_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_2_s1_c_RNIO52I_LC_8_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_2_s1_c_RNIO52I_LC_8_15_3  (
            .in0(_gnd_net_),
            .in1(N__12751),
            .in2(N__6947),
            .in3(N__5423),
            .lcout(\DUT.uart_inst0.rx_countdown_3_s1_3 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_countdown_3_cry_2_s1 ),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_s1_c_RNIQBCS_LC_8_15_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_s1_c_RNIQBCS_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_s1_c_RNIQBCS_LC_8_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_3_s1_c_RNIQBCS_LC_8_15_4  (
            .in0(_gnd_net_),
            .in1(N__12752),
            .in2(N__7019),
            .in3(N__5420),
            .lcout(\DUT.uart_inst0.rx_countdown_3_s1_4 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_countdown_3_cry_3_s1 ),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_4_s1_c_RNISHMM_LC_8_15_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_4_s1_c_RNISHMM_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_4_s1_c_RNISHMM_LC_8_15_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_4_s1_c_RNISHMM_LC_8_15_5  (
            .in0(_gnd_net_),
            .in1(N__6400),
            .in2(_gnd_net_),
            .in3(N__5585),
            .lcout(\DUT.uart_inst0.rx_countdown_3_s1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_1_2_LC_8_15_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_1_2_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_1_2_LC_8_15_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_1_2_LC_8_15_6  (
            .in0(N__5582),
            .in1(N__5576),
            .in2(N__5546),
            .in3(N__7899),
            .lcout(\DUT.uart_inst0.N_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_1_LC_8_15_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_1_LC_8_15_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_1_LC_8_15_7 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \DUT.uart_inst0.recv_state_1_LC_8_15_7  (
            .in0(N__7900),
            .in1(N__6182),
            .in2(N__5564),
            .in3(N__5555),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13049),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_12_2_LC_8_16_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_12_2_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_12_2_LC_8_16_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_12_2_LC_8_16_0  (
            .in0(N__6479),
            .in1(N__6871),
            .in2(N__6420),
            .in3(N__6686),
            .lcout(),
            .ltout(\DUT.uart_inst0.m4_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_5_2_LC_8_16_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_5_2_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_5_2_LC_8_16_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_5_2_LC_8_16_1  (
            .in0(N__5468),
            .in1(N__7030),
            .in2(N__5549),
            .in3(N__6940),
            .lcout(\DUT.uart_inst0.N_18_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_1_LC_8_16_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_1_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_1_LC_8_16_2 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_0_1_LC_8_16_2  (
            .in0(N__6480),
            .in1(N__7925),
            .in2(N__10046),
            .in3(N__6251),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_297_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_1_LC_8_16_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_1_LC_8_16_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_1_LC_8_16_3 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \DUT.uart_inst0.rx_countdown_1_LC_8_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5537),
            .in3(N__9541),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13044),
            .ce(N__12000),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_11_2_LC_8_16_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_11_2_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_11_2_LC_8_16_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_11_2_LC_8_16_4  (
            .in0(N__5506),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10146),
            .lcout(\DUT.uart_inst0.N_15_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNIPHLT1_5_LC_8_16_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNIPHLT1_5_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNIPHLT1_5_LC_8_16_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNIPHLT1_5_LC_8_16_5  (
            .in0(N__6685),
            .in1(N__6939),
            .in2(N__6424),
            .in3(N__6478),
            .lcout(),
            .ltout(\DUT.uart_inst0.g0_0_i_a3_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNI7CGS2_2_LC_8_16_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNI7CGS2_2_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNI7CGS2_2_LC_8_16_6 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNI7CGS2_2_LC_8_16_6  (
            .in0(N__7031),
            .in1(_gnd_net_),
            .in2(N__5672),
            .in3(N__6872),
            .lcout(\DUT.uart_inst0.g0_0_i_a3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNIEQQU_5_LC_8_16_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNIEQQU_5_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNIEQQU_5_LC_8_16_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNIEQQU_5_LC_8_16_7  (
            .in0(_gnd_net_),
            .in1(N__6396),
            .in2(_gnd_net_),
            .in3(N__6477),
            .lcout(\DUT.uart_inst0.N_13_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNI8P9F_2_LC_8_17_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNI8P9F_2_LC_8_17_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNI8P9F_2_LC_8_17_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNI8P9F_2_LC_8_17_0  (
            .in0(_gnd_net_),
            .in1(N__12064),
            .in2(_gnd_net_),
            .in3(N__5643),
            .lcout(\DUT.uart_inst0.m11_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNISAK33_LC_8_17_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNISAK33_LC_8_17_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNISAK33_LC_8_17_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNISAK33_LC_8_17_2  (
            .in0(N__6565),
            .in1(N__6140),
            .in2(N__6335),
            .in3(N__6250),
            .lcout(\DUT.uart_inst0.m10_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.wPllLocked_i_LC_8_17_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.wPllLocked_i_LC_8_17_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.wPllLocked_i_LC_8_17_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \DUT.uart_inst0.wPllLocked_i_LC_8_17_7  (
            .in0(N__12065),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(wPllLocked_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_LC_8_18_0 .C_ON=1'b1;
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_LC_8_18_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_LC_8_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_LC_8_18_0  (
            .in0(_gnd_net_),
            .in1(N__7148),
            .in2(N__7076),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_18_0_),
            .carryout(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_1_LC_8_18_1 .C_ON=1'b1;
    defparam \DUT.fifo_rx_inst.rFifoCount_1_LC_8_18_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoCount_1_LC_8_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_1_LC_8_18_1  (
            .in0(_gnd_net_),
            .in1(N__7233),
            .in2(N__5684),
            .in3(N__5591),
            .lcout(\DUT.fifo_rx_inst.rFifoCountZ0Z_1 ),
            .ltout(),
            .carryin(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0 ),
            .carryout(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1 ),
            .clk(N__13038),
            .ce(),
            .sr(N__10527));
    defparam \DUT.fifo_rx_inst.rFifoCount_2_LC_8_18_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_2_LC_8_18_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoCount_2_LC_8_18_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_2_LC_8_18_2  (
            .in0(_gnd_net_),
            .in1(N__5696),
            .in2(_gnd_net_),
            .in3(N__5588),
            .lcout(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13038),
            .ce(),
            .sr(N__10527));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_2_1_LC_8_19_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_2_1_LC_8_19_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_2_1_LC_8_19_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI96D91_2_1_LC_8_19_0  (
            .in0(N__5800),
            .in1(N__7130),
            .in2(N__5833),
            .in3(N__7271),
            .lcout(\DUT.fifo_rx_inst.rFifoData_awe3 ),
            .ltout(\DUT.fifo_rx_inst.rFifoData_awe3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1_1_LC_8_19_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1_1_LC_8_19_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1_1_LC_8_19_1 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1_1_LC_8_19_1  (
            .in0(N__12070),
            .in1(_gnd_net_),
            .in2(N__5702),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.un1_i11_i ),
            .ltout(\DUT.fifo_rx_inst.un1_i11_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_0_LC_8_19_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_0_LC_8_19_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rWritePtr_0_LC_8_19_2 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_0_LC_8_19_2  (
            .in0(N__5822),
            .in1(_gnd_net_),
            .in2(N__5699),
            .in3(N__5857),
            .lcout(\DUT.fifo_rx_inst.rWritePtrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13033),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNO_0_2_LC_8_19_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNO_0_2_LC_8_19_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNO_0_2_LC_8_19_3 .LUT_INIT=16'b1100110011000110;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNO_0_2_LC_8_19_3  (
            .in0(N__10653),
            .in1(N__7273),
            .in2(N__7141),
            .in3(N__8223),
            .lcout(\DUT.fifo_rx_inst.un1_rFifoCount_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_LC_8_19_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_LC_8_19_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_LC_8_19_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_LC_8_19_4  (
            .in0(N__7272),
            .in1(N__7229),
            .in2(_gnd_net_),
            .in3(N__7072),
            .lcout(N_92_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_1_LC_8_19_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_1_LC_8_19_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rWritePtr_1_LC_8_19_6 .LUT_INIT=16'b0001001000100010;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_1_LC_8_19_6  (
            .in0(N__5801),
            .in1(N__5690),
            .in2(N__5834),
            .in3(N__5858),
            .lcout(\DUT.fifo_rx_inst.rWritePtrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13033),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIK3G92_1_LC_8_19_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIK3G92_1_LC_8_19_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIK3G92_1_LC_8_19_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNIK3G92_1_LC_8_19_7  (
            .in0(N__7131),
            .in1(N__10652),
            .in2(N__7235),
            .in3(N__8222),
            .lcout(\DUT.fifo_rx_inst.rFifoCount_RNIK3G92Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_8_20_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_8_20_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_8_20_1 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_8_20_1  (
            .in0(N__5803),
            .in1(_gnd_net_),
            .in2(N__5840),
            .in3(N__5855),
            .lcout(\DUT.fifo_rx_inst.rFifoData_awe0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_8_20_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_8_20_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_8_20_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_8_20_3  (
            .in0(_gnd_net_),
            .in1(N__7106),
            .in2(_gnd_net_),
            .in3(N__7274),
            .lcout(\DUT.fifo_rx_inst.rWritePtr16 ),
            .ltout(\DUT.fifo_rx_inst.rWritePtr16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_8_20_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_8_20_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_8_20_4 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_8_20_4  (
            .in0(_gnd_net_),
            .in1(N__5835),
            .in2(N__5675),
            .in3(N__5802),
            .lcout(\DUT.fifo_rx_inst.rFifoData_awe1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_1_LC_8_20_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_1_LC_8_20_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_1_LC_8_20_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_0_1_LC_8_20_5  (
            .in0(N__11437),
            .in1(N__11606),
            .in2(_gnd_net_),
            .in3(N__11686),
            .lcout(\DUT.uart_inst0.N_8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_8_20_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_8_20_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_8_20_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_8_20_6  (
            .in0(N__5856),
            .in1(N__5839),
            .in2(_gnd_net_),
            .in3(N__5804),
            .lcout(\DUT.fifo_rx_inst.rFifoData_awe2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_8_20_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_8_20_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_8_20_7 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_8_20_7  (
            .in0(N__8977),
            .in1(N__5783),
            .in2(N__6017),
            .in3(N__8182),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rTxByte_esr_6_LC_8_21_0.C_ON=1'b0;
    defparam rTxByte_esr_6_LC_8_21_0.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_6_LC_8_21_0.LUT_INIT=16'b1010000011011101;
    LogicCell40 rTxByte_esr_6_LC_8_21_0 (
            .in0(N__9017),
            .in1(N__7610),
            .in2(N__5777),
            .in3(N__5720),
            .lcout(rTxByteZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13022),
            .ce(N__8877),
            .sr(N__8844));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_8_21_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_8_21_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_8_21_1 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_8_21_1  (
            .in0(N__5765),
            .in1(N__9010),
            .in2(N__5996),
            .in3(N__8197),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rTxByte_esr_4_LC_8_21_2.C_ON=1'b0;
    defparam rTxByte_esr_4_LC_8_21_2.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_4_LC_8_21_2.LUT_INIT=16'b1000111110000101;
    LogicCell40 rTxByte_esr_4_LC_8_21_2 (
            .in0(N__9015),
            .in1(N__5756),
            .in2(N__5747),
            .in3(N__7715),
            .lcout(rTxByteZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13022),
            .ce(N__8877),
            .sr(N__8844));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_8_21_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_8_21_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_8_21_3 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_8_21_3  (
            .in0(N__5744),
            .in1(N__9011),
            .in2(N__5984),
            .in3(N__8198),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rTxByte_esr_5_LC_8_21_4.C_ON=1'b0;
    defparam rTxByte_esr_5_LC_8_21_4.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_5_LC_8_21_4.LUT_INIT=16'b1010110100001101;
    LogicCell40 rTxByte_esr_5_LC_8_21_4 (
            .in0(N__9016),
            .in1(N__7664),
            .in2(N__5738),
            .in3(N__5735),
            .lcout(rTxByteZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13022),
            .ce(N__8877),
            .sr(N__8844));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_8_21_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_8_21_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_8_21_5 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_8_21_5  (
            .in0(N__5726),
            .in1(N__9009),
            .in2(N__5972),
            .in3(N__8195),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_8_21_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_8_21_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_8_21_6 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_8_21_6  (
            .in0(N__8196),
            .in1(N__6005),
            .in2(N__9025),
            .in3(N__5711),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rTxByte_esr_3_LC_8_21_7.C_ON=1'b0;
    defparam rTxByte_esr_3_LC_8_21_7.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_3_LC_8_21_7.LUT_INIT=16'b1100101000001111;
    LogicCell40 rTxByte_esr_3_LC_8_21_7 (
            .in0(N__7766),
            .in1(N__5948),
            .in2(N__5939),
            .in3(N__9018),
            .lcout(rTxByteZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13022),
            .ce(N__8877),
            .sr(N__8844));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_8_22_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_8_22_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_8_22_0 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_8_22_0  (
            .in0(N__8194),
            .in1(N__5873),
            .in2(N__5936),
            .in3(N__9019),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rTxByte_esr_0_LC_8_22_1.C_ON=1'b0;
    defparam rTxByte_esr_0_LC_8_22_1.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_0_LC_8_22_1.LUT_INIT=16'b1100101000001111;
    LogicCell40 rTxByte_esr_0_LC_8_22_1 (
            .in0(N__7385),
            .in1(N__5927),
            .in2(N__5915),
            .in3(N__9005),
            .lcout(rTxByteZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13016),
            .ce(N__8879),
            .sr(N__8852));
    defparam rTxByte_esr_7_LC_8_22_2.C_ON=1'b0;
    defparam rTxByte_esr_7_LC_8_22_2.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_7_LC_8_22_2.LUT_INIT=16'b1011100000110011;
    LogicCell40 rTxByte_esr_7_LC_8_22_2 (
            .in0(N__5912),
            .in1(N__7556),
            .in2(N__7598),
            .in3(N__9020),
            .lcout(rTxByteZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13016),
            .ce(N__8879),
            .sr(N__8852));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_8_22_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_8_22_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_8_22_5 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_8_22_5  (
            .in0(N__5900),
            .in1(N__9004),
            .in2(N__5867),
            .in3(N__8193),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rTxByte_esr_2_LC_8_22_6.C_ON=1'b0;
    defparam rTxByte_esr_2_LC_8_22_6.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_2_LC_8_22_6.LUT_INIT=16'b1011001110000011;
    LogicCell40 rTxByte_esr_2_LC_8_22_6 (
            .in0(N__5894),
            .in1(N__5882),
            .in2(N__9024),
            .in3(N__7280),
            .lcout(rTxByteZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13016),
            .ce(N__8879),
            .sr(N__8852));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_8_23_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_8_23_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_8_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_8_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7427),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13011),
            .ce(N__7511),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_8_23_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_8_23_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_8_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_8_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7375),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13011),
            .ce(N__7511),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_8_23_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_8_23_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_8_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_8_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7328),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13011),
            .ce(N__7511),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_8_23_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_8_23_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_8_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_8_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7814),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13011),
            .ce(N__7511),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_8_23_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_8_23_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_8_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_8_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7759),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13011),
            .ce(N__7511),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_8_23_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_8_23_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_8_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_8_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7708),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13011),
            .ce(N__7511),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_8_23_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_8_23_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_8_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_8_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7654),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13011),
            .ce(N__7511),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_8_23_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_8_23_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_8_23_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_8_23_7  (
            .in0(N__10492),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13011),
            .ce(N__7511),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_4_4_LC_9_13_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_4_4_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_4_4_LC_9_13_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_4_4_LC_9_13_0  (
            .in0(N__6954),
            .in1(N__6425),
            .in2(N__7018),
            .in3(N__6494),
            .lcout(\DUT.uart_inst0.N_81_mux_i_i_a5_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_4_LC_9_13_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_4_LC_9_13_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_4_LC_9_13_1 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_4_LC_9_13_1  (
            .in0(N__6143),
            .in1(N__9938),
            .in2(N__7923),
            .in3(N__6998),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13053),
            .ce(N__11980),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_4_2_LC_9_13_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_4_2_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_4_2_LC_9_13_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_4_2_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__6994),
            .in2(_gnd_net_),
            .in3(N__6953),
            .lcout(\DUT.uart_inst0.G_9_i_o4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_9_13_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_9_13_4 .LUT_INIT=16'b0100000001000011;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_9_13_4  (
            .in0(N__5954),
            .in1(N__7895),
            .in2(N__6733),
            .in3(N__6344),
            .lcout(),
            .ltout(\DUT.uart_inst0.G_21_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_2_LC_9_13_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_2_LC_9_13_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_2_LC_9_13_5 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_2_LC_9_13_5  (
            .in0(N__6176),
            .in1(N__9566),
            .in2(N__6170),
            .in3(N__6068),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13053),
            .ce(N__11980),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_2_LC_9_13_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_2_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_2_LC_9_13_6 .LUT_INIT=16'b0100010001000010;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_1_2_LC_9_13_6  (
            .in0(N__6077),
            .in1(N__7894),
            .in2(N__6732),
            .in3(N__6167),
            .lcout(\DUT.uart_inst0.g0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_s1_c_RNIMT2J1_LC_9_14_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_s1_c_RNIMT2J1_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_s1_c_RNIMT2J1_LC_9_14_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_3_s1_c_RNIMT2J1_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__6125),
            .in2(_gnd_net_),
            .in3(N__6790),
            .lcout(),
            .ltout(\DUT.uart_inst0.G_16_i_a3_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNIA4I1B_0_LC_9_14_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNIA4I1B_0_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNIA4I1B_0_LC_9_14_1 .LUT_INIT=16'b0011111101010101;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNIA4I1B_0_LC_9_14_1  (
            .in0(N__6503),
            .in1(N__6269),
            .in2(N__6155),
            .in3(N__7893),
            .lcout(\DUT.uart_inst0.N_45 ),
            .ltout(\DUT.uart_inst0.N_45_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_5_LC_9_14_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_5_LC_9_14_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_5_LC_9_14_2 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \DUT.uart_inst0.recv_state_5_LC_9_14_2  (
            .in0(N__8328),
            .in1(_gnd_net_),
            .in2(N__6152),
            .in3(N__6149),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13050),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_5_2_LC_9_14_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_5_2_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_5_2_LC_9_14_3 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_5_2_LC_9_14_3  (
            .in0(N__6124),
            .in1(N__6558),
            .in2(N__6253),
            .in3(N__6696),
            .lcout(\DUT.uart_inst0.N_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNI7H9R3_10_LC_9_14_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI7H9R3_10_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI7H9R3_10_LC_9_14_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNI7H9R3_10_LC_9_14_4  (
            .in0(N__7958),
            .in1(N__7829),
            .in2(N__7823),
            .in3(N__7943),
            .lcout(\DUT.uart_inst0.un2_rx_clk_divider_0 ),
            .ltout(\DUT.uart_inst0.un2_rx_clk_divider_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_9_14_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_9_14_5 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_9_14_5  (
            .in0(N__10019),
            .in1(N__6325),
            .in2(N__6071),
            .in3(N__6854),
            .lcout(\DUT.uart_inst0.G_21_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_0_LC_9_14_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_0_LC_9_14_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_0_LC_9_14_6 .LUT_INIT=16'b0010111111111111;
    LogicCell40 \DUT.uart_inst0.recv_state_0_LC_9_14_6  (
            .in0(N__6062),
            .in1(N__6046),
            .in2(N__8348),
            .in3(N__6029),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13050),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNI69LM2_0_LC_9_14_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNI69LM2_0_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNI69LM2_0_LC_9_14_7 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNI69LM2_0_LC_9_14_7  (
            .in0(N__6238),
            .in1(N__6559),
            .in2(N__6332),
            .in3(N__6695),
            .lcout(\DUT.uart_inst0.G_16_i_a3_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_5_LC_9_15_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_5_LC_9_15_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_5_LC_9_15_1 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_5_LC_9_15_1  (
            .in0(N__6781),
            .in1(N__9937),
            .in2(N__6426),
            .in3(N__7920),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13045),
            .ce(N__11989),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_7_2_LC_9_15_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_7_2_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_7_2_LC_9_15_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_7_2_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__6412),
            .in2(_gnd_net_),
            .in3(N__6487),
            .lcout(\DUT.uart_inst0.g1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_0_LC_9_15_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_0_LC_9_15_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_0_LC_9_15_3 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \DUT.uart_inst0.rx_countdown_0_LC_9_15_3  (
            .in0(N__6688),
            .in1(N__9936),
            .in2(_gnd_net_),
            .in3(N__7918),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13045),
            .ce(N__11989),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNI2GC23_0_LC_9_15_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNI2GC23_0_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNI2GC23_0_LC_9_15_4 .LUT_INIT=16'b0000000001001111;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNI2GC23_0_LC_9_15_4  (
            .in0(N__6234),
            .in1(N__6687),
            .in2(N__6890),
            .in3(N__6780),
            .lcout(\DUT.uart_inst0.N_15_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_3_LC_9_15_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_3_LC_9_15_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_3_LC_9_15_5 .LUT_INIT=16'b1111111111010111;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_3_LC_9_15_5  (
            .in0(N__9564),
            .in1(N__9181),
            .in2(N__9167),
            .in3(N__7919),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13045),
            .ce(N__11989),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIMQ571_1_LC_9_15_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIMQ571_1_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIMQ571_1_LC_9_15_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIMQ571_1_LC_9_15_6  (
            .in0(N__9180),
            .in1(N__9646),
            .in2(N__9491),
            .in3(N__9219),
            .lcout(\DUT.uart_inst0.un2_rx_clk_divider_a_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_LC_9_15_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_1_LC_9_15_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_LC_9_15_7 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_LC_9_15_7  (
            .in0(N__9220),
            .in1(N__9206),
            .in2(_gnd_net_),
            .in3(N__9580),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13045),
            .ce(N__11989),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_2_1_LC_9_16_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_2_1_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_2_1_LC_9_16_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_2_1_LC_9_16_0  (
            .in0(N__9539),
            .in1(N__6405),
            .in2(N__6575),
            .in3(N__6483),
            .lcout(\DUT.uart_inst0.N_81_mux_i_i_a5_1_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_4_1_LC_9_16_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_4_1_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_4_1_LC_9_16_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_4_1_LC_9_16_1  (
            .in0(N__6863),
            .in1(N__6937),
            .in2(N__7034),
            .in3(N__6679),
            .lcout(\DUT.uart_inst0.N_81_mux_i_i_a5_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_3_LC_9_16_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_3_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_3_LC_9_16_2 .LUT_INIT=16'b0000000100001101;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_0_3_LC_9_16_2  (
            .in0(N__6938),
            .in1(N__7924),
            .in2(N__10045),
            .in3(N__6564),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_300_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_LC_9_16_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_LC_9_16_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_3_LC_9_16_3 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6509),
            .in3(N__9540),
            .lcout(\DUT.uart_inst0.rx_countdownZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13041),
            .ce(N__11993),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNI237O_0_LC_9_16_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNI237O_0_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNI237O_0_LC_9_16_4 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \DUT.uart_inst0.recv_state_RNI237O_0_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(N__10145),
            .in2(_gnd_net_),
            .in3(N__9969),
            .lcout(\DUT.uart_inst0.N_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNIPHLT1_2_LC_9_16_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNIPHLT1_2_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNIPHLT1_2_LC_9_16_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNIPHLT1_2_LC_9_16_5  (
            .in0(N__6862),
            .in1(N__6935),
            .in2(N__7032),
            .in3(N__6678),
            .lcout(),
            .ltout(\DUT.uart_inst0.G_16_i_a3_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNI7CGS2_5_LC_9_16_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNI7CGS2_5_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNI7CGS2_5_LC_9_16_6 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNI7CGS2_5_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(N__6404),
            .in2(N__6506),
            .in3(N__6481),
            .lcout(\DUT.uart_inst0.G_16_i_a3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_3_2_LC_9_16_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_3_2_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_3_2_LC_9_16_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_3_2_LC_9_16_7  (
            .in0(N__6482),
            .in1(N__6419),
            .in2(N__7033),
            .in3(N__6936),
            .lcout(\DUT.uart_inst0.N_11_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_0_LC_9_17_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_0_LC_9_17_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rWritePtr_0_LC_9_17_0 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_0_LC_9_17_0  (
            .in0(N__8568),
            .in1(N__7043),
            .in2(_gnd_net_),
            .in3(N__8485),
            .lcout(\DUT.fifo_tx_inst.rWritePtrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13039),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_2_1_LC_9_17_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_2_1_LC_9_17_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_2_1_LC_9_17_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_RNIN79A_2_1_LC_9_17_1  (
            .in0(N__8530),
            .in1(N__10663),
            .in2(N__8570),
            .in3(N__10571),
            .lcout(\DUT.fifo_tx_inst.rFifoData_awe3 ),
            .ltout(\DUT.fifo_tx_inst.rFifoData_awe3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIJLJC_1_LC_9_17_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIJLJC_1_LC_9_17_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIJLJC_1_LC_9_17_2 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_RNIJLJC_1_LC_9_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7046),
            .in3(N__12061),
            .lcout(\DUT.fifo_tx_inst.un1_i11_i ),
            .ltout(\DUT.fifo_tx_inst.un1_i11_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_1_LC_9_17_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_1_LC_9_17_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rWritePtr_1_LC_9_17_3 .LUT_INIT=16'b0000011100001000;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_1_LC_9_17_3  (
            .in0(N__8486),
            .in1(N__8569),
            .in2(N__7037),
            .in3(N__8531),
            .lcout(\DUT.fifo_tx_inst.rWritePtrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13039),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNI323D2_2_LC_9_17_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNI323D2_2_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNI323D2_2_LC_9_17_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNI323D2_2_LC_9_17_4  (
            .in0(N__7029),
            .in1(N__6941),
            .in2(N__6889),
            .in3(N__6870),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_8_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNIV8RM6_0_LC_9_17_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNIV8RM6_0_LC_9_17_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNIV8RM6_0_LC_9_17_5 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNIV8RM6_0_LC_9_17_5  (
            .in0(N__6800),
            .in1(N__6719),
            .in2(N__6605),
            .in3(N__6602),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNIG3R3E_2_LC_9_17_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNIG3R3E_2_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNIG3R3E_2_LC_9_17_6 .LUT_INIT=16'b1000000000100000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNIG3R3E_2_LC_9_17_6  (
            .in0(N__6596),
            .in1(N__6587),
            .in2(N__6578),
            .in3(N__7926),
            .lcout(\DUT.uart_inst0.rx_bits_remaining_2_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_0_LC_9_18_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_0_LC_9_18_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_0_LC_9_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_0_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7351),
            .lcout(\DUT.wRxByte_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13034),
            .ce(N__7160),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_1_LC_9_18_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_1_LC_9_18_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_1_LC_9_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_1_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7303),
            .lcout(\DUT.wRxByte_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13034),
            .ce(N__7160),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_2_LC_9_18_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_2_LC_9_18_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_2_LC_9_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_2_LC_9_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7787),
            .lcout(\DUT.wRxByte_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13034),
            .ce(N__7160),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_3_LC_9_18_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_3_LC_9_18_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_3_LC_9_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_3_LC_9_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7731),
            .lcout(\DUT.wRxByte_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13034),
            .ce(N__7160),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_4_LC_9_18_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_4_LC_9_18_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_4_LC_9_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_4_LC_9_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7680),
            .lcout(\DUT.wRxByte_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13034),
            .ce(N__7160),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_5_LC_9_18_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_5_LC_9_18_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_5_LC_9_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_5_LC_9_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7628),
            .lcout(\DUT.wRxByte_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13034),
            .ce(N__7160),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_6_LC_9_18_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_6_LC_9_18_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_6_LC_9_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_6_LC_9_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10469),
            .lcout(\DUT.wRxByte_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13034),
            .ce(N__7160),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_7_LC_9_18_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_7_LC_9_18_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_7_LC_9_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_7_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10111),
            .lcout(\DUT.wRxByte_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13034),
            .ce(N__7160),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIPTFQ1_0_LC_9_19_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIPTFQ1_0_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIPTFQ1_0_LC_9_19_0 .LUT_INIT=16'b1101110110011001;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNIPTFQ1_0_LC_9_19_0  (
            .in0(N__7138),
            .in1(N__10647),
            .in2(_gnd_net_),
            .in3(N__8221),
            .lcout(\DUT.fifo_rx_inst.N_87 ),
            .ltout(\DUT.fifo_rx_inst.N_87_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_9_19_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_9_19_1 .LUT_INIT=16'b0000001100001111;
    LogicCell40 \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_9_19_1  (
            .in0(N__7071),
            .in1(N__7139),
            .in2(N__7151),
            .in3(N__7265),
            .lcout(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_0_LC_9_19_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_0_LC_9_19_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoCount_0_LC_9_19_2 .LUT_INIT=16'b1111100000000111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_0_LC_9_19_2  (
            .in0(N__7266),
            .in1(N__7140),
            .in2(N__7088),
            .in3(N__7070),
            .lcout(\DUT.fifo_rx_inst.rFifoCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13028),
            .ce(),
            .sr(N__10525));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_0_LC_9_19_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_0_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_0_LC_9_19_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_0_LC_9_19_4  (
            .in0(N__7264),
            .in1(N__7228),
            .in2(_gnd_net_),
            .in3(N__7068),
            .lcout(\DUT.fifo_rx_inst.N_92 ),
            .ltout(\DUT.fifo_rx_inst.N_92_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rReadPtr_RNI8B9Q1_0_LC_9_19_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rReadPtr_RNI8B9Q1_0_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rReadPtr_RNI8B9Q1_0_LC_9_19_5 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \DUT.fifo_rx_inst.rReadPtr_RNI8B9Q1_0_LC_9_19_5  (
            .in0(N__10648),
            .in1(_gnd_net_),
            .in2(N__7079),
            .in3(N__8163),
            .lcout(\DUT.fifo_rx_inst.CO0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rRxRead_LC_9_19_7.C_ON=1'b0;
    defparam rRxRead_LC_9_19_7.SEQ_MODE=4'b1000;
    defparam rRxRead_LC_9_19_7.LUT_INIT=16'b1111111111101110;
    LogicCell40 rRxRead_LC_9_19_7 (
            .in0(N__7069),
            .in1(N__7267),
            .in2(_gnd_net_),
            .in3(N__7234),
            .lcout(rRxReadZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13028),
            .ce(),
            .sr(N__10525));
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_LC_9_20_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_LC_9_20_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_LC_9_20_0  (
            .in0(N__8575),
            .in1(N__8534),
            .in2(_gnd_net_),
            .in3(N__8476),
            .lcout(\DUT.fifo_tx_inst.rFifoData_awe2 ),
            .ltout(\DUT.fifo_tx_inst.rFifoData_awe2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_LC_9_20_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_LC_9_20_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_LC_9_20_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_2_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7193),
            .in3(N__7181),
            .lcout(\DUT.fifo_tx_inst.rFifoDataro_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13023),
            .ce(),
            .sr(N__10524));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_3_LC_9_20_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_3_LC_9_20_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_3_LC_9_20_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_3_LC_9_20_2  (
            .in0(N__7190),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12523),
            .lcout(\DUT.fifo_tx_inst.rFifoDataro_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13023),
            .ce(),
            .sr(N__10524));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_9_20_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_9_20_3 .LUT_INIT=16'b0010111101111111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_9_20_3  (
            .in0(N__10901),
            .in1(N__7189),
            .in2(N__10852),
            .in3(N__7180),
            .lcout(\DUT.rFifoDataror_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_1_LC_9_20_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_1_LC_9_20_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_1_LC_9_20_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_1_LC_9_20_5  (
            .in0(_gnd_net_),
            .in1(N__8437),
            .in2(_gnd_net_),
            .in3(N__12861),
            .lcout(\DUT.fifo_tx_inst.rFifoDataro_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13023),
            .ce(),
            .sr(N__10524));
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_1_LC_9_20_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_1_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_1_LC_9_20_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_1_LC_9_20_6  (
            .in0(N__8574),
            .in1(N__8533),
            .in2(_gnd_net_),
            .in3(N__8475),
            .lcout(\DUT.fifo_tx_inst.rFifoData_awe0 ),
            .ltout(\DUT.fifo_tx_inst.rFifoData_awe0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_LC_9_20_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_LC_9_20_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_LC_9_20_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_0_LC_9_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7172),
            .in3(N__8450),
            .lcout(\DUT.fifo_tx_inst.rFifoDataro_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13023),
            .ce(),
            .sr(N__10524));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNI0AQO1_LC_9_21_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNI0AQO1_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNI0AQO1_LC_9_21_0 .LUT_INIT=16'b1111001011110111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_0_RNI0AQO1_LC_9_21_0  (
            .in0(N__8161),
            .in1(N__7495),
            .in2(N__8968),
            .in3(N__7168),
            .lcout(\DUT.fifo_rx_inst.rTxByte_42_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_LC_9_21_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_LC_9_21_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_LC_9_21_1 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_0_LC_9_21_1  (
            .in0(N__7169),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10424),
            .lcout(\DUT.fifo_rx_inst.rFifoDataro_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13017),
            .ce(),
            .sr(N__10523));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_1_LC_9_21_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_1_LC_9_21_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_1_LC_9_21_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_1_LC_9_21_2  (
            .in0(_gnd_net_),
            .in1(N__7507),
            .in2(_gnd_net_),
            .in3(N__7496),
            .lcout(\DUT.fifo_rx_inst.rFifoDataro_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13017),
            .ce(),
            .sr(N__10523));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_3_LC_9_21_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_3_LC_9_21_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_3_LC_9_21_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_3_LC_9_21_3  (
            .in0(N__7469),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7585),
            .lcout(\DUT.fifo_rx_inst.rFifoDataro_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13017),
            .ce(),
            .sr(N__10523));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_LC_9_21_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_LC_9_21_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_LC_9_21_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_2_LC_9_21_4  (
            .in0(_gnd_net_),
            .in1(N__7459),
            .in2(_gnd_net_),
            .in3(N__7480),
            .lcout(\DUT.fifo_rx_inst.rFifoDataro_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13017),
            .ce(),
            .sr(N__10523));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_9_21_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_9_21_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_9_21_5 .LUT_INIT=16'b0111011100111111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_9_21_5  (
            .in0(N__7468),
            .in1(N__8946),
            .in2(N__7460),
            .in3(N__8162),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rTxByte_42_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNIHJV05_LC_9_21_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNIHJV05_LC_9_21_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNIHJV05_LC_9_21_6 .LUT_INIT=16'b0101010111010101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_0_RNIHJV05_LC_9_21_6  (
            .in0(N__12072),
            .in1(N__7448),
            .in2(N__7442),
            .in3(N__8228),
            .lcout(rFifoDatarff_0_RNIHJV05),
            .ltout(rFifoDatarff_0_RNIHJV05_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI250E6_0_LC_9_21_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI250E6_0_LC_9_21_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI250E6_0_LC_9_21_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNI250E6_0_LC_9_21_7  (
            .in0(N__7439),
            .in1(_gnd_net_),
            .in2(N__7430),
            .in3(_gnd_net_),
            .lcout(N_92_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_9_22_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_9_22_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_9_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_9_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7426),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13012),
            .ce(N__7589),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_9_22_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_9_22_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_9_22_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_9_22_1  (
            .in0(N__7370),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13012),
            .ce(N__7589),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_9_22_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_9_22_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_9_22_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_9_22_2  (
            .in0(N__7319),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13012),
            .ce(N__7589),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_9_22_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_9_22_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_9_22_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_9_22_3  (
            .in0(N__7802),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13012),
            .ce(N__7589),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_9_22_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_9_22_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_9_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_9_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7760),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13012),
            .ce(N__7589),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_9_22_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_9_22_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_9_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_9_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7709),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13012),
            .ce(N__7589),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_9_22_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_9_22_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_9_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_9_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7653),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13012),
            .ce(N__7589),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_9_22_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_9_22_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_9_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_9_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10490),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13012),
            .ce(N__7589),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_9_23_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_9_23_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_9_23_0 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_9_23_0  (
            .in0(N__8192),
            .in1(N__10451),
            .in2(N__9026),
            .in3(N__7562),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ft2232h_inst.rFifoState_1_LC_10_12_5 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rFifoState_1_LC_10_12_5 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rFifoState_1_LC_10_12_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_inst.ft2232h_inst.rFifoState_1_LC_10_12_5  (
            .in0(N__11121),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11010),
            .lcout(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13051),
            .ce(),
            .sr(N__10529));
    defparam \fifo_inst.ft2232h_inst.rRx_n_LC_10_12_6 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rRx_n_LC_10_12_6 .SEQ_MODE=4'b1001;
    defparam \fifo_inst.ft2232h_inst.rRx_n_LC_10_12_6 .LUT_INIT=16'b1111110101110000;
    LogicCell40 \fifo_inst.ft2232h_inst.rRx_n_LC_10_12_6  (
            .in0(N__11011),
            .in1(N__11122),
            .in2(N__8819),
            .in3(N__7522),
            .lcout(P1A3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13051),
            .ce(),
            .sr(N__10529));
    defparam \fifo_inst.ft2232h_inst.rFifoState_2_LC_10_12_7 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rFifoState_2_LC_10_12_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rFifoState_2_LC_10_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.ft2232h_inst.rFifoState_2_LC_10_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7949),
            .lcout(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13051),
            .ce(),
            .sr(N__10529));
    defparam \DUT.uart_inst0.rx_clk_divider_RNI6B671_5_LC_10_13_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI6B671_5_LC_10_13_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI6B671_5_LC_10_13_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNI6B671_5_LC_10_13_0  (
            .in0(N__9090),
            .in1(N__9114),
            .in2(N__9065),
            .in3(N__9141),
            .lcout(\DUT.uart_inst0.un2_rx_clk_divider_a_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_7_LC_10_13_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_7_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_7_LC_10_13_1 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_7_LC_10_13_1  (
            .in0(N__9092),
            .in1(N__9074),
            .in2(_gnd_net_),
            .in3(N__9591),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13046),
            .ce(N__11976),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_5_LC_10_13_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_5_LC_10_13_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_5_LC_10_13_2 .LUT_INIT=16'b1111111110011111;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_5_LC_10_13_2  (
            .in0(N__9128),
            .in1(N__9142),
            .in2(N__9613),
            .in3(N__7921),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13046),
            .ce(N__11976),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_6_LC_10_13_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_6_LC_10_13_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_6_LC_10_13_3 .LUT_INIT=16'b1111101110111111;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_6_LC_10_13_3  (
            .in0(N__7922),
            .in1(N__9599),
            .in2(N__9119),
            .in3(N__9101),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13046),
            .ce(N__11976),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_8_LC_10_13_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_8_LC_10_13_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_8_LC_10_13_4 .LUT_INIT=16'b1010000001010000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_8_LC_10_13_4  (
            .in0(N__9063),
            .in1(_gnd_net_),
            .in2(N__9612),
            .in3(N__9047),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13046),
            .ce(N__11976),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_11_LC_10_13_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_11_LC_10_13_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_11_LC_10_13_5 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_11_LC_10_13_5  (
            .in0(N__9359),
            .in1(N__9341),
            .in2(_gnd_net_),
            .in3(N__9590),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13046),
            .ce(N__11976),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIB99J_10_LC_10_13_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIB99J_10_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIB99J_10_LC_10_13_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIB99J_10_LC_10_13_6  (
            .in0(N__9357),
            .in1(N__9384),
            .in2(N__9416),
            .in3(N__9676),
            .lcout(\DUT.uart_inst0.un2_rx_clk_divider_a_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_9_LC_10_13_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_9_LC_10_13_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_9_LC_10_13_7 .LUT_INIT=16'b1100001100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_9_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(N__9414),
            .in2(N__9398),
            .in3(N__9595),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13046),
            .ce(N__11976),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNI3ALC_17_LC_10_14_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI3ALC_17_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI3ALC_17_LC_10_14_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNI3ALC_17_LC_10_14_0  (
            .in0(N__9276),
            .in1(N__9303),
            .in2(N__9698),
            .in3(N__9327),
            .lcout(\DUT.uart_inst0.un2_rx_clk_divider_a_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_13_LC_10_14_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_13_LC_10_14_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_13_LC_10_14_1 .LUT_INIT=16'b1010000001010000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_13_LC_10_14_1  (
            .in0(N__9328),
            .in1(_gnd_net_),
            .in2(N__9614),
            .in3(N__9314),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13042),
            .ce(N__11978),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_14_LC_10_14_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_14_LC_10_14_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_14_LC_10_14_2 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_14_LC_10_14_2  (
            .in0(N__9305),
            .in1(N__9287),
            .in2(_gnd_net_),
            .in3(N__9605),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13042),
            .ce(N__11978),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_15_LC_10_14_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_15_LC_10_14_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_15_LC_10_14_3 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_15_LC_10_14_3  (
            .in0(N__9606),
            .in1(N__9263),
            .in2(_gnd_net_),
            .in3(N__9277),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13042),
            .ce(N__11978),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_0_LC_10_14_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_0_LC_10_14_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_0_LC_10_14_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_0_LC_10_14_4  (
            .in0(N__8590),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9600),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13042),
            .ce(N__11978),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIJI4K1_16_LC_10_14_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIJI4K1_16_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIJI4K1_16_LC_10_14_5 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIJI4K1_16_LC_10_14_5  (
            .in0(N__9252),
            .in1(N__8589),
            .in2(_gnd_net_),
            .in3(N__7964),
            .lcout(\DUT.uart_inst0.un2_rx_clk_divider_a_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_16_LC_10_14_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_16_LC_10_14_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_16_LC_10_14_6 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_16_LC_10_14_6  (
            .in0(N__9254),
            .in1(N__9236),
            .in2(_gnd_net_),
            .in3(N__9607),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13042),
            .ce(N__11978),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_10_LC_10_14_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_10_LC_10_14_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_10_LC_10_14_7 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_10_LC_10_14_7  (
            .in0(N__9601),
            .in1(N__9368),
            .in2(_gnd_net_),
            .in3(N__9386),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13042),
            .ce(N__11978),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_10_15_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_10_15_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_10_15_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_10_15_0  (
            .in0(N__9734),
            .in1(N__9782),
            .in2(_gnd_net_),
            .in3(N__9856),
            .lcout(),
            .ltout(\DUT.uart_inst0.un1_N_5_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_3_LC_10_15_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_3_LC_10_15_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_bits_remaining_3_LC_10_15_1 .LUT_INIT=16'b1101110101111101;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_3_LC_10_15_1  (
            .in0(N__7970),
            .in1(N__9897),
            .in2(N__7952),
            .in3(N__9752),
            .lcout(\DUT.uart_inst0.tx_bits_remainingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13040),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_5_3_LC_10_15_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_5_3_LC_10_15_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_5_3_LC_10_15_2 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_5_3_LC_10_15_2  (
            .in0(N__11414),
            .in1(N__11834),
            .in2(N__11593),
            .in3(N__11924),
            .lcout(),
            .ltout(\DUT.uart_inst0.g0_i_o6_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_10_15_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_10_15_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_10_15_3 .LUT_INIT=16'b0000000011111100;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(N__7979),
            .in2(N__7982),
            .in3(N__11885),
            .lcout(\DUT.uart_inst0.g0_i_a6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_6_3_LC_10_15_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_6_3_LC_10_15_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_6_3_LC_10_15_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_6_3_LC_10_15_4  (
            .in0(N__9732),
            .in1(N__9780),
            .in2(N__9901),
            .in3(N__9852),
            .lcout(\DUT.uart_inst0.g0_i_o6_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_4_2_LC_10_15_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_4_2_LC_10_15_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_4_2_LC_10_15_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_4_2_LC_10_15_5  (
            .in0(N__9781),
            .in1(N__9896),
            .in2(N__9857),
            .in3(N__9733),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_139_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_2_LC_10_15_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_2_LC_10_15_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_2_LC_10_15_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_0_2_LC_10_15_6  (
            .in0(N__11415),
            .in1(N__11536),
            .in2(N__7973),
            .in3(N__11777),
            .lcout(\DUT.uart_inst0.g0_11_a4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_1_3_LC_10_15_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_1_3_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_1_3_LC_10_15_7 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNO_1_3_LC_10_15_7  (
            .in0(N__11537),
            .in1(N__11416),
            .in2(N__12073),
            .in3(N__11680),
            .lcout(\DUT.uart_inst0.tx_bits_remaining_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_0_LC_10_16_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_0_LC_10_16_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_state_0_LC_10_16_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DUT.uart_inst0.tx_state_0_LC_10_16_0  (
            .in0(N__8123),
            .in1(N__10180),
            .in2(_gnd_net_),
            .in3(N__9424),
            .lcout(\DUT.tx_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13035),
            .ce(),
            .sr(N__10526));
    defparam \DUT.uart_inst0.tx_state_1_LC_10_16_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_1_LC_10_16_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_state_1_LC_10_16_1 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \DUT.uart_inst0.tx_state_1_LC_10_16_1  (
            .in0(N__9425),
            .in1(N__11408),
            .in2(N__10184),
            .in3(N__10235),
            .lcout(\DUT.uart_inst0.tx_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13035),
            .ce(),
            .sr(N__10526));
    defparam \DUT.uart_inst0.tx_data_0_LC_10_17_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_0_LC_10_17_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_0_LC_10_17_0 .LUT_INIT=16'b1100000011100010;
    LogicCell40 \DUT.uart_inst0.tx_data_0_LC_10_17_0  (
            .in0(N__10388),
            .in1(N__11545),
            .in2(N__8060),
            .in3(N__8389),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13030),
            .ce(N__8002),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNINQKO8_0_0_LC_10_17_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNINQKO8_0_0_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNINQKO8_0_0_LC_10_17_1 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \DUT.uart_inst0.tx_state_RNINQKO8_0_0_LC_10_17_1  (
            .in0(N__9801),
            .in1(N__9825),
            .in2(N__11595),
            .in3(N__10232),
            .lcout(\DUT.uart_inst0.N_22_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_1_LC_10_17_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_1_LC_10_17_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_1_LC_10_17_2 .LUT_INIT=16'b1100111000000010;
    LogicCell40 \DUT.uart_inst0.tx_data_1_LC_10_17_2  (
            .in0(N__10355),
            .in1(N__11548),
            .in2(N__8396),
            .in3(N__8051),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13030),
            .ce(N__8002),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_2_LC_10_17_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_2_LC_10_17_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_2_LC_10_17_3 .LUT_INIT=16'b1100010111000000;
    LogicCell40 \DUT.uart_inst0.tx_data_2_LC_10_17_3  (
            .in0(N__8387),
            .in1(N__8045),
            .in2(N__11596),
            .in3(N__8099),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13030),
            .ce(N__8002),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_3_LC_10_17_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_3_LC_10_17_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_3_LC_10_17_4 .LUT_INIT=16'b1100000011100010;
    LogicCell40 \DUT.uart_inst0.tx_data_3_LC_10_17_4  (
            .in0(N__8069),
            .in1(N__11546),
            .in2(N__8039),
            .in3(N__8390),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13030),
            .ce(N__8002),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_4_LC_10_17_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_4_LC_10_17_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_4_LC_10_17_5 .LUT_INIT=16'b1100010111000000;
    LogicCell40 \DUT.uart_inst0.tx_data_4_LC_10_17_5  (
            .in0(N__8388),
            .in1(N__8030),
            .in2(N__11597),
            .in3(N__10328),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13030),
            .ce(N__8002),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_5_LC_10_17_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_5_LC_10_17_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_5_LC_10_17_6 .LUT_INIT=16'b1100000011100010;
    LogicCell40 \DUT.uart_inst0.tx_data_5_LC_10_17_6  (
            .in0(N__10934),
            .in1(N__11547),
            .in2(N__8021),
            .in3(N__8391),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13030),
            .ce(N__8002),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_6_LC_10_17_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_6_LC_10_17_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_6_LC_10_17_7 .LUT_INIT=16'b1100000011001010;
    LogicCell40 \DUT.uart_inst0.tx_data_6_LC_10_17_7  (
            .in0(N__10748),
            .in1(N__8012),
            .in2(N__11598),
            .in3(N__8395),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13030),
            .ce(N__8002),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_7_LC_10_18_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_7_LC_10_18_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_7_LC_10_18_0 .LUT_INIT=16'b0000001000100010;
    LogicCell40 \DUT.uart_inst0.tx_data_7_LC_10_18_0  (
            .in0(N__10280),
            .in1(N__11576),
            .in2(N__8423),
            .in3(N__8411),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13025),
            .ce(N__8003),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_5_LC_10_18_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_5_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_5_LC_10_18_1 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_1_5_LC_10_18_1  (
            .in0(N__11412),
            .in1(_gnd_net_),
            .in2(N__11603),
            .in3(N__11664),
            .lcout(\DUT.uart_inst0.N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_3_2_LC_10_18_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_3_2_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_3_2_LC_10_18_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_3_2_LC_10_18_2  (
            .in0(N__11665),
            .in1(N__11566),
            .in2(_gnd_net_),
            .in3(N__11413),
            .lcout(\DUT.uart_inst0.N_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNICU6U_1_LC_10_18_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNICU6U_1_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNICU6U_1_LC_10_18_3 .LUT_INIT=16'b1111101011111111;
    LogicCell40 \DUT.uart_inst0.tx_state_RNICU6U_1_LC_10_18_3  (
            .in0(N__11410),
            .in1(_gnd_net_),
            .in2(N__11601),
            .in3(N__11662),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_79_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNI5PJS2_1_LC_10_18_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNI5PJS2_1_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNI5PJS2_1_LC_10_18_4 .LUT_INIT=16'b1111111101011111;
    LogicCell40 \DUT.uart_inst0.tx_state_RNI5PJS2_1_LC_10_18_4  (
            .in0(N__12063),
            .in1(_gnd_net_),
            .in2(N__8126),
            .in3(N__12227),
            .lcout(\DUT.uart_inst0.N_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNO_0_0_LC_10_18_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNO_0_0_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNO_0_0_LC_10_18_5 .LUT_INIT=16'b1010101010101111;
    LogicCell40 \DUT.uart_inst0.tx_state_RNO_0_0_LC_10_18_5  (
            .in0(N__11411),
            .in1(_gnd_net_),
            .in2(N__11602),
            .in3(N__11663),
            .lcout(\DUT.uart_inst0.tx_state_ns_i_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNI3R8C_1_LC_10_18_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNI3R8C_1_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNI3R8C_1_LC_10_18_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \DUT.uart_inst0.tx_state_RNI3R8C_1_LC_10_18_6  (
            .in0(N__12062),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11409),
            .lcout(\DUT.rTransmitc_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNIBTN81_0_LC_10_18_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNIBTN81_0_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNIBTN81_0_LC_10_18_7 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \DUT.uart_inst0.tx_state_RNIBTN81_0_LC_10_18_7  (
            .in0(N__11565),
            .in1(N__9872),
            .in2(_gnd_net_),
            .in3(N__11661),
            .lcout(\DUT.uart_inst0.N_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_10_19_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_10_19_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_10_19_0  (
            .in0(N__8090),
            .in1(N__10826),
            .in2(N__12461),
            .in3(N__10903),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_10_19_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_10_19_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_10_19_1  (
            .in0(N__10830),
            .in1(N__12095),
            .in2(N__8114),
            .in3(N__8111),
            .lcout(\DUT.rFifoDatarx_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_10_19_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_10_19_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_10_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_10_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12499),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13019),
            .ce(N__13189),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_10_19_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_10_19_3 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_10_19_3  (
            .in0(N__10904),
            .in1(N__12410),
            .in2(N__10853),
            .in3(N__8456),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_10_19_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_10_19_4 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_10_19_4  (
            .in0(N__12086),
            .in1(N__8084),
            .in2(N__8072),
            .in3(N__10831),
            .lcout(\DUT.rFifoDatarx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_10_19_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_10_19_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_10_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_10_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12438),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13019),
            .ce(N__13189),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_RNI86BE_LC_10_19_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_RNI86BE_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_RNI86BE_LC_10_19_6 .LUT_INIT=16'b1100111111011101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_0_RNI86BE_LC_10_19_6  (
            .in0(N__8449),
            .in1(N__10825),
            .in2(N__8438),
            .in3(N__10902),
            .lcout(\DUT.rFifoDataror_1 ),
            .ltout(\DUT.rFifoDataror_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_RNIKCMS_LC_10_19_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_RNIKCMS_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_RNIKCMS_LC_10_19_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_0_RNIKCMS_LC_10_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8414),
            .in3(N__8407),
            .lcout(\DUT.rFifoDataror_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.rTransmit_LC_10_20_0 .C_ON=1'b0;
    defparam \DUT.rTransmit_LC_10_20_0 .SEQ_MODE=4'b1000;
    defparam \DUT.rTransmit_LC_10_20_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \DUT.rTransmit_LC_10_20_0  (
            .in0(N__8492),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11605),
            .lcout(\DUT.rTransmitZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13014),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rReadPtr_1_LC_10_20_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rReadPtr_1_LC_10_20_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rReadPtr_1_LC_10_20_1 .LUT_INIT=16'b0000000001011010;
    LogicCell40 \DUT.fifo_rx_inst.rReadPtr_1_LC_10_20_1  (
            .in0(N__8246),
            .in1(_gnd_net_),
            .in2(N__9003),
            .in3(N__8237),
            .lcout(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13014),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rReadPtr_1_LC_10_20_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rReadPtr_1_LC_10_20_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rReadPtr_1_LC_10_20_2 .LUT_INIT=16'b0000100100001100;
    LogicCell40 \DUT.fifo_tx_inst.rReadPtr_1_LC_10_20_2  (
            .in0(N__10598),
            .in1(N__10851),
            .in2(N__9038),
            .in3(N__10915),
            .lcout(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13014),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rReadPtr_0_LC_10_20_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rReadPtr_0_LC_10_20_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rReadPtr_0_LC_10_20_3 .LUT_INIT=16'b0010001000010001;
    LogicCell40 \DUT.fifo_tx_inst.rReadPtr_0_LC_10_20_3  (
            .in0(N__10914),
            .in1(N__9034),
            .in2(_gnd_net_),
            .in3(N__10597),
            .lcout(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13014),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rReadPtr_RNI4NC92_1_LC_10_20_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rReadPtr_RNI4NC92_1_LC_10_20_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rReadPtr_RNI4NC92_1_LC_10_20_4 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \DUT.fifo_rx_inst.rReadPtr_RNI4NC92_1_LC_10_20_4  (
            .in0(N__8332),
            .in1(N__8964),
            .in2(_gnd_net_),
            .in3(N__8245),
            .lcout(\DUT.fifo_rx_inst.un1_i11_2_i ),
            .ltout(\DUT.fifo_rx_inst.un1_i11_2_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rReadPtr_0_LC_10_20_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rReadPtr_0_LC_10_20_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rReadPtr_0_LC_10_20_5 .LUT_INIT=16'b0000101000000110;
    LogicCell40 \DUT.fifo_rx_inst.rReadPtr_0_LC_10_20_5  (
            .in0(N__8176),
            .in1(N__10654),
            .in2(N__8231),
            .in3(N__8227),
            .lcout(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13014),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_0_1_LC_10_20_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_0_1_LC_10_20_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_0_1_LC_10_20_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_RNIN79A_0_1_LC_10_20_6  (
            .in0(N__8576),
            .in1(N__8532),
            .in2(_gnd_net_),
            .in3(N__8474),
            .lcout(\DUT.fifo_tx_inst.rFifoData_awe1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNI8CH01_1_LC_10_20_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNI8CH01_1_LC_10_20_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNI8CH01_1_LC_10_20_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \DUT.uart_inst0.tx_state_RNI8CH01_1_LC_10_20_7  (
            .in0(N__11604),
            .in1(N__11438),
            .in2(N__12074),
            .in3(N__11660),
            .lcout(\DUT.uart_inst0.N_65_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_10_21_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_10_21_0 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_10_21_0  (
            .in0(N__10555),
            .in1(N__10658),
            .in2(N__10736),
            .in3(N__8501),
            .lcout(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIME2J_0_LC_10_21_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIME2J_0_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIME2J_0_LC_10_21_1 .LUT_INIT=16'b0101010101010111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNIME2J_0_LC_10_21_1  (
            .in0(N__11636),
            .in1(N__10682),
            .in2(N__10734),
            .in3(N__10553),
            .lcout(\DUT.fifo_tx_inst.N_83 ),
            .ltout(\DUT.fifo_tx_inst.N_83_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIDGST_0_LC_10_21_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIDGST_0_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIDGST_0_LC_10_21_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNIDGST_0_LC_10_21_2  (
            .in0(_gnd_net_),
            .in1(N__10655),
            .in2(N__8504),
            .in3(N__11637),
            .lcout(\DUT.fifo_tx_inst.N_88 ),
            .ltout(\DUT.fifo_tx_inst.N_88_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_0_LC_10_21_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_0_LC_10_21_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoCount_0_LC_10_21_3 .LUT_INIT=16'b1111100000000111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_0_LC_10_21_3  (
            .in0(N__10659),
            .in1(N__10557),
            .in2(N__8495),
            .in3(N__10730),
            .lcout(\DUT.rFifoCount_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13008),
            .ce(),
            .sr(N__10522));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIBPFM_1_LC_10_21_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIBPFM_1_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIBPFM_1_LC_10_21_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNIBPFM_1_LC_10_21_4  (
            .in0(N__10684),
            .in1(N__10594),
            .in2(_gnd_net_),
            .in3(N__10657),
            .lcout(\DUT.fifo_tx_inst.rFifoCount_RNIBPFMZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.rTransmit_RNO_0_LC_10_21_5 .C_ON=1'b0;
    defparam \DUT.rTransmit_RNO_0_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \DUT.rTransmit_RNO_0_LC_10_21_5 .LUT_INIT=16'b1010101010101011;
    LogicCell40 \DUT.rTransmit_RNO_0_LC_10_21_5  (
            .in0(N__9830),
            .in1(N__10683),
            .in2(N__10735),
            .in3(N__10556),
            .lcout(\DUT.rTransmitc ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIMBD3_2_LC_10_21_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIMBD3_2_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIMBD3_2_LC_10_21_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNIMBD3_2_LC_10_21_6  (
            .in0(N__10554),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10656),
            .lcout(\DUT.fifo_tx_inst.rWritePtr16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rReadPtr_RNILV421_0_LC_10_21_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rReadPtr_RNILV421_0_LC_10_21_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rReadPtr_RNILV421_0_LC_10_21_7 .LUT_INIT=16'b0111001100110011;
    LogicCell40 \DUT.fifo_tx_inst.rReadPtr_RNILV421_0_LC_10_21_7  (
            .in0(N__10595),
            .in1(N__12071),
            .in2(N__10916),
            .in3(N__10850),
            .lcout(\DUT.fifo_tx_inst.un1_i11_2_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rTxByte_esr_1_LC_10_22_3.C_ON=1'b0;
    defparam rTxByte_esr_1_LC_10_22_3.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_1_LC_10_22_3.LUT_INIT=16'b1000100011110101;
    LogicCell40 rTxByte_esr_1_LC_10_22_3 (
            .in0(N__8976),
            .in1(N__8909),
            .in2(N__8897),
            .in3(N__8888),
            .lcout(rTxByteZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13005),
            .ce(N__8878),
            .sr(N__8851));
    defparam \fifo_inst.ft2232h_inst.rFifoState_4_LC_11_12_0 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rFifoState_4_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rFifoState_4_LC_11_12_0 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \fifo_inst.ft2232h_inst.rFifoState_4_LC_11_12_0  (
            .in0(N__8612),
            .in1(N__8637),
            .in2(_gnd_net_),
            .in3(N__8761),
            .lcout(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13047),
            .ce(),
            .sr(N__10528));
    defparam \fifo_inst.ft2232h_inst.rFifoState_0_LC_11_12_1 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rFifoState_0_LC_11_12_1 .SEQ_MODE=4'b1001;
    defparam \fifo_inst.ft2232h_inst.rFifoState_0_LC_11_12_1 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \fifo_inst.ft2232h_inst.rFifoState_0_LC_11_12_1  (
            .in0(N__8638),
            .in1(N__8815),
            .in2(N__8617),
            .in3(N__10982),
            .lcout(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13047),
            .ce(),
            .sr(N__10528));
    defparam \fifo_inst.ft2232h_inst.rTx_n_LC_11_12_2 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rTx_n_LC_11_12_2 .SEQ_MODE=4'b1001;
    defparam \fifo_inst.ft2232h_inst.rTx_n_LC_11_12_2 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \fifo_inst.ft2232h_inst.rTx_n_LC_11_12_2  (
            .in0(N__8639),
            .in1(N__8762),
            .in2(N__8618),
            .in3(N__8775),
            .lcout(P1A4_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13047),
            .ce(),
            .sr(N__10528));
    defparam \fifo_inst.ft2232h_inst.rFifoState_3_LC_11_12_3 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rFifoState_3_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rFifoState_3_LC_11_12_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \fifo_inst.ft2232h_inst.rFifoState_3_LC_11_12_3  (
            .in0(N__11120),
            .in1(N__11066),
            .in2(_gnd_net_),
            .in3(N__11009),
            .lcout(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13047),
            .ce(),
            .sr(N__10528));
    defparam \fifo_inst.ft2232h_inst.rTxBusReady_LC_11_12_4 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rTxBusReady_LC_11_12_4 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rTxBusReady_LC_11_12_4 .LUT_INIT=16'b1111111101110000;
    LogicCell40 \fifo_inst.ft2232h_inst.rTxBusReady_LC_11_12_4  (
            .in0(N__8613),
            .in1(N__8635),
            .in2(N__8679),
            .in3(N__9911),
            .lcout(rTxBusReady),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13047),
            .ce(),
            .sr(N__10528));
    defparam \fifo_inst.ft2232h_inst.rTxRdEn_LC_11_12_6 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rTxRdEn_LC_11_12_6 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rTxRdEn_LC_11_12_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \fifo_inst.ft2232h_inst.rTxRdEn_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(N__8608),
            .in2(_gnd_net_),
            .in3(N__8636),
            .lcout(\fifo_inst.ft2232h_inst.rTxRdEnZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13047),
            .ce(),
            .sr(N__10528));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_11_13_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_11_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__8591),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_11_13_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_11_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(N__9227),
            .in2(N__12842),
            .in3(N__9194),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_0 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_11_13_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_11_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(N__9647),
            .in2(N__12846),
            .in3(N__9191),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_1 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_2_THRU_LUT4_0_LC_11_13_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_2_THRU_LUT4_0_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_2_THRU_LUT4_0_LC_11_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_2_THRU_LUT4_0_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__9188),
            .in2(N__12843),
            .in3(N__9149),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_2 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_11_13_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_11_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(N__9490),
            .in2(N__12847),
            .in3(N__9146),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_3 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_4_THRU_LUT4_0_LC_11_13_5 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_4_THRU_LUT4_0_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_4_THRU_LUT4_0_LC_11_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_4_THRU_LUT4_0_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(N__9143),
            .in2(N__12844),
            .in3(N__9122),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_4 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_5_THRU_LUT4_0_LC_11_13_6 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_5_THRU_LUT4_0_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_5_THRU_LUT4_0_LC_11_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_5_THRU_LUT4_0_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(N__9118),
            .in2(N__12848),
            .in3(N__9095),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_5 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_11_13_7 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_11_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(N__9091),
            .in2(N__12845),
            .in3(N__9068),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_6 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_11_14_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_11_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(N__9064),
            .in2(N__12817),
            .in3(N__9041),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_11_14_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_11_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(N__9415),
            .in2(N__12814),
            .in3(N__9389),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_8 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_LUT4_0_LC_11_14_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_LUT4_0_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_LUT4_0_LC_11_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_LUT4_0_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(N__9385),
            .in2(N__12818),
            .in3(N__9362),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_9 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_LUT4_0_LC_11_14_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_LUT4_0_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_LUT4_0_LC_11_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_LUT4_0_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(N__9358),
            .in2(N__12811),
            .in3(N__9335),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_10 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_LUT4_0_LC_11_14_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_LUT4_0_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_LUT4_0_LC_11_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_LUT4_0_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(N__9677),
            .in2(N__12815),
            .in3(N__9332),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_11 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_LUT4_0_LC_11_14_5 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_LUT4_0_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_LUT4_0_LC_11_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_LUT4_0_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(N__9329),
            .in2(N__12812),
            .in3(N__9308),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_12 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_LUT4_0_LC_11_14_6 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_LUT4_0_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_LUT4_0_LC_11_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_LUT4_0_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(N__9304),
            .in2(N__12816),
            .in3(N__9281),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_13 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_LUT4_0_LC_11_14_7 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_LUT4_0_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_LUT4_0_LC_11_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_LUT4_0_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(N__9278),
            .in2(N__12813),
            .in3(N__9257),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_14 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_LUT4_0_LC_11_15_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_LUT4_0_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_LUT4_0_LC_11_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_LUT4_0_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(N__9253),
            .in2(N__12763),
            .in3(N__9230),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_17_LC_11_15_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_17_LC_11_15_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_17_LC_11_15_1 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_17_LC_11_15_1  (
            .in0(N__9609),
            .in1(N__9697),
            .in2(_gnd_net_),
            .in3(N__9701),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13036),
            .ce(N__11979),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_12_LC_11_15_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_12_LC_11_15_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_12_LC_11_15_2 .LUT_INIT=16'b1000100001000100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_12_LC_11_15_2  (
            .in0(N__9683),
            .in1(N__9608),
            .in2(_gnd_net_),
            .in3(N__9675),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13036),
            .ce(N__11979),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_2_LC_11_15_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_2_LC_11_15_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_2_LC_11_15_3 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_2_LC_11_15_3  (
            .in0(N__9610),
            .in1(N__9656),
            .in2(_gnd_net_),
            .in3(N__9645),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13036),
            .ce(N__11979),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_4_LC_11_15_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_4_LC_11_15_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_4_LC_11_15_4 .LUT_INIT=16'b1000100001000100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_4_LC_11_15_4  (
            .in0(N__9623),
            .in1(N__9611),
            .in2(_gnd_net_),
            .in3(N__9486),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13036),
            .ce(N__11979),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_RNO_1_LC_11_16_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_RNO_1_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_out_RNO_1_LC_11_16_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \DUT.uart_inst0.tx_out_RNO_1_LC_11_16_0  (
            .in0(N__11407),
            .in1(N__9431),
            .in2(N__11600),
            .in3(N__10234),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_98_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_LC_11_16_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_LC_11_16_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_out_LC_11_16_1 .LUT_INIT=16'b1111101011111000;
    LogicCell40 \DUT.uart_inst0.tx_out_LC_11_16_1  (
            .in0(N__9448),
            .in1(N__9806),
            .in2(N__9464),
            .in3(N__10211),
            .lcout(P1A7_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13031),
            .ce(N__11985),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_RNO_2_LC_11_16_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_RNO_2_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_out_RNO_2_LC_11_16_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.uart_inst0.tx_out_RNO_2_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(N__9873),
            .in2(_gnd_net_),
            .in3(N__10246),
            .lcout(\DUT.uart_inst0.N_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNISP995_0_LC_11_16_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNISP995_0_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNISP995_0_LC_11_16_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \DUT.uart_inst0.tx_state_RNISP995_0_LC_11_16_3  (
            .in0(N__9874),
            .in1(N__11150),
            .in2(N__11594),
            .in3(N__12221),
            .lcout(\DUT.uart_inst0.N_99 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNISP995_0_0_LC_11_16_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNISP995_0_0_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNISP995_0_0_LC_11_16_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \DUT.uart_inst0.tx_state_RNISP995_0_0_LC_11_16_4  (
            .in0(N__12222),
            .in1(N__9875),
            .in2(N__11599),
            .in3(N__11222),
            .lcout(\DUT.uart_inst0.N_100 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNIHH651_0_LC_11_16_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNIHH651_0_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNIHH651_0_LC_11_16_6 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \DUT.uart_inst0.recv_state_RNIHH651_0_LC_11_16_6  (
            .in0(N__10170),
            .in1(N__10040),
            .in2(_gnd_net_),
            .in3(N__9977),
            .lcout(\DUT.uart_inst0.N_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ft2232h_inst.rFifoState_RNIRPB71_0_LC_11_16_7 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rFifoState_RNIRPB71_0_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ft2232h_inst.rFifoState_RNIRPB71_0_LC_11_16_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \fifo_inst.ft2232h_inst.rFifoState_RNIRPB71_0_LC_11_16_7  (
            .in0(N__11061),
            .in1(N__11108),
            .in2(_gnd_net_),
            .in3(N__11015),
            .lcout(\fifo_inst.ft2232h_inst.rFifoStatec_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_3_LC_11_17_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_3_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_3_LC_11_17_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_3_LC_11_17_1  (
            .in0(N__9843),
            .in1(N__9716),
            .in2(N__9902),
            .in3(N__9769),
            .lcout(\DUT.uart_inst0.N_139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_2_LC_11_17_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_2_LC_11_17_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_bits_remaining_2_LC_11_17_2 .LUT_INIT=16'b1100110011001001;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_2_LC_11_17_2  (
            .in0(N__9772),
            .in1(N__9844),
            .in2(N__9731),
            .in3(N__9748),
            .lcout(\DUT.uart_inst0.tx_bits_remainingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13026),
            .ce(),
            .sr(N__10265));
    defparam \DUT.uart_inst0.tx_countdown_RNI3MLP6_1_LC_11_17_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNI3MLP6_1_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNI3MLP6_1_LC_11_17_3 .LUT_INIT=16'b0011001110101010;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNI3MLP6_1_LC_11_17_3  (
            .in0(N__11221),
            .in1(N__11149),
            .in2(_gnd_net_),
            .in3(N__12199),
            .lcout(\DUT.uart_inst0.N_85 ),
            .ltout(\DUT.uart_inst0.N_85_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNINQKO8_0_LC_11_17_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNINQKO8_0_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNINQKO8_0_LC_11_17_4 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \DUT.uart_inst0.tx_state_RNINQKO8_0_LC_11_17_4  (
            .in0(N__11541),
            .in1(N__9829),
            .in2(N__9809),
            .in3(N__9802),
            .lcout(\DUT.uart_inst0.N_22 ),
            .ltout(\DUT.uart_inst0.N_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_0_LC_11_17_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_0_LC_11_17_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_bits_remaining_0_LC_11_17_5 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_0_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9785),
            .in3(N__9770),
            .lcout(\DUT.uart_inst0.tx_bits_remainingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13026),
            .ce(),
            .sr(N__10265));
    defparam \DUT.uart_inst0.tx_bits_remaining_1_LC_11_17_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_1_LC_11_17_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_bits_remaining_1_LC_11_17_6 .LUT_INIT=16'b1111000010100101;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_1_LC_11_17_6  (
            .in0(N__9771),
            .in1(_gnd_net_),
            .in2(N__9730),
            .in3(N__9747),
            .lcout(\DUT.uart_inst0.tx_bits_remainingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13026),
            .ce(),
            .sr(N__10265));
    defparam \DUT.uart_inst0.tx_out_RNO_0_LC_11_17_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_RNO_0_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_out_RNO_0_LC_11_17_7 .LUT_INIT=16'b1110111011100100;
    LogicCell40 \DUT.uart_inst0.tx_out_RNO_0_LC_11_17_7  (
            .in0(N__11564),
            .in1(N__11406),
            .in2(N__10250),
            .in3(N__10233),
            .lcout(\DUT.uart_inst0.N_89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_11_18_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_11_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(N__11240),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_1_LC_11_18_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_1_LC_11_18_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_1_LC_11_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_1_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(N__11252),
            .in2(N__12759),
            .in3(N__10205),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_1 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_0 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_1 ),
            .clk(N__13020),
            .ce(),
            .sr(N__11268));
    defparam \DUT.uart_inst0.tx_clk_divider_2_LC_11_18_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_2_LC_11_18_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_2_LC_11_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_2_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(N__12350),
            .in2(N__12741),
            .in3(N__10202),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_2 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_1 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_2 ),
            .clk(N__13020),
            .ce(),
            .sr(N__11268));
    defparam \DUT.uart_inst0.tx_clk_divider_3_LC_11_18_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_3_LC_11_18_3 .SEQ_MODE=4'b1001;
    defparam \DUT.uart_inst0.tx_clk_divider_3_LC_11_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_3_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(N__12311),
            .in2(N__12760),
            .in3(N__10199),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_3 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_2 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_3 ),
            .clk(N__13020),
            .ce(),
            .sr(N__11268));
    defparam \DUT.uart_inst0.tx_clk_divider_4_LC_11_18_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_4_LC_11_18_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_4_LC_11_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_4_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(N__12338),
            .in2(N__12742),
            .in3(N__10196),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_4 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_3 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_4 ),
            .clk(N__13020),
            .ce(),
            .sr(N__11268));
    defparam \DUT.uart_inst0.tx_clk_divider_5_LC_11_18_5 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_5_LC_11_18_5 .SEQ_MODE=4'b1001;
    defparam \DUT.uart_inst0.tx_clk_divider_5_LC_11_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_5_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(N__12325),
            .in2(N__12761),
            .in3(N__10193),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_5 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_4 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_5 ),
            .clk(N__13020),
            .ce(),
            .sr(N__11268));
    defparam \DUT.uart_inst0.tx_clk_divider_6_LC_11_18_6 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_6_LC_11_18_6 .SEQ_MODE=4'b1001;
    defparam \DUT.uart_inst0.tx_clk_divider_6_LC_11_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_6_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(N__12260),
            .in2(N__12743),
            .in3(N__10190),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_6 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_5 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_6 ),
            .clk(N__13020),
            .ce(),
            .sr(N__11268));
    defparam \DUT.uart_inst0.tx_clk_divider_7_LC_11_18_7 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_7_LC_11_18_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_7_LC_11_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_7_LC_11_18_7  (
            .in0(_gnd_net_),
            .in1(N__12287),
            .in2(N__12762),
            .in3(N__10187),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_7 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_6 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_7 ),
            .clk(N__13020),
            .ce(),
            .sr(N__11268));
    defparam \DUT.uart_inst0.tx_clk_divider_8_LC_11_19_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_8_LC_11_19_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_8_LC_11_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_8_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(N__11288),
            .in2(N__12758),
            .in3(N__10310),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_8 ),
            .ltout(),
            .carryin(bfn_11_19_0_),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_8 ),
            .clk(N__13015),
            .ce(),
            .sr(N__11272));
    defparam \DUT.uart_inst0.tx_clk_divider_9_LC_11_19_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_9_LC_11_19_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_9_LC_11_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_9_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(N__12702),
            .in2(N__11333),
            .in3(N__10307),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_9 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_8 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_9 ),
            .clk(N__13015),
            .ce(),
            .sr(N__11272));
    defparam \DUT.uart_inst0.tx_clk_divider_10_LC_11_19_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_10_LC_11_19_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_10_LC_11_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_10_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(N__11318),
            .in2(N__12756),
            .in3(N__10304),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_10 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_9 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_10 ),
            .clk(N__13015),
            .ce(),
            .sr(N__11272));
    defparam \DUT.uart_inst0.tx_clk_divider_11_LC_11_19_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_11_LC_11_19_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_11_LC_11_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_11_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(N__12695),
            .in2(N__11306),
            .in3(N__10301),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_11 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_10 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_11 ),
            .clk(N__13015),
            .ce(),
            .sr(N__11272));
    defparam \DUT.uart_inst0.tx_clk_divider_12_LC_11_19_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_12_LC_11_19_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_12_LC_11_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_12_LC_11_19_4  (
            .in0(_gnd_net_),
            .in1(N__12299),
            .in2(N__12757),
            .in3(N__10298),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_12 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_11 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_12 ),
            .clk(N__13015),
            .ce(),
            .sr(N__11272));
    defparam \DUT.uart_inst0.tx_clk_divider_13_LC_11_19_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_13_LC_11_19_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_13_LC_11_19_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_13_LC_11_19_5  (
            .in0(_gnd_net_),
            .in1(N__12274),
            .in2(_gnd_net_),
            .in3(N__10295),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13015),
            .ce(),
            .sr(N__11272));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_11_20_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_11_20_0 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_11_20_0  (
            .in0(N__10907),
            .in1(N__13283),
            .in2(N__10855),
            .in3(N__10271),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_11_20_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_11_20_1 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_11_20_1  (
            .in0(N__10292),
            .in1(N__12533),
            .in2(N__10283),
            .in3(N__10841),
            .lcout(\DUT.rFifoDatarx_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_11_20_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_11_20_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_11_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_11_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13320),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13009),
            .ce(N__13190),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_11_20_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_11_20_3 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_11_20_3  (
            .in0(N__10376),
            .in1(N__10832),
            .in2(N__13067),
            .in3(N__10905),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_11_20_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_11_20_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_11_20_4  (
            .in0(N__10839),
            .in1(N__12107),
            .in2(N__10403),
            .in3(N__10400),
            .lcout(\DUT.rFifoDatarxZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_11_20_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_11_20_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_11_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_11_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13098),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13009),
            .ce(N__13190),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_11_20_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_11_20_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_11_20_6 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_11_20_6  (
            .in0(N__10906),
            .in1(N__12506),
            .in2(N__10854),
            .in3(N__13235),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_11_20_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_11_20_7 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_11_20_7  (
            .in0(N__12101),
            .in1(N__10370),
            .in2(N__10358),
            .in3(N__10840),
            .lcout(\DUT.rFifoDatarx_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_11_21_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_11_21_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_11_21_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_11_21_0  (
            .in0(N__10316),
            .in1(N__10842),
            .in2(N__12368),
            .in3(N__10908),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_11_21_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_11_21_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_11_21_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_11_21_1  (
            .in0(N__10847),
            .in1(N__12569),
            .in2(N__10343),
            .in3(N__10340),
            .lcout(\DUT.rFifoDatarx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_11_21_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_11_21_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_11_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_11_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12390),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13006),
            .ce(N__13187),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_11_21_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_11_21_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_11_21_3 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_11_21_3  (
            .in0(N__10909),
            .in1(N__13115),
            .in2(N__10856),
            .in3(N__10922),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_11_21_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_11_21_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_11_21_4 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_11_21_4  (
            .in0(N__12557),
            .in1(N__10949),
            .in2(N__10937),
            .in3(N__10848),
            .lcout(\DUT.rFifoDatarx_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_11_21_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_11_21_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_11_21_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_11_21_5  (
            .in0(N__13140),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13006),
            .ce(N__13187),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_11_21_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_11_21_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_11_21_6 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_11_21_6  (
            .in0(N__13196),
            .in1(N__10846),
            .in2(N__12359),
            .in3(N__10910),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_11_21_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_11_21_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_11_21_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_11_21_7  (
            .in0(N__10849),
            .in1(N__12545),
            .in2(N__10763),
            .in3(N__10760),
            .lcout(\DUT.rFifoDatarx_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_11_22_0 .C_ON=1'b1;
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_11_22_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_11_22_0  (
            .in0(_gnd_net_),
            .in1(N__10729),
            .in2(N__10703),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_22_0_),
            .carryout(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_1_LC_11_22_1 .C_ON=1'b1;
    defparam \DUT.fifo_tx_inst.rFifoCount_1_LC_11_22_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoCount_1_LC_11_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_1_LC_11_22_1  (
            .in0(_gnd_net_),
            .in1(N__10685),
            .in2(N__10694),
            .in3(N__10667),
            .lcout(\DUT.rFifoCount_1 ),
            .ltout(),
            .carryin(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0 ),
            .carryout(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1 ),
            .clk(N__13003),
            .ce(),
            .sr(N__10521));
    defparam \DUT.fifo_tx_inst.rFifoCount_2_LC_11_22_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_2_LC_11_22_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoCount_2_LC_11_22_2 .LUT_INIT=16'b0001111011100001;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_2_LC_11_22_2  (
            .in0(N__10664),
            .in1(N__10596),
            .in2(N__10567),
            .in3(N__10574),
            .lcout(\DUT.rFifoCount_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13003),
            .ce(),
            .sr(N__10521));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_11_23_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_11_23_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_11_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_11_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10496),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13001),
            .ce(N__10442),
            .sr(_gnd_net_));
    defparam \fifo_inst.ft2232h_inst.rFifoState_RNO_0_0_LC_12_12_1 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rFifoState_RNO_0_0_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ft2232h_inst.rFifoState_RNO_0_0_LC_12_12_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \fifo_inst.ft2232h_inst.rFifoState_RNO_0_0_LC_12_12_1  (
            .in0(N__11123),
            .in1(N__11065),
            .in2(_gnd_net_),
            .in3(N__11005),
            .lcout(\fifo_inst.ft2232h_inst.N_101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_7_3_LC_12_15_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_7_3_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_7_3_LC_12_15_0 .LUT_INIT=16'b0101010101000100;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_7_3_LC_12_15_0  (
            .in0(N__11882),
            .in1(N__11719),
            .in2(_gnd_net_),
            .in3(N__11765),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_4_3_LC_12_15_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_4_3_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_4_3_LC_12_15_1 .LUT_INIT=16'b1111000111110000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_4_3_LC_12_15_1  (
            .in0(N__11609),
            .in1(N__11431),
            .in2(N__10976),
            .in3(N__11687),
            .lcout(),
            .ltout(\DUT.uart_inst0.g0_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_12_15_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_12_15_2 .LUT_INIT=16'b1111000011110010;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_12_15_2  (
            .in0(N__12170),
            .in1(N__11879),
            .in2(N__10973),
            .in3(N__12223),
            .lcout(),
            .ltout(\DUT.uart_inst0.g0_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_3_LC_12_15_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_3_LC_12_15_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_3_LC_12_15_3 .LUT_INIT=16'b0000001100000101;
    LogicCell40 \DUT.uart_inst0.tx_countdown_3_LC_12_15_3  (
            .in0(N__10958),
            .in1(N__10970),
            .in2(N__10961),
            .in3(N__12116),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13029),
            .ce(N__11975),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_2_3_LC_12_15_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_2_3_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_2_3_LC_12_15_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_2_3_LC_12_15_4  (
            .in0(N__11880),
            .in1(N__11724),
            .in2(_gnd_net_),
            .in3(N__11768),
            .lcout(\DUT.uart_inst0.g0_i_a6_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_4_LC_12_15_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_4_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_4_LC_12_15_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_0_4_LC_12_15_5  (
            .in0(N__11767),
            .in1(N__11881),
            .in2(N__11728),
            .in3(N__12169),
            .lcout(\DUT.uart_inst0.g0_i_o2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_2_5_LC_12_15_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_2_5_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_2_5_LC_12_15_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_2_5_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(N__11878),
            .in2(_gnd_net_),
            .in3(N__11766),
            .lcout(),
            .ltout(\DUT.uart_inst0.g0_i_o2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_5_LC_12_15_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_5_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_5_LC_12_15_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_0_5_LC_12_15_7  (
            .in0(N__11723),
            .in1(N__11919),
            .in2(N__10952),
            .in3(N__12168),
            .lcout(\DUT.uart_inst0.g0_i_o2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNI67HK1_5_LC_12_16_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNI67HK1_5_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNI67HK1_5_LC_12_16_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNI67HK1_5_LC_12_16_0  (
            .in0(N__11910),
            .in1(N__11868),
            .in2(N__11829),
            .in3(N__11717),
            .lcout(\DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0 ),
            .ltout(\DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNIJKPE2_1_LC_12_16_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNIJKPE2_1_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNIJKPE2_1_LC_12_16_1 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNIJKPE2_1_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__11764),
            .in2(N__11225),
            .in3(N__12154),
            .lcout(\DUT.uart_inst0.N_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_4_LC_12_16_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_4_LC_12_16_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_4_LC_12_16_2 .LUT_INIT=16'b0011000000010010;
    LogicCell40 \DUT.uart_inst0.tx_countdown_4_LC_12_16_2  (
            .in0(N__12225),
            .in1(N__11342),
            .in2(N__11920),
            .in3(N__11210),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13024),
            .ce(N__11977),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_5_LC_12_16_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_5_LC_12_16_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_5_LC_12_16_3 .LUT_INIT=16'b0000100100001100;
    LogicCell40 \DUT.uart_inst0.tx_countdown_5_LC_12_16_3  (
            .in0(N__11204),
            .in1(N__11821),
            .in2(N__11198),
            .in3(N__12226),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13024),
            .ce(N__11977),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_2_LC_12_16_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_2_LC_12_16_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_2_LC_12_16_4 .LUT_INIT=16'b1111110111110101;
    LogicCell40 \DUT.uart_inst0.tx_countdown_2_LC_12_16_4  (
            .in0(N__11693),
            .in1(N__11183),
            .in2(N__11171),
            .in3(N__11786),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13024),
            .ce(N__11977),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNIUUGK1_2_LC_12_16_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNIUUGK1_2_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNIUUGK1_2_LC_12_16_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNIUUGK1_2_LC_12_16_5  (
            .in0(N__11718),
            .in1(N__11763),
            .in2(N__11883),
            .in3(N__12153),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_state_ns_i_i_o2_a0_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNIJKPE2_5_LC_12_16_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNIJKPE2_5_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNIJKPE2_5_LC_12_16_6 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNIJKPE2_5_LC_12_16_6  (
            .in0(N__11911),
            .in1(_gnd_net_),
            .in2(N__11153),
            .in3(N__11822),
            .lcout(\DUT.uart_inst0.N_71_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_1_LC_12_16_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_1_LC_12_16_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_1_LC_12_16_7 .LUT_INIT=16'b0000100100001010;
    LogicCell40 \DUT.uart_inst0.tx_countdown_1_LC_12_16_7  (
            .in0(N__11773),
            .in1(N__12155),
            .in2(N__11138),
            .in3(N__12224),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13024),
            .ce(N__11977),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_0_LC_12_17_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_0_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_0_LC_12_17_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_0_0_LC_12_17_0  (
            .in0(N__11608),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11684),
            .lcout(),
            .ltout(\DUT.uart_inst0.g0_i_a3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_0_LC_12_17_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_0_LC_12_17_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_0_LC_12_17_1 .LUT_INIT=16'b0110011000000110;
    LogicCell40 \DUT.uart_inst0.tx_countdown_0_LC_12_17_1  (
            .in0(N__12217),
            .in1(N__12167),
            .in2(N__12077),
            .in3(N__11433),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13018),
            .ce(N__11981),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_5_2_LC_12_17_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_5_2_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_5_2_LC_12_17_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_5_2_LC_12_17_2  (
            .in0(N__11918),
            .in1(N__11884),
            .in2(N__11833),
            .in3(N__12156),
            .lcout(),
            .ltout(\DUT.uart_inst0.g0_11_a3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_2_2_LC_12_17_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_2_2_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_2_2_LC_12_17_3 .LUT_INIT=16'b1010000010110001;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_2_2_LC_12_17_3  (
            .in0(N__12216),
            .in1(N__11795),
            .in2(N__11789),
            .in3(N__12166),
            .lcout(\DUT.uart_inst0.N_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_2_LC_12_17_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_2_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_2_LC_12_17_4 .LUT_INIT=16'b0001111000001111;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_1_2_LC_12_17_4  (
            .in0(N__11772),
            .in1(N__12157),
            .in2(N__11729),
            .in3(N__12215),
            .lcout(\DUT.uart_inst0.N_6_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_4_LC_12_17_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_4_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_4_LC_12_17_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_1_4_LC_12_17_7  (
            .in0(N__11685),
            .in1(N__11607),
            .in2(_gnd_net_),
            .in3(N__11432),
            .lcout(\DUT.uart_inst0.N_11_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_8_LC_12_18_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_8_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_8_LC_12_18_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_8_LC_12_18_0  (
            .in0(N__11329),
            .in1(N__11317),
            .in2(N__11305),
            .in3(N__11287),
            .lcout(\DUT.uart_inst0.un1_tx_clk_divider_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_0_LC_12_18_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_0_LC_12_18_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_0_LC_12_18_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_0_LC_12_18_1  (
            .in0(N__11239),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12636),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13013),
            .ce(),
            .sr(N__11276));
    defparam \DUT.uart_inst0.tx_clk_divider_RNIBPK2_0_LC_12_18_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNIBPK2_0_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNIBPK2_0_LC_12_18_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNIBPK2_0_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(N__11251),
            .in2(_gnd_net_),
            .in3(N__11238),
            .lcout(\DUT.uart_inst0.un1_tx_clk_divider_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_RNI2V95_2_LC_12_18_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI2V95_2_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI2V95_2_LC_12_18_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNI2V95_2_LC_12_18_3  (
            .in0(N__12349),
            .in1(N__12337),
            .in2(N__12326),
            .in3(N__12310),
            .lcout(\DUT.uart_inst0.un1_tx_clk_divider_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_13_LC_12_18_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_13_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_13_LC_12_18_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_13_LC_12_18_4  (
            .in0(N__12298),
            .in1(N__12286),
            .in2(N__12275),
            .in3(N__12259),
            .lcout(),
            .ltout(\DUT.uart_inst0.un1_tx_clk_divider_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_RNITC2S1_0_LC_12_18_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNITC2S1_0_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNITC2S1_0_LC_12_18_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNITC2S1_0_LC_12_18_5  (
            .in0(N__12248),
            .in1(N__12242),
            .in2(N__12236),
            .in3(N__12233),
            .lcout(\DUT.uart_inst0.un1_tx_clk_divider_0 ),
            .ltout(\DUT.uart_inst0.un1_tx_clk_divider_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_3_3_LC_12_18_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_3_3_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_3_3_LC_12_18_6 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_3_3_LC_12_18_6  (
            .in0(N__12158),
            .in1(_gnd_net_),
            .in2(N__12119),
            .in3(_gnd_net_),
            .lcout(\DUT.uart_inst0.N_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_12_19_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_12_19_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_12_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_12_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13106),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13007),
            .ce(N__12527),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_12_19_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_12_19_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_12_19_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_12_19_1  (
            .in0(N__13276),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13007),
            .ce(N__12527),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_12_19_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_12_19_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_12_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_12_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12500),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13007),
            .ce(N__12527),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_12_19_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_12_19_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_12_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12446),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13007),
            .ce(N__12527),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_12_19_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_12_19_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_12_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_12_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12398),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13007),
            .ce(N__12527),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_12_19_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_12_19_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_12_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_12_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13148),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13007),
            .ce(N__12527),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_12_19_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_12_19_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_12_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_12_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13229),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13007),
            .ce(N__12527),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_12_19_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_12_19_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_12_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_12_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13322),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13007),
            .ce(N__12527),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_12_20_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_12_20_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_12_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_12_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13275),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13004),
            .ce(N__12879),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_12_20_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_12_20_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_12_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_12_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12498),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13004),
            .ce(N__12879),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_12_20_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_12_20_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_12_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_12_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12445),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13004),
            .ce(N__12879),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_12_20_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_12_20_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_12_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_12_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12397),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13004),
            .ce(N__12879),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_12_20_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_12_20_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_12_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_12_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13228),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13004),
            .ce(N__12879),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_12_20_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_12_20_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_12_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_12_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13321),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13004),
            .ce(N__12879),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_12_21_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_12_21_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_12_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_12_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13274),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13002),
            .ce(N__13188),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_12_21_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_12_21_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_12_21_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_12_21_1  (
            .in0(_gnd_net_),
            .in1(N__13216),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13002),
            .ce(N__13188),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_12_22_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_12_22_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_12_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_12_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13147),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13000),
            .ce(N__12884),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_13_20_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_13_20_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_13_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_13_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13105),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__13010),
            .ce(N__12883),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_14_21_2.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_14_21_2.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_14_21_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_14_21_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // top
