-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Mar 29 2020 11:31:56

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    ioFifoData : inout std_logic_vector(7 downto 0);
    P1A9 : out std_logic;
    P1A1 : in std_logic;
    P1A8 : out std_logic;
    oRx_n : out std_logic;
    P1A7 : out std_logic;
    P1A3 : out std_logic;
    iTxE_n : in std_logic;
    iRxF_n : in std_logic;
    iClk : in std_logic;
    P1A2 : out std_logic;
    BTN_N : in std_logic;
    BTN1 : in std_logic;
    oTx_n : out std_logic;
    P1A4 : out std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__13366\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13315\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13252\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13242\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13233\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13207\ : std_logic;
signal \N__13206\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13158\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13147\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13108\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13083\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13049\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13034\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13004\ : std_logic;
signal \N__13003\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12996\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12973\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12965\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12950\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12939\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12901\ : std_logic;
signal \N__12898\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12883\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12877\ : std_logic;
signal \N__12874\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12848\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12839\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12830\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12824\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12820\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12814\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12803\ : std_logic;
signal \N__12802\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12793\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12787\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12784\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12781\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12779\ : std_logic;
signal \N__12778\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12775\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12769\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12637\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12613\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12565\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12552\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12454\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12410\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12383\ : std_logic;
signal \N__12380\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12353\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12347\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12344\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12289\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12281\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12272\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12257\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12136\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12100\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11950\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11240\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10947\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10684\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10292\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9807\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9753\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9707\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9300\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9219\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9210\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7972\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7895\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7775\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7713\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7657\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7648\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7371\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7326\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7131\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6633\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6351\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \BTN_N_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_0\ : std_logic;
signal \bfn_12_4_0_\ : std_logic;
signal \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0\ : std_logic;
signal \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1\ : std_logic;
signal \un1_oRxFlag_0_i_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoCount_RNITA8H2Z0Z_1\ : std_logic;
signal \rFifoCount_RNIHH0D1_0_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0\ : std_logic;
signal \ioFifoData_in_6\ : std_logic;
signal \ioFifoData_in_0\ : std_logic;
signal \ioFifoData_in_4\ : std_logic;
signal \wRxFifoData_0\ : std_logic;
signal \DUT.rFifoDatarx_0\ : std_logic;
signal \wRxFifoData_4\ : std_logic;
signal \wRxFifoData_6\ : std_logic;
signal \DUT.rFifoDatarx_6\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDataro_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDataro_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_6\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_7\ : std_logic;
signal \DUT.fifo_rx_inst.rReadPtr_RNIDU4H2Z0Z_0_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_6\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6\ : std_logic;
signal \DUT.fifo_rx_inst.rReadPtr_RNIDU4H2Z0Z_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_4\ : std_logic;
signal \DUT.rFifoDatarx_0_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_5\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_5\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_6\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_4\ : std_logic;
signal \wPllLocked_i\ : std_logic;
signal \DUT.uart_inst0.N_275_cascade_\ : std_logic;
signal \DUT.uart_inst0.g0_0_5_cascade_\ : std_logic;
signal \DUT.uart_inst0.g0_6_cascade_\ : std_logic;
signal \DUT.uart_inst0.g0_1_0\ : std_logic;
signal \DUT.uart_inst0.g3_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.g0_0_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoCountZ0Z_1\ : std_logic;
signal \DUT.fifo_rx_inst.N_148\ : std_logic;
signal \ioFifoData_in_7\ : std_logic;
signal \ioFifoData_in_1\ : std_logic;
signal \ioFifoData_in_3\ : std_logic;
signal \ioFifoData_in_5\ : std_logic;
signal \ioFifoData_in_2\ : std_logic;
signal \wRxFifoData_1\ : std_logic;
signal \wRxFifoData_2\ : std_logic;
signal \wRxFifoData_3\ : std_logic;
signal \DUT.rFifoDatarx_0_5\ : std_logic;
signal \wRxFifoData_5\ : std_logic;
signal \DUT.rFifoDatarx_0_7\ : std_logic;
signal \wRxFifoData_7\ : std_logic;
signal \un1_oRxFlag_0_i_0\ : std_logic;
signal \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1\ : std_logic;
signal \DUT.rFifoDatarx_0_1\ : std_logic;
signal \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1\ : std_logic;
signal \DUT.wRcvd\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoCountZ0Z_2\ : std_logic;
signal \DUT.fifo_rx_inst.N_194_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2_cascade_\ : std_logic;
signal \DUT.rFifoDatarx_0_2\ : std_logic;
signal \DUT.rFifoDataror_0_0_cascade_\ : std_logic;
signal \DUT.rFifoDataror_1\ : std_logic;
signal \DUT.uart_inst0.N_257\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_\ : std_logic;
signal \DUT.rFifoDatarx_3\ : std_logic;
signal \DUT.fifo_rx_inst.rReadPtrZ0Z_0\ : std_logic;
signal \DUT.fifo_rx_inst.rReadPtrZ0Z_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_awe0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_5\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_5_i_a2_1_3\ : std_logic;
signal \DUT.uart_inst0.N_222_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_5_i_a2_11_0_5_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_5_i_a2_11_5\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_5_i_a2_11_5_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_221\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_0_0_c_RNOZ0\ : std_logic;
signal \bfn_14_3_0_\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_0Z0Z_0\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_0\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_1Z0Z_0\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_1\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_RNIP8N2BZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_2\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_2Z0Z_0\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_3\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_4\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_5_cascade_\ : std_logic;
signal \DUT.uart_inst0.g3_4\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_i_3\ : std_logic;
signal \DUT.uart_inst0.N_275\ : std_logic;
signal \DUT.uart_inst0.N_196_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_33_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_3_0_c_RNIP8IZ0Z482\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remaining_RNO_0Z0Z_1\ : std_logic;
signal \DUT.uart_inst0.g0_8_1\ : std_logic;
signal \P1A2_c_0_0\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_4\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rFifoState_0_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_6\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_awe3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDataro_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_awe2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDataro_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_awe1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_awe3_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.un1_i11_i\ : std_logic;
signal \DUT.fifo_tx_inst.un1_i11_i_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.N_194\ : std_logic;
signal \DUT.fifo_rx_inst.rWritePtrZ0Z_0\ : std_logic;
signal \DUT.fifo_rx_inst.rWritePtrZ0Z_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_5\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_awe1\ : std_logic;
signal \bfn_15_1_0_\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_0\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_1\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_3\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_2\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_4\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_3\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_5\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_4\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_6\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_6\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_5\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_7\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_6\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_7\ : std_logic;
signal \bfn_15_2_0_\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_8\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_9\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_10\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_11\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_12\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_14\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_13\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_15\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_15\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_14\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_15\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_16\ : std_logic;
signal \bfn_15_3_0_\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_16\ : std_logic;
signal \DUT.uart_inst0.recv_state_RNO_2Z0Z_4_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa_0_a2_0_a2_0_a3_1\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_8_i_0_o2_1_2_2_cascade_\ : std_logic;
signal \DUT.uart_inst0.recv_state_ns_0_i_0_0_o2_0_3\ : std_logic;
signal \DUT.uart_inst0.G_9_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.G_11_i_a4_0_4\ : std_logic;
signal \DUT.uart_inst0.N_4_i_1\ : std_logic;
signal \DUT.wRxByte_1\ : std_logic;
signal \DUT.wRxByte_0\ : std_logic;
signal \DUT.wRxByte_4\ : std_logic;
signal \DUT.wRxByte_5\ : std_logic;
signal \DUT.wRxByte_6\ : std_logic;
signal \DUT.wRxByte_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_awe3\ : std_logic;
signal \rTxByteZ0Z_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_0\ : std_logic;
signal \rTxByteZ0Z_1\ : std_logic;
signal \rTxByteZ0Z_3\ : std_logic;
signal \rTxByteZ0Z_6\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_4\ : std_logic;
signal \rTxByteZ0Z_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_\ : std_logic;
signal \rTxByteZ0Z_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_6\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_6\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoDataro_3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoDataro_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoDataro_1\ : std_logic;
signal \DUT.rFifoDataror_0_0_0\ : std_logic;
signal \DUT.rFifoDataror_1_0_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_6\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_6\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6\ : std_logic;
signal \DUT.fifo_tx_inst.rWritePtrZ0Z_0\ : std_logic;
signal \DUT.fifo_tx_inst.N_79_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rWritePtrZ0Z_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_awe2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoDataro_2\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rWrDelayZ0\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_3\ : std_logic;
signal \P1A4_c\ : std_logic;
signal \rTxBusReady\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_8\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_8\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_9\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_9\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_11\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_11\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_12\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_12\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_7\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_1\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ1Z_1\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_1\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_2\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.g0_0_3\ : std_logic;
signal \DUT.uart_inst0.g1\ : std_logic;
signal \DUT.uart_inst0.g0_0_0\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_17\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_17\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_10\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_10\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_13\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_13\ : std_logic;
signal \DUT.uart_inst0.N_199_0\ : std_logic;
signal \N_1239_i\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_5_i_a2_12_1_5\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_16\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_5_i_a2_12_4_5\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_14\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_5_i_a2_12_5\ : std_logic;
signal \DUT.uart_inst0.N_31_0\ : std_logic;
signal \DUT.uart_inst0.N_203\ : std_logic;
signal \DUT.uart_inst0.recv_state_ns_0_i_0_0_a3_0_0_3\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remainingZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remainingZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remainingZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remainingZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.N_215_4\ : std_logic;
signal \DUT.uart_inst0.N_215_4_cascade_\ : std_logic;
signal \DUT.uart_inst0.recv_state_srsts_1_2_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_193\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.g0_0\ : std_logic;
signal \DUT.wRxByte_3\ : std_logic;
signal \DUT.wRxByte_2\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_3\ : std_logic;
signal \DUT.rFifoDatarx_0_0\ : std_logic;
signal \DUT.uart_inst0.tx_out_6_iv_0_1\ : std_logic;
signal \DUT.rFifoDatarx_1\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_1\ : std_logic;
signal \DUT.rFifoDatarx_2\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_2\ : std_logic;
signal \DUT.rFifoDatarx_0_3\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_7\ : std_logic;
signal \DUT.uart_inst0.tx_out_6_iv_0_a3_0_1\ : std_logic;
signal \DUT.uart_inst0.N_101\ : std_logic;
signal \DUT.rFifoDatarx_5\ : std_logic;
signal \DUT.rFifoDatarx_0_6\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_6\ : std_logic;
signal \DUT.rFifoDatarx_4\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_4\ : std_logic;
signal \DUT.rFifoDatarx_7\ : std_logic;
signal \DUT.uart_inst0.N_145\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_7\ : std_logic;
signal \DUT.uart_inst0.N_22_i\ : std_logic;
signal \DUT.fifo_tx_inst.N_83_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_0\ : std_logic;
signal \P1A7_c\ : std_logic;
signal \DUT.uart_inst0.N_98\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rFifoStatec_0\ : std_logic;
signal \DUT.fifo_tx_inst.N_79\ : std_logic;
signal \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoCountZ0Z_0\ : std_logic;
signal \bfn_16_11_0_\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoCount_RNISSQ21Z0Z_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoCountZ0Z_1\ : std_logic;
signal \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0\ : std_logic;
signal \DUT.fifo_tx_inst.N_83\ : std_logic;
signal \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoCountZ0Z_2\ : std_logic;
signal \P1A1_c\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.g0_1\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_4\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_5\ : std_logic;
signal \DUT.uart_inst0.recv_state_RNO_2Z0Z_1\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_0\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_2\ : std_logic;
signal \DUT.uart_inst0.G_10_i_a4_0_4_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_3\ : std_logic;
signal \DUT.uart_inst0.N_4_i_0_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_149\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_1\ : std_logic;
signal \rRxReadZ0\ : std_logic;
signal \DUT.fifo_rx_inst.N_206\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoCountZ0Z_0\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1\ : std_logic;
signal \P1A2_c\ : std_logic;
signal \rFifoCount_RNIHH0D1_0\ : std_logic;
signal \rTxWriteZ0\ : std_logic;
signal \P1A3_c\ : std_logic;
signal \rTxByteZ0Z_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_2\ : std_logic;
signal \rTxByteZ0Z_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_awe0\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remainingZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remainingZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remainingZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.N_142_cascade_\ : std_logic;
signal \wPllLocked\ : std_logic;
signal \DUT.uart_inst0.N_84_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_22\ : std_logic;
signal \DUT.uart_inst0.N_22_cascade_\ : std_logic;
signal \DUT.uart_inst0.un1_tx_bits_remaining_c3\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remainingZ0Z_3\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2\ : std_logic;
signal \fifo_inst.ftdi_output_inst.N_78_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_142\ : std_logic;
signal \DUT.uart_inst0.N_144\ : std_logic;
signal \DUT.uart_inst0.N_74_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_143\ : std_logic;
signal \DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_75\ : std_logic;
signal \DUT.uart_inst0.N_75_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_7s2_0_0\ : std_logic;
signal \DUT.uart_inst0.tx_state_ns_i_i_o2_a0_3_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_69_i\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_30_3_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_84\ : std_logic;
signal \DUT.uart_inst0.N_30_1\ : std_logic;
signal \N_1242_i\ : std_logic;
signal \N_1240_i\ : std_logic;
signal \rTxBusReady_rep1_i_ess\ : std_logic;
signal \rTxBusReady_rep3_i_ess\ : std_logic;
signal \rTxBusReady_rep0_i_ess\ : std_logic;
signal \iTxE_n_c\ : std_logic;
signal \fifo_inst.ftdi_output_inst.N_68_0\ : std_logic;
signal \wPllLocked_i_g\ : std_logic;
signal \fifo_inst.ftdi_output_inst.un1_oTx_n_1_sqmuxa_0_i_cascade_\ : std_logic;
signal \fifo_inst.ftdi_output_inst.un1_oTx_n_1_sqmuxa_0_i_0\ : std_logic;
signal \iRxF_n_c\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0\ : std_logic;
signal \fifo_inst.ftdi_output_inst.N_80\ : std_logic;
signal \DUT.uart_inst0.N_77_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_state_RNI8CH01Z0Z_1\ : std_logic;
signal \DUT.uart_inst0.tx_state_RNI8CH01Z0Z_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_59_i\ : std_logic;
signal \DUT.N_93\ : std_logic;
signal \DUT.tx_state_1\ : std_logic;
signal \DUT.rTransmitZ0\ : std_logic;
signal \DUT.fifo_tx_inst.rReadPtrZ0Z_1\ : std_logic;
signal \DUT.fifo_tx_inst.un1_i11_2_i\ : std_logic;
signal \DUT.fifo_tx_inst.rReadPtr11\ : std_logic;
signal \DUT.fifo_tx_inst.un1_i11_2_i_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rReadPtrZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.N_74\ : std_logic;
signal \DUT.tx_state_0\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_7_1_2\ : std_logic;
signal \DUT.uart_inst0.N_91\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_0_c4_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_7_ns_1_4\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_7_ns_1_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_0_c4\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_7_ns_1_5\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_7_m1_0_o2_1_2_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.N_68\ : std_logic;
signal \DUT.uart_inst0.N_146\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_7_sm0_0\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_7_ns_1_3\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_3\ : std_logic;
signal \rTxBusReady_rep2_i_ess\ : std_logic;
signal \N_1241_i\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_9\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_6_cascade_\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_0_cascade_\ : std_logic;
signal \wPllLocked_g\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_8\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_7\ : std_logic;
signal \DUT.uart_inst0.N_77\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_0\ : std_logic;
signal \DUT.uart_inst0.N_147\ : std_logic;
signal \bfn_21_9_0_\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_0\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_1\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_2\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_3\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_4\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_6\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_5\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_7\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_6\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_7\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_8\ : std_logic;
signal \bfn_21_10_0_\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_9\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_8\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_10\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_9\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_11\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_10\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_12\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_11\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_12\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_13\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_0\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_48mhz : std_logic;
signal \DUT.uart_inst0.N_20\ : std_logic;

signal \iClk_wire\ : std_logic;
signal \P1A8_wire\ : std_logic;
signal \P1A4_wire\ : std_logic;
signal \oRx_n_wire\ : std_logic;
signal \P1A2_wire\ : std_logic;
signal \iRxF_n_wire\ : std_logic;
signal \P1A3_wire\ : std_logic;
signal \P1A7_wire\ : std_logic;
signal \BTN_N_wire\ : std_logic;
signal \oTx_n_wire\ : std_logic;
signal \iTxE_n_wire\ : std_logic;
signal \P1A1_wire\ : std_logic;
signal \P1A9_wire\ : std_logic;
signal \top_pll_inst.top_pll_inst_pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \iClk_wire\ <= iClk;
    P1A8 <= \P1A8_wire\;
    P1A4 <= \P1A4_wire\;
    oRx_n <= \oRx_n_wire\;
    P1A2 <= \P1A2_wire\;
    \iRxF_n_wire\ <= iRxF_n;
    P1A3 <= \P1A3_wire\;
    P1A7 <= \P1A7_wire\;
    \BTN_N_wire\ <= BTN_N;
    oTx_n <= \oTx_n_wire\;
    \iTxE_n_wire\ <= iTxE_n;
    \P1A1_wire\ <= P1A1;
    P1A9 <= \P1A9_wire\;
    \top_pll_inst.top_pll_inst_pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \top_pll_inst.top_pll_inst_pll\ : PLL40
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "0111111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            PLLOUTGLOBAL => clk_48mhz,
            SDI => \GNDG0\,
            BYPASS => \GNDG0\,
            RESETB => \N__5089\,
            PLLOUTCORE => OPEN,
            LOCK => \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO\,
            SDO => OPEN,
            SCLK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            EXTFEEDBACK => \GNDG0\,
            DYNAMICDELAY => \top_pll_inst.top_pll_inst_pll_DYNAMICDELAY_wire\,
            PLLIN => \N__13366\
        );

    \top_pll_inst.top_pll_inst_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \VCCG0\,
            DIN => '0',
            DOUT => \N__13366\,
            PACKAGEPIN => \iClk_wire\
        );

    \P1A8_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13352\,
            DIN => \N__13351\,
            DOUT => \N__13350\,
            PACKAGEPIN => \P1A8_wire\
        );

    \P1A8_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13352\,
            PADOUT => \N__13351\,
            PADIN => \N__13350\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13343\,
            DIN => \N__13342\,
            DOUT => \N__13341\,
            PACKAGEPIN => ioFifoData(6)
        );

    \ioFifoData_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13343\,
            PADOUT => \N__13342\,
            PADIN => \N__13341\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7830\,
            DIN0 => \ioFifoData_in_6\,
            DOUT0 => \N__12960\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13334\,
            DIN => \N__13333\,
            DOUT => \N__13332\,
            PACKAGEPIN => ioFifoData(3)
        );

    \ioFifoData_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13334\,
            PADOUT => \N__13333\,
            PADIN => \N__13332\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10819\,
            DIN0 => \ioFifoData_in_3\,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A4_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13325\,
            DIN => \N__13324\,
            DOUT => \N__13323\,
            PACKAGEPIN => \P1A4_wire\
        );

    \P1A4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13325\,
            PADOUT => \N__13324\,
            PADIN => \N__13323\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7873\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \oRx_n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13316\,
            DIN => \N__13315\,
            DOUT => \N__13314\,
            PACKAGEPIN => \oRx_n_wire\
        );

    \oRx_n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13316\,
            PADOUT => \N__13315\,
            PADIN => \N__13314\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10182\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13307\,
            DIN => \N__13306\,
            DOUT => \N__13305\,
            PACKAGEPIN => \P1A2_wire\
        );

    \P1A2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13307\,
            PADOUT => \N__13306\,
            PADIN => \N__13305\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10351\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13298\,
            DIN => \N__13297\,
            DOUT => \N__13296\,
            PACKAGEPIN => ioFifoData(0)
        );

    \ioFifoData_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13298\,
            PADOUT => \N__13297\,
            PADIN => \N__13296\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__8296\,
            DIN0 => \ioFifoData_in_0\,
            DOUT0 => \N__13041\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \iRxF_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13289\,
            DIN => \N__13288\,
            DOUT => \N__13287\,
            PACKAGEPIN => \iRxF_n_wire\
        );

    \iRxF_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13289\,
            PADOUT => \N__13288\,
            PADIN => \N__13287\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \iRxF_n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13280\,
            DIN => \N__13279\,
            DOUT => \N__13278\,
            PACKAGEPIN => \P1A3_wire\
        );

    \P1A3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13280\,
            PADOUT => \N__13279\,
            PADIN => \N__13278\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10195\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A7_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13271\,
            DIN => \N__13270\,
            DOUT => \N__13269\,
            PACKAGEPIN => \P1A7_wire\
        );

    \P1A7_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13271\,
            PADOUT => \N__13270\,
            PADIN => \N__13269\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9060\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13262\,
            DIN => \N__13261\,
            DOUT => \N__13260\,
            PACKAGEPIN => ioFifoData(7)
        );

    \ioFifoData_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13262\,
            PADOUT => \N__13261\,
            PADIN => \N__13260\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7831\,
            DIN0 => \ioFifoData_in_7\,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BTN_N_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13253\,
            DIN => \N__13252\,
            DOUT => \N__13251\,
            PACKAGEPIN => \BTN_N_wire\
        );

    \BTN_N_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13253\,
            PADOUT => \N__13252\,
            PADIN => \N__13251\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \BTN_N_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13244\,
            DIN => \N__13243\,
            DOUT => \N__13242\,
            PACKAGEPIN => ioFifoData(4)
        );

    \ioFifoData_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13244\,
            PADOUT => \N__13243\,
            PADIN => \N__13242\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7829\,
            DIN0 => \ioFifoData_in_4\,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13235\,
            DIN => \N__13234\,
            DOUT => \N__13233\,
            PACKAGEPIN => ioFifoData(1)
        );

    \ioFifoData_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13235\,
            PADOUT => \N__13234\,
            PADIN => \N__13233\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__10807\,
            DIN0 => \ioFifoData_in_1\,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13226\,
            DIN => \N__13225\,
            DOUT => \N__13224\,
            PACKAGEPIN => ioFifoData(5)
        );

    \ioFifoData_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13226\,
            PADOUT => \N__13225\,
            PADIN => \N__13224\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__7819\,
            DIN0 => \ioFifoData_in_5\,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \oTx_n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13217\,
            DIN => \N__13216\,
            DOUT => \N__13215\,
            PACKAGEPIN => \oTx_n_wire\
        );

    \oTx_n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13217\,
            PADOUT => \N__13216\,
            PADIN => \N__13215\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7869\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \iTxE_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13208\,
            DIN => \N__13207\,
            DOUT => \N__13206\,
            PACKAGEPIN => \iTxE_n_wire\
        );

    \iTxE_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13208\,
            PADOUT => \N__13207\,
            PADIN => \N__13206\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \iTxE_n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13199\,
            DIN => \N__13198\,
            DOUT => \N__13197\,
            PACKAGEPIN => \P1A1_wire\
        );

    \P1A1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13199\,
            PADOUT => \N__13198\,
            PADIN => \N__13197\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \P1A1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13190\,
            DIN => \N__13189\,
            DOUT => \N__13188\,
            PACKAGEPIN => ioFifoData(2)
        );

    \ioFifoData_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13190\,
            PADOUT => \N__13189\,
            PADIN => \N__13188\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__12466\,
            DIN0 => \ioFifoData_in_2\,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A9_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13181\,
            DIN => \N__13180\,
            DOUT => \N__13179\,
            PACKAGEPIN => \P1A9_wire\
        );

    \P1A9_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13181\,
            PADOUT => \N__13180\,
            PADIN => \N__13179\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__3123\ : CascadeMux
    port map (
            O => \N__13162\,
            I => \N__13159\
        );

    \I__3122\ : InMux
    port map (
            O => \N__13159\,
            I => \N__13155\
        );

    \I__3121\ : InMux
    port map (
            O => \N__13158\,
            I => \N__13152\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__13155\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_9\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__13152\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_9\
        );

    \I__3118\ : InMux
    port map (
            O => \N__13147\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_8\
        );

    \I__3117\ : InMux
    port map (
            O => \N__13144\,
            I => \N__13140\
        );

    \I__3116\ : InMux
    port map (
            O => \N__13143\,
            I => \N__13137\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__13140\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_10\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__13137\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_10\
        );

    \I__3113\ : InMux
    port map (
            O => \N__13132\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_9\
        );

    \I__3112\ : CascadeMux
    port map (
            O => \N__13129\,
            I => \N__13125\
        );

    \I__3111\ : CascadeMux
    port map (
            O => \N__13128\,
            I => \N__13122\
        );

    \I__3110\ : InMux
    port map (
            O => \N__13125\,
            I => \N__13119\
        );

    \I__3109\ : InMux
    port map (
            O => \N__13122\,
            I => \N__13116\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__13119\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_11\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__13116\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_11\
        );

    \I__3106\ : InMux
    port map (
            O => \N__13111\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_10\
        );

    \I__3105\ : InMux
    port map (
            O => \N__13108\,
            I => \N__13104\
        );

    \I__3104\ : InMux
    port map (
            O => \N__13107\,
            I => \N__13101\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__13104\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_12\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__13101\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_12\
        );

    \I__3101\ : InMux
    port map (
            O => \N__13096\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_11\
        );

    \I__3100\ : InMux
    port map (
            O => \N__13093\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_12\
        );

    \I__3099\ : InMux
    port map (
            O => \N__13090\,
            I => \N__13086\
        );

    \I__3098\ : InMux
    port map (
            O => \N__13089\,
            I => \N__13083\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__13086\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_13\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__13083\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_13\
        );

    \I__3095\ : CascadeMux
    port map (
            O => \N__13078\,
            I => \N__13068\
        );

    \I__3094\ : CascadeMux
    port map (
            O => \N__13077\,
            I => \N__13065\
        );

    \I__3093\ : CascadeMux
    port map (
            O => \N__13076\,
            I => \N__13062\
        );

    \I__3092\ : CascadeMux
    port map (
            O => \N__13075\,
            I => \N__13059\
        );

    \I__3091\ : CascadeMux
    port map (
            O => \N__13074\,
            I => \N__13056\
        );

    \I__3090\ : CascadeMux
    port map (
            O => \N__13073\,
            I => \N__13052\
        );

    \I__3089\ : CascadeMux
    port map (
            O => \N__13072\,
            I => \N__13049\
        );

    \I__3088\ : CascadeMux
    port map (
            O => \N__13071\,
            I => \N__13046\
        );

    \I__3087\ : InMux
    port map (
            O => \N__13068\,
            I => \N__13034\
        );

    \I__3086\ : InMux
    port map (
            O => \N__13065\,
            I => \N__13034\
        );

    \I__3085\ : InMux
    port map (
            O => \N__13062\,
            I => \N__13034\
        );

    \I__3084\ : InMux
    port map (
            O => \N__13059\,
            I => \N__13023\
        );

    \I__3083\ : InMux
    port map (
            O => \N__13056\,
            I => \N__13023\
        );

    \I__3082\ : InMux
    port map (
            O => \N__13055\,
            I => \N__13023\
        );

    \I__3081\ : InMux
    port map (
            O => \N__13052\,
            I => \N__13023\
        );

    \I__3080\ : InMux
    port map (
            O => \N__13049\,
            I => \N__13023\
        );

    \I__3079\ : InMux
    port map (
            O => \N__13046\,
            I => \N__13020\
        );

    \I__3078\ : CascadeMux
    port map (
            O => \N__13045\,
            I => \N__13017\
        );

    \I__3077\ : CascadeMux
    port map (
            O => \N__13044\,
            I => \N__13013\
        );

    \I__3076\ : CascadeMux
    port map (
            O => \N__13043\,
            I => \N__13009\
        );

    \I__3075\ : CascadeMux
    port map (
            O => \N__13042\,
            I => \N__13005\
        );

    \I__3074\ : IoInMux
    port map (
            O => \N__13041\,
            I => \N__12999\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__13034\,
            I => \N__12993\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__13023\,
            I => \N__12988\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__13020\,
            I => \N__12988\
        );

    \I__3070\ : InMux
    port map (
            O => \N__13017\,
            I => \N__12973\
        );

    \I__3069\ : InMux
    port map (
            O => \N__13016\,
            I => \N__12973\
        );

    \I__3068\ : InMux
    port map (
            O => \N__13013\,
            I => \N__12973\
        );

    \I__3067\ : InMux
    port map (
            O => \N__13012\,
            I => \N__12973\
        );

    \I__3066\ : InMux
    port map (
            O => \N__13009\,
            I => \N__12973\
        );

    \I__3065\ : InMux
    port map (
            O => \N__13008\,
            I => \N__12973\
        );

    \I__3064\ : InMux
    port map (
            O => \N__13005\,
            I => \N__12973\
        );

    \I__3063\ : CascadeMux
    port map (
            O => \N__13004\,
            I => \N__12969\
        );

    \I__3062\ : CascadeMux
    port map (
            O => \N__13003\,
            I => \N__12966\
        );

    \I__3061\ : CascadeMux
    port map (
            O => \N__13002\,
            I => \N__12962\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__12999\,
            I => \N__12957\
        );

    \I__3059\ : CascadeMux
    port map (
            O => \N__12998\,
            I => \N__12954\
        );

    \I__3058\ : CascadeMux
    port map (
            O => \N__12997\,
            I => \N__12950\
        );

    \I__3057\ : CascadeMux
    port map (
            O => \N__12996\,
            I => \N__12946\
        );

    \I__3056\ : Span4Mux_v
    port map (
            O => \N__12993\,
            I => \N__12939\
        );

    \I__3055\ : Span4Mux_v
    port map (
            O => \N__12988\,
            I => \N__12939\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__12973\,
            I => \N__12936\
        );

    \I__3053\ : InMux
    port map (
            O => \N__12972\,
            I => \N__12923\
        );

    \I__3052\ : InMux
    port map (
            O => \N__12969\,
            I => \N__12923\
        );

    \I__3051\ : InMux
    port map (
            O => \N__12966\,
            I => \N__12923\
        );

    \I__3050\ : InMux
    port map (
            O => \N__12965\,
            I => \N__12923\
        );

    \I__3049\ : InMux
    port map (
            O => \N__12962\,
            I => \N__12923\
        );

    \I__3048\ : InMux
    port map (
            O => \N__12961\,
            I => \N__12923\
        );

    \I__3047\ : IoInMux
    port map (
            O => \N__12960\,
            I => \N__12920\
        );

    \I__3046\ : Span4Mux_s0_v
    port map (
            O => \N__12957\,
            I => \N__12917\
        );

    \I__3045\ : InMux
    port map (
            O => \N__12954\,
            I => \N__12912\
        );

    \I__3044\ : InMux
    port map (
            O => \N__12953\,
            I => \N__12912\
        );

    \I__3043\ : InMux
    port map (
            O => \N__12950\,
            I => \N__12901\
        );

    \I__3042\ : InMux
    port map (
            O => \N__12949\,
            I => \N__12901\
        );

    \I__3041\ : InMux
    port map (
            O => \N__12946\,
            I => \N__12901\
        );

    \I__3040\ : InMux
    port map (
            O => \N__12945\,
            I => \N__12901\
        );

    \I__3039\ : InMux
    port map (
            O => \N__12944\,
            I => \N__12901\
        );

    \I__3038\ : Span4Mux_v
    port map (
            O => \N__12939\,
            I => \N__12898\
        );

    \I__3037\ : Span4Mux_h
    port map (
            O => \N__12936\,
            I => \N__12893\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__12923\,
            I => \N__12893\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__12920\,
            I => \N__12890\
        );

    \I__3034\ : Sp12to4
    port map (
            O => \N__12917\,
            I => \N__12883\
        );

    \I__3033\ : LocalMux
    port map (
            O => \N__12912\,
            I => \N__12883\
        );

    \I__3032\ : LocalMux
    port map (
            O => \N__12901\,
            I => \N__12883\
        );

    \I__3031\ : Span4Mux_v
    port map (
            O => \N__12898\,
            I => \N__12880\
        );

    \I__3030\ : Span4Mux_v
    port map (
            O => \N__12893\,
            I => \N__12877\
        );

    \I__3029\ : IoSpan4Mux
    port map (
            O => \N__12890\,
            I => \N__12874\
        );

    \I__3028\ : Span12Mux_s11_h
    port map (
            O => \N__12883\,
            I => \N__12871\
        );

    \I__3027\ : Sp12to4
    port map (
            O => \N__12880\,
            I => \N__12866\
        );

    \I__3026\ : Sp12to4
    port map (
            O => \N__12877\,
            I => \N__12866\
        );

    \I__3025\ : Span4Mux_s3_v
    port map (
            O => \N__12874\,
            I => \N__12863\
        );

    \I__3024\ : Span12Mux_v
    port map (
            O => \N__12871\,
            I => \N__12858\
        );

    \I__3023\ : Span12Mux_s11_h
    port map (
            O => \N__12866\,
            I => \N__12858\
        );

    \I__3022\ : Span4Mux_v
    port map (
            O => \N__12863\,
            I => \N__12855\
        );

    \I__3021\ : Odrv12
    port map (
            O => \N__12858\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3020\ : Odrv4
    port map (
            O => \N__12855\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3019\ : InMux
    port map (
            O => \N__12850\,
            I => \N__12845\
        );

    \I__3018\ : InMux
    port map (
            O => \N__12849\,
            I => \N__12842\
        );

    \I__3017\ : InMux
    port map (
            O => \N__12848\,
            I => \N__12839\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__12845\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_0\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__12842\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_0\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__12839\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_0\
        );

    \I__3013\ : ClkMux
    port map (
            O => \N__12832\,
            I => \N__12640\
        );

    \I__3012\ : ClkMux
    port map (
            O => \N__12831\,
            I => \N__12640\
        );

    \I__3011\ : ClkMux
    port map (
            O => \N__12830\,
            I => \N__12640\
        );

    \I__3010\ : ClkMux
    port map (
            O => \N__12829\,
            I => \N__12640\
        );

    \I__3009\ : ClkMux
    port map (
            O => \N__12828\,
            I => \N__12640\
        );

    \I__3008\ : ClkMux
    port map (
            O => \N__12827\,
            I => \N__12640\
        );

    \I__3007\ : ClkMux
    port map (
            O => \N__12826\,
            I => \N__12640\
        );

    \I__3006\ : ClkMux
    port map (
            O => \N__12825\,
            I => \N__12640\
        );

    \I__3005\ : ClkMux
    port map (
            O => \N__12824\,
            I => \N__12640\
        );

    \I__3004\ : ClkMux
    port map (
            O => \N__12823\,
            I => \N__12640\
        );

    \I__3003\ : ClkMux
    port map (
            O => \N__12822\,
            I => \N__12640\
        );

    \I__3002\ : ClkMux
    port map (
            O => \N__12821\,
            I => \N__12640\
        );

    \I__3001\ : ClkMux
    port map (
            O => \N__12820\,
            I => \N__12640\
        );

    \I__3000\ : ClkMux
    port map (
            O => \N__12819\,
            I => \N__12640\
        );

    \I__2999\ : ClkMux
    port map (
            O => \N__12818\,
            I => \N__12640\
        );

    \I__2998\ : ClkMux
    port map (
            O => \N__12817\,
            I => \N__12640\
        );

    \I__2997\ : ClkMux
    port map (
            O => \N__12816\,
            I => \N__12640\
        );

    \I__2996\ : ClkMux
    port map (
            O => \N__12815\,
            I => \N__12640\
        );

    \I__2995\ : ClkMux
    port map (
            O => \N__12814\,
            I => \N__12640\
        );

    \I__2994\ : ClkMux
    port map (
            O => \N__12813\,
            I => \N__12640\
        );

    \I__2993\ : ClkMux
    port map (
            O => \N__12812\,
            I => \N__12640\
        );

    \I__2992\ : ClkMux
    port map (
            O => \N__12811\,
            I => \N__12640\
        );

    \I__2991\ : ClkMux
    port map (
            O => \N__12810\,
            I => \N__12640\
        );

    \I__2990\ : ClkMux
    port map (
            O => \N__12809\,
            I => \N__12640\
        );

    \I__2989\ : ClkMux
    port map (
            O => \N__12808\,
            I => \N__12640\
        );

    \I__2988\ : ClkMux
    port map (
            O => \N__12807\,
            I => \N__12640\
        );

    \I__2987\ : ClkMux
    port map (
            O => \N__12806\,
            I => \N__12640\
        );

    \I__2986\ : ClkMux
    port map (
            O => \N__12805\,
            I => \N__12640\
        );

    \I__2985\ : ClkMux
    port map (
            O => \N__12804\,
            I => \N__12640\
        );

    \I__2984\ : ClkMux
    port map (
            O => \N__12803\,
            I => \N__12640\
        );

    \I__2983\ : ClkMux
    port map (
            O => \N__12802\,
            I => \N__12640\
        );

    \I__2982\ : ClkMux
    port map (
            O => \N__12801\,
            I => \N__12640\
        );

    \I__2981\ : ClkMux
    port map (
            O => \N__12800\,
            I => \N__12640\
        );

    \I__2980\ : ClkMux
    port map (
            O => \N__12799\,
            I => \N__12640\
        );

    \I__2979\ : ClkMux
    port map (
            O => \N__12798\,
            I => \N__12640\
        );

    \I__2978\ : ClkMux
    port map (
            O => \N__12797\,
            I => \N__12640\
        );

    \I__2977\ : ClkMux
    port map (
            O => \N__12796\,
            I => \N__12640\
        );

    \I__2976\ : ClkMux
    port map (
            O => \N__12795\,
            I => \N__12640\
        );

    \I__2975\ : ClkMux
    port map (
            O => \N__12794\,
            I => \N__12640\
        );

    \I__2974\ : ClkMux
    port map (
            O => \N__12793\,
            I => \N__12640\
        );

    \I__2973\ : ClkMux
    port map (
            O => \N__12792\,
            I => \N__12640\
        );

    \I__2972\ : ClkMux
    port map (
            O => \N__12791\,
            I => \N__12640\
        );

    \I__2971\ : ClkMux
    port map (
            O => \N__12790\,
            I => \N__12640\
        );

    \I__2970\ : ClkMux
    port map (
            O => \N__12789\,
            I => \N__12640\
        );

    \I__2969\ : ClkMux
    port map (
            O => \N__12788\,
            I => \N__12640\
        );

    \I__2968\ : ClkMux
    port map (
            O => \N__12787\,
            I => \N__12640\
        );

    \I__2967\ : ClkMux
    port map (
            O => \N__12786\,
            I => \N__12640\
        );

    \I__2966\ : ClkMux
    port map (
            O => \N__12785\,
            I => \N__12640\
        );

    \I__2965\ : ClkMux
    port map (
            O => \N__12784\,
            I => \N__12640\
        );

    \I__2964\ : ClkMux
    port map (
            O => \N__12783\,
            I => \N__12640\
        );

    \I__2963\ : ClkMux
    port map (
            O => \N__12782\,
            I => \N__12640\
        );

    \I__2962\ : ClkMux
    port map (
            O => \N__12781\,
            I => \N__12640\
        );

    \I__2961\ : ClkMux
    port map (
            O => \N__12780\,
            I => \N__12640\
        );

    \I__2960\ : ClkMux
    port map (
            O => \N__12779\,
            I => \N__12640\
        );

    \I__2959\ : ClkMux
    port map (
            O => \N__12778\,
            I => \N__12640\
        );

    \I__2958\ : ClkMux
    port map (
            O => \N__12777\,
            I => \N__12640\
        );

    \I__2957\ : ClkMux
    port map (
            O => \N__12776\,
            I => \N__12640\
        );

    \I__2956\ : ClkMux
    port map (
            O => \N__12775\,
            I => \N__12640\
        );

    \I__2955\ : ClkMux
    port map (
            O => \N__12774\,
            I => \N__12640\
        );

    \I__2954\ : ClkMux
    port map (
            O => \N__12773\,
            I => \N__12640\
        );

    \I__2953\ : ClkMux
    port map (
            O => \N__12772\,
            I => \N__12640\
        );

    \I__2952\ : ClkMux
    port map (
            O => \N__12771\,
            I => \N__12640\
        );

    \I__2951\ : ClkMux
    port map (
            O => \N__12770\,
            I => \N__12640\
        );

    \I__2950\ : ClkMux
    port map (
            O => \N__12769\,
            I => \N__12640\
        );

    \I__2949\ : GlobalMux
    port map (
            O => \N__12640\,
            I => clk_48mhz
        );

    \I__2948\ : SRMux
    port map (
            O => \N__12637\,
            I => \N__12633\
        );

    \I__2947\ : SRMux
    port map (
            O => \N__12636\,
            I => \N__12630\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__12633\,
            I => \N__12627\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__12630\,
            I => \N__12624\
        );

    \I__2944\ : Span4Mux_v
    port map (
            O => \N__12627\,
            I => \N__12621\
        );

    \I__2943\ : Span4Mux_h
    port map (
            O => \N__12624\,
            I => \N__12618\
        );

    \I__2942\ : Odrv4
    port map (
            O => \N__12621\,
            I => \DUT.uart_inst0.N_20\
        );

    \I__2941\ : Odrv4
    port map (
            O => \N__12618\,
            I => \DUT.uart_inst0.N_20\
        );

    \I__2940\ : InMux
    port map (
            O => \N__12613\,
            I => \N__12609\
        );

    \I__2939\ : InMux
    port map (
            O => \N__12612\,
            I => \N__12606\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__12609\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_1\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__12606\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_1\
        );

    \I__2936\ : InMux
    port map (
            O => \N__12601\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_0\
        );

    \I__2935\ : CascadeMux
    port map (
            O => \N__12598\,
            I => \N__12595\
        );

    \I__2934\ : InMux
    port map (
            O => \N__12595\,
            I => \N__12591\
        );

    \I__2933\ : InMux
    port map (
            O => \N__12594\,
            I => \N__12588\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__12591\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_2\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__12588\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_2\
        );

    \I__2930\ : InMux
    port map (
            O => \N__12583\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_1\
        );

    \I__2929\ : CascadeMux
    port map (
            O => \N__12580\,
            I => \N__12576\
        );

    \I__2928\ : InMux
    port map (
            O => \N__12579\,
            I => \N__12573\
        );

    \I__2927\ : InMux
    port map (
            O => \N__12576\,
            I => \N__12570\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__12573\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_3\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__12570\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_3\
        );

    \I__2924\ : InMux
    port map (
            O => \N__12565\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_2\
        );

    \I__2923\ : CascadeMux
    port map (
            O => \N__12562\,
            I => \N__12559\
        );

    \I__2922\ : InMux
    port map (
            O => \N__12559\,
            I => \N__12555\
        );

    \I__2921\ : InMux
    port map (
            O => \N__12558\,
            I => \N__12552\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__12555\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_4\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__12552\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_4\
        );

    \I__2918\ : InMux
    port map (
            O => \N__12547\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_3\
        );

    \I__2917\ : InMux
    port map (
            O => \N__12544\,
            I => \N__12540\
        );

    \I__2916\ : InMux
    port map (
            O => \N__12543\,
            I => \N__12537\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__12540\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_5\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__12537\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_5\
        );

    \I__2913\ : InMux
    port map (
            O => \N__12532\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_4\
        );

    \I__2912\ : CascadeMux
    port map (
            O => \N__12529\,
            I => \N__12526\
        );

    \I__2911\ : InMux
    port map (
            O => \N__12526\,
            I => \N__12522\
        );

    \I__2910\ : InMux
    port map (
            O => \N__12525\,
            I => \N__12519\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__12522\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_6\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__12519\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_6\
        );

    \I__2907\ : InMux
    port map (
            O => \N__12514\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_5\
        );

    \I__2906\ : CascadeMux
    port map (
            O => \N__12511\,
            I => \N__12507\
        );

    \I__2905\ : InMux
    port map (
            O => \N__12510\,
            I => \N__12504\
        );

    \I__2904\ : InMux
    port map (
            O => \N__12507\,
            I => \N__12501\
        );

    \I__2903\ : LocalMux
    port map (
            O => \N__12504\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_7\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__12501\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_7\
        );

    \I__2901\ : InMux
    port map (
            O => \N__12496\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_6\
        );

    \I__2900\ : InMux
    port map (
            O => \N__12493\,
            I => \N__12489\
        );

    \I__2899\ : InMux
    port map (
            O => \N__12492\,
            I => \N__12486\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__12489\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_8\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__12486\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_8\
        );

    \I__2896\ : InMux
    port map (
            O => \N__12481\,
            I => \bfn_21_10_0_\
        );

    \I__2895\ : InMux
    port map (
            O => \N__12478\,
            I => \N__12475\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__12475\,
            I => \N__12472\
        );

    \I__2893\ : Span4Mux_s3_v
    port map (
            O => \N__12472\,
            I => \N__12469\
        );

    \I__2892\ : Odrv4
    port map (
            O => \N__12469\,
            I => \rTxBusReady_rep2_i_ess\
        );

    \I__2891\ : IoInMux
    port map (
            O => \N__12466\,
            I => \N__12463\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__12463\,
            I => \N__12460\
        );

    \I__2889\ : Span4Mux_s1_v
    port map (
            O => \N__12460\,
            I => \N__12457\
        );

    \I__2888\ : Odrv4
    port map (
            O => \N__12457\,
            I => \N_1241_i\
        );

    \I__2887\ : InMux
    port map (
            O => \N__12454\,
            I => \N__12451\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__12451\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_9\
        );

    \I__2885\ : CascadeMux
    port map (
            O => \N__12448\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_6_cascade_\
        );

    \I__2884\ : CascadeMux
    port map (
            O => \N__12445\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0_cascade_\
        );

    \I__2883\ : CascadeMux
    port map (
            O => \N__12442\,
            I => \N__12434\
        );

    \I__2882\ : CascadeMux
    port map (
            O => \N__12441\,
            I => \N__12429\
        );

    \I__2881\ : CascadeMux
    port map (
            O => \N__12440\,
            I => \N__12425\
        );

    \I__2880\ : InMux
    port map (
            O => \N__12439\,
            I => \N__12418\
        );

    \I__2879\ : InMux
    port map (
            O => \N__12438\,
            I => \N__12415\
        );

    \I__2878\ : InMux
    port map (
            O => \N__12437\,
            I => \N__12410\
        );

    \I__2877\ : InMux
    port map (
            O => \N__12434\,
            I => \N__12410\
        );

    \I__2876\ : InMux
    port map (
            O => \N__12433\,
            I => \N__12407\
        );

    \I__2875\ : InMux
    port map (
            O => \N__12432\,
            I => \N__12404\
        );

    \I__2874\ : InMux
    port map (
            O => \N__12429\,
            I => \N__12401\
        );

    \I__2873\ : InMux
    port map (
            O => \N__12428\,
            I => \N__12398\
        );

    \I__2872\ : InMux
    port map (
            O => \N__12425\,
            I => \N__12395\
        );

    \I__2871\ : InMux
    port map (
            O => \N__12424\,
            I => \N__12392\
        );

    \I__2870\ : InMux
    port map (
            O => \N__12423\,
            I => \N__12389\
        );

    \I__2869\ : InMux
    port map (
            O => \N__12422\,
            I => \N__12386\
        );

    \I__2868\ : InMux
    port map (
            O => \N__12421\,
            I => \N__12383\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__12418\,
            I => \N__12380\
        );

    \I__2866\ : LocalMux
    port map (
            O => \N__12415\,
            I => \N__12377\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__12410\,
            I => \N__12372\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__12407\,
            I => \N__12369\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__12404\,
            I => \N__12366\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__12401\,
            I => \N__12363\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__12398\,
            I => \N__12360\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__12395\,
            I => \N__12357\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__12392\,
            I => \N__12354\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__12389\,
            I => \N__12350\
        );

    \I__2857\ : LocalMux
    port map (
            O => \N__12386\,
            I => \N__12347\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__12383\,
            I => \N__12341\
        );

    \I__2855\ : Glb2LocalMux
    port map (
            O => \N__12380\,
            I => \N__12301\
        );

    \I__2854\ : Glb2LocalMux
    port map (
            O => \N__12377\,
            I => \N__12301\
        );

    \I__2853\ : CEMux
    port map (
            O => \N__12376\,
            I => \N__12301\
        );

    \I__2852\ : CEMux
    port map (
            O => \N__12375\,
            I => \N__12301\
        );

    \I__2851\ : Glb2LocalMux
    port map (
            O => \N__12372\,
            I => \N__12301\
        );

    \I__2850\ : Glb2LocalMux
    port map (
            O => \N__12369\,
            I => \N__12301\
        );

    \I__2849\ : Glb2LocalMux
    port map (
            O => \N__12366\,
            I => \N__12301\
        );

    \I__2848\ : Glb2LocalMux
    port map (
            O => \N__12363\,
            I => \N__12301\
        );

    \I__2847\ : Glb2LocalMux
    port map (
            O => \N__12360\,
            I => \N__12301\
        );

    \I__2846\ : Glb2LocalMux
    port map (
            O => \N__12357\,
            I => \N__12301\
        );

    \I__2845\ : Glb2LocalMux
    port map (
            O => \N__12354\,
            I => \N__12301\
        );

    \I__2844\ : CEMux
    port map (
            O => \N__12353\,
            I => \N__12301\
        );

    \I__2843\ : Glb2LocalMux
    port map (
            O => \N__12350\,
            I => \N__12301\
        );

    \I__2842\ : Glb2LocalMux
    port map (
            O => \N__12347\,
            I => \N__12301\
        );

    \I__2841\ : CEMux
    port map (
            O => \N__12346\,
            I => \N__12301\
        );

    \I__2840\ : CEMux
    port map (
            O => \N__12345\,
            I => \N__12301\
        );

    \I__2839\ : CEMux
    port map (
            O => \N__12344\,
            I => \N__12301\
        );

    \I__2838\ : Glb2LocalMux
    port map (
            O => \N__12341\,
            I => \N__12301\
        );

    \I__2837\ : CEMux
    port map (
            O => \N__12340\,
            I => \N__12301\
        );

    \I__2836\ : GlobalMux
    port map (
            O => \N__12301\,
            I => \N__12298\
        );

    \I__2835\ : gio2CtrlBuf
    port map (
            O => \N__12298\,
            I => \wPllLocked_g\
        );

    \I__2834\ : InMux
    port map (
            O => \N__12295\,
            I => \N__12292\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__12292\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_8\
        );

    \I__2832\ : InMux
    port map (
            O => \N__12289\,
            I => \N__12286\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__12286\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_7\
        );

    \I__2830\ : InMux
    port map (
            O => \N__12283\,
            I => \N__12278\
        );

    \I__2829\ : InMux
    port map (
            O => \N__12282\,
            I => \N__12275\
        );

    \I__2828\ : InMux
    port map (
            O => \N__12281\,
            I => \N__12272\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__12278\,
            I => \N__12269\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__12275\,
            I => \N__12266\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__12272\,
            I => \N__12263\
        );

    \I__2824\ : Span4Mux_v
    port map (
            O => \N__12269\,
            I => \N__12260\
        );

    \I__2823\ : Span4Mux_h
    port map (
            O => \N__12266\,
            I => \N__12257\
        );

    \I__2822\ : Odrv4
    port map (
            O => \N__12263\,
            I => \DUT.uart_inst0.N_77\
        );

    \I__2821\ : Odrv4
    port map (
            O => \N__12260\,
            I => \DUT.uart_inst0.N_77\
        );

    \I__2820\ : Odrv4
    port map (
            O => \N__12257\,
            I => \DUT.uart_inst0.N_77\
        );

    \I__2819\ : CascadeMux
    port map (
            O => \N__12250\,
            I => \N__12240\
        );

    \I__2818\ : InMux
    port map (
            O => \N__12249\,
            I => \N__12237\
        );

    \I__2817\ : CascadeMux
    port map (
            O => \N__12248\,
            I => \N__12234\
        );

    \I__2816\ : CascadeMux
    port map (
            O => \N__12247\,
            I => \N__12231\
        );

    \I__2815\ : InMux
    port map (
            O => \N__12246\,
            I => \N__12225\
        );

    \I__2814\ : InMux
    port map (
            O => \N__12245\,
            I => \N__12225\
        );

    \I__2813\ : InMux
    port map (
            O => \N__12244\,
            I => \N__12218\
        );

    \I__2812\ : InMux
    port map (
            O => \N__12243\,
            I => \N__12218\
        );

    \I__2811\ : InMux
    port map (
            O => \N__12240\,
            I => \N__12215\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__12237\,
            I => \N__12212\
        );

    \I__2809\ : InMux
    port map (
            O => \N__12234\,
            I => \N__12205\
        );

    \I__2808\ : InMux
    port map (
            O => \N__12231\,
            I => \N__12205\
        );

    \I__2807\ : InMux
    port map (
            O => \N__12230\,
            I => \N__12205\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__12225\,
            I => \N__12202\
        );

    \I__2805\ : InMux
    port map (
            O => \N__12224\,
            I => \N__12197\
        );

    \I__2804\ : InMux
    port map (
            O => \N__12223\,
            I => \N__12197\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__12218\,
            I => \N__12193\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__12215\,
            I => \N__12190\
        );

    \I__2801\ : Span4Mux_h
    port map (
            O => \N__12212\,
            I => \N__12187\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__12205\,
            I => \N__12180\
        );

    \I__2799\ : Span4Mux_v
    port map (
            O => \N__12202\,
            I => \N__12180\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__12197\,
            I => \N__12180\
        );

    \I__2797\ : InMux
    port map (
            O => \N__12196\,
            I => \N__12177\
        );

    \I__2796\ : Span4Mux_h
    port map (
            O => \N__12193\,
            I => \N__12174\
        );

    \I__2795\ : Odrv12
    port map (
            O => \N__12190\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0\
        );

    \I__2794\ : Odrv4
    port map (
            O => \N__12187\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0\
        );

    \I__2793\ : Odrv4
    port map (
            O => \N__12180\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__12177\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0\
        );

    \I__2791\ : Odrv4
    port map (
            O => \N__12174\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0\
        );

    \I__2790\ : CascadeMux
    port map (
            O => \N__12163\,
            I => \N__12159\
        );

    \I__2789\ : InMux
    port map (
            O => \N__12162\,
            I => \N__12154\
        );

    \I__2788\ : InMux
    port map (
            O => \N__12159\,
            I => \N__12147\
        );

    \I__2787\ : InMux
    port map (
            O => \N__12158\,
            I => \N__12147\
        );

    \I__2786\ : InMux
    port map (
            O => \N__12157\,
            I => \N__12147\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__12154\,
            I => \N__12142\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__12147\,
            I => \N__12142\
        );

    \I__2783\ : Odrv4
    port map (
            O => \N__12142\,
            I => \DUT.uart_inst0.N_147\
        );

    \I__2782\ : CascadeMux
    port map (
            O => \N__12139\,
            I => \N__12136\
        );

    \I__2781\ : InMux
    port map (
            O => \N__12136\,
            I => \N__12127\
        );

    \I__2780\ : InMux
    port map (
            O => \N__12135\,
            I => \N__12127\
        );

    \I__2779\ : InMux
    port map (
            O => \N__12134\,
            I => \N__12124\
        );

    \I__2778\ : InMux
    port map (
            O => \N__12133\,
            I => \N__12119\
        );

    \I__2777\ : InMux
    port map (
            O => \N__12132\,
            I => \N__12119\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__12127\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_2\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__12124\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_2\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__12119\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_2\
        );

    \I__2773\ : CascadeMux
    port map (
            O => \N__12112\,
            I => \DUT.uart_inst0.tx_countdown_0_c4_cascade_\
        );

    \I__2772\ : InMux
    port map (
            O => \N__12109\,
            I => \N__12106\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__12106\,
            I => \DUT.uart_inst0.tx_countdown_7_ns_1_4\
        );

    \I__2770\ : CascadeMux
    port map (
            O => \N__12103\,
            I => \DUT.uart_inst0.tx_countdown_7_ns_1_1_cascade_\
        );

    \I__2769\ : CascadeMux
    port map (
            O => \N__12100\,
            I => \N__12097\
        );

    \I__2768\ : InMux
    port map (
            O => \N__12097\,
            I => \N__12094\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__12094\,
            I => \DUT.uart_inst0.tx_countdown_0_c4\
        );

    \I__2766\ : InMux
    port map (
            O => \N__12091\,
            I => \N__12088\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__12088\,
            I => \DUT.uart_inst0.tx_countdown_7_ns_1_5\
        );

    \I__2764\ : InMux
    port map (
            O => \N__12085\,
            I => \N__12075\
        );

    \I__2763\ : InMux
    port map (
            O => \N__12084\,
            I => \N__12070\
        );

    \I__2762\ : InMux
    port map (
            O => \N__12083\,
            I => \N__12070\
        );

    \I__2761\ : InMux
    port map (
            O => \N__12082\,
            I => \N__12063\
        );

    \I__2760\ : InMux
    port map (
            O => \N__12081\,
            I => \N__12063\
        );

    \I__2759\ : InMux
    port map (
            O => \N__12080\,
            I => \N__12063\
        );

    \I__2758\ : InMux
    port map (
            O => \N__12079\,
            I => \N__12058\
        );

    \I__2757\ : InMux
    port map (
            O => \N__12078\,
            I => \N__12058\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__12075\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__12070\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__2754\ : LocalMux
    port map (
            O => \N__12063\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__12058\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__2752\ : CascadeMux
    port map (
            O => \N__12049\,
            I => \N__12039\
        );

    \I__2751\ : InMux
    port map (
            O => \N__12048\,
            I => \N__12034\
        );

    \I__2750\ : InMux
    port map (
            O => \N__12047\,
            I => \N__12034\
        );

    \I__2749\ : InMux
    port map (
            O => \N__12046\,
            I => \N__12029\
        );

    \I__2748\ : InMux
    port map (
            O => \N__12045\,
            I => \N__12029\
        );

    \I__2747\ : InMux
    port map (
            O => \N__12044\,
            I => \N__12024\
        );

    \I__2746\ : InMux
    port map (
            O => \N__12043\,
            I => \N__12024\
        );

    \I__2745\ : InMux
    port map (
            O => \N__12042\,
            I => \N__12019\
        );

    \I__2744\ : InMux
    port map (
            O => \N__12039\,
            I => \N__12019\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__12034\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__2742\ : LocalMux
    port map (
            O => \N__12029\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__12024\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__12019\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__2739\ : CascadeMux
    port map (
            O => \N__12010\,
            I => \N__12003\
        );

    \I__2738\ : InMux
    port map (
            O => \N__12009\,
            I => \N__12000\
        );

    \I__2737\ : InMux
    port map (
            O => \N__12008\,
            I => \N__11995\
        );

    \I__2736\ : InMux
    port map (
            O => \N__12007\,
            I => \N__11995\
        );

    \I__2735\ : InMux
    port map (
            O => \N__12006\,
            I => \N__11990\
        );

    \I__2734\ : InMux
    port map (
            O => \N__12003\,
            I => \N__11990\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__12000\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_5\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__11995\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_5\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__11990\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_5\
        );

    \I__2730\ : CascadeMux
    port map (
            O => \N__11983\,
            I => \DUT.uart_inst0.tx_countdown_7_m1_0_o2_1_2_cascade_\
        );

    \I__2729\ : InMux
    port map (
            O => \N__11980\,
            I => \N__11972\
        );

    \I__2728\ : InMux
    port map (
            O => \N__11979\,
            I => \N__11965\
        );

    \I__2727\ : InMux
    port map (
            O => \N__11978\,
            I => \N__11965\
        );

    \I__2726\ : InMux
    port map (
            O => \N__11977\,
            I => \N__11965\
        );

    \I__2725\ : InMux
    port map (
            O => \N__11976\,
            I => \N__11960\
        );

    \I__2724\ : InMux
    port map (
            O => \N__11975\,
            I => \N__11960\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__11972\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_4\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__11965\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_4\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__11960\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_4\
        );

    \I__2720\ : InMux
    port map (
            O => \N__11953\,
            I => \N__11950\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__11950\,
            I => \N__11947\
        );

    \I__2718\ : Odrv4
    port map (
            O => \N__11947\,
            I => \DUT.uart_inst0.N_68\
        );

    \I__2717\ : InMux
    port map (
            O => \N__11944\,
            I => \N__11935\
        );

    \I__2716\ : InMux
    port map (
            O => \N__11943\,
            I => \N__11935\
        );

    \I__2715\ : InMux
    port map (
            O => \N__11942\,
            I => \N__11935\
        );

    \I__2714\ : LocalMux
    port map (
            O => \N__11935\,
            I => \N__11932\
        );

    \I__2713\ : Span4Mux_h
    port map (
            O => \N__11932\,
            I => \N__11929\
        );

    \I__2712\ : Odrv4
    port map (
            O => \N__11929\,
            I => \DUT.uart_inst0.N_146\
        );

    \I__2711\ : CascadeMux
    port map (
            O => \N__11926\,
            I => \N__11922\
        );

    \I__2710\ : InMux
    port map (
            O => \N__11925\,
            I => \N__11914\
        );

    \I__2709\ : InMux
    port map (
            O => \N__11922\,
            I => \N__11911\
        );

    \I__2708\ : InMux
    port map (
            O => \N__11921\,
            I => \N__11902\
        );

    \I__2707\ : InMux
    port map (
            O => \N__11920\,
            I => \N__11902\
        );

    \I__2706\ : InMux
    port map (
            O => \N__11919\,
            I => \N__11902\
        );

    \I__2705\ : InMux
    port map (
            O => \N__11918\,
            I => \N__11902\
        );

    \I__2704\ : InMux
    port map (
            O => \N__11917\,
            I => \N__11899\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__11914\,
            I => \DUT.uart_inst0.tx_countdown_7_sm0_0\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__11911\,
            I => \DUT.uart_inst0.tx_countdown_7_sm0_0\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__11902\,
            I => \DUT.uart_inst0.tx_countdown_7_sm0_0\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__11899\,
            I => \DUT.uart_inst0.tx_countdown_7_sm0_0\
        );

    \I__2699\ : InMux
    port map (
            O => \N__11890\,
            I => \N__11887\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__11887\,
            I => \DUT.uart_inst0.tx_countdown_7_ns_1_3\
        );

    \I__2697\ : CascadeMux
    port map (
            O => \N__11884\,
            I => \N__11879\
        );

    \I__2696\ : CascadeMux
    port map (
            O => \N__11883\,
            I => \N__11876\
        );

    \I__2695\ : InMux
    port map (
            O => \N__11882\,
            I => \N__11870\
        );

    \I__2694\ : InMux
    port map (
            O => \N__11879\,
            I => \N__11867\
        );

    \I__2693\ : InMux
    port map (
            O => \N__11876\,
            I => \N__11862\
        );

    \I__2692\ : InMux
    port map (
            O => \N__11875\,
            I => \N__11862\
        );

    \I__2691\ : InMux
    port map (
            O => \N__11874\,
            I => \N__11857\
        );

    \I__2690\ : InMux
    port map (
            O => \N__11873\,
            I => \N__11857\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__11870\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__11867\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__11862\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__11857\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__2685\ : CascadeMux
    port map (
            O => \N__11848\,
            I => \DUT.uart_inst0.tx_state_RNI8CH01Z0Z_1_cascade_\
        );

    \I__2684\ : SRMux
    port map (
            O => \N__11845\,
            I => \N__11842\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__11842\,
            I => \DUT.uart_inst0.N_59_i\
        );

    \I__2682\ : InMux
    port map (
            O => \N__11839\,
            I => \N__11836\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__11836\,
            I => \N__11833\
        );

    \I__2680\ : Span4Mux_h
    port map (
            O => \N__11833\,
            I => \N__11829\
        );

    \I__2679\ : InMux
    port map (
            O => \N__11832\,
            I => \N__11826\
        );

    \I__2678\ : Odrv4
    port map (
            O => \N__11829\,
            I => \DUT.N_93\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__11826\,
            I => \DUT.N_93\
        );

    \I__2676\ : InMux
    port map (
            O => \N__11821\,
            I => \N__11815\
        );

    \I__2675\ : CascadeMux
    port map (
            O => \N__11820\,
            I => \N__11812\
        );

    \I__2674\ : CascadeMux
    port map (
            O => \N__11819\,
            I => \N__11809\
        );

    \I__2673\ : CascadeMux
    port map (
            O => \N__11818\,
            I => \N__11805\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__11815\,
            I => \N__11798\
        );

    \I__2671\ : InMux
    port map (
            O => \N__11812\,
            I => \N__11795\
        );

    \I__2670\ : InMux
    port map (
            O => \N__11809\,
            I => \N__11792\
        );

    \I__2669\ : InMux
    port map (
            O => \N__11808\,
            I => \N__11789\
        );

    \I__2668\ : InMux
    port map (
            O => \N__11805\,
            I => \N__11784\
        );

    \I__2667\ : InMux
    port map (
            O => \N__11804\,
            I => \N__11784\
        );

    \I__2666\ : InMux
    port map (
            O => \N__11803\,
            I => \N__11779\
        );

    \I__2665\ : InMux
    port map (
            O => \N__11802\,
            I => \N__11779\
        );

    \I__2664\ : InMux
    port map (
            O => \N__11801\,
            I => \N__11776\
        );

    \I__2663\ : Span4Mux_v
    port map (
            O => \N__11798\,
            I => \N__11773\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__11795\,
            I => \N__11764\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__11792\,
            I => \N__11764\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__11789\,
            I => \N__11764\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__11784\,
            I => \N__11764\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__11779\,
            I => \DUT.tx_state_1\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__11776\,
            I => \DUT.tx_state_1\
        );

    \I__2656\ : Odrv4
    port map (
            O => \N__11773\,
            I => \DUT.tx_state_1\
        );

    \I__2655\ : Odrv4
    port map (
            O => \N__11764\,
            I => \DUT.tx_state_1\
        );

    \I__2654\ : CascadeMux
    port map (
            O => \N__11755\,
            I => \N__11750\
        );

    \I__2653\ : InMux
    port map (
            O => \N__11754\,
            I => \N__11743\
        );

    \I__2652\ : InMux
    port map (
            O => \N__11753\,
            I => \N__11740\
        );

    \I__2651\ : InMux
    port map (
            O => \N__11750\,
            I => \N__11737\
        );

    \I__2650\ : InMux
    port map (
            O => \N__11749\,
            I => \N__11730\
        );

    \I__2649\ : InMux
    port map (
            O => \N__11748\,
            I => \N__11730\
        );

    \I__2648\ : InMux
    port map (
            O => \N__11747\,
            I => \N__11730\
        );

    \I__2647\ : InMux
    port map (
            O => \N__11746\,
            I => \N__11727\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__11743\,
            I => \N__11724\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__11740\,
            I => \N__11719\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__11737\,
            I => \N__11719\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__11730\,
            I => \N__11716\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__11727\,
            I => \N__11713\
        );

    \I__2641\ : Span4Mux_v
    port map (
            O => \N__11724\,
            I => \N__11708\
        );

    \I__2640\ : Span4Mux_v
    port map (
            O => \N__11719\,
            I => \N__11705\
        );

    \I__2639\ : Span4Mux_h
    port map (
            O => \N__11716\,
            I => \N__11702\
        );

    \I__2638\ : Span4Mux_h
    port map (
            O => \N__11713\,
            I => \N__11699\
        );

    \I__2637\ : InMux
    port map (
            O => \N__11712\,
            I => \N__11696\
        );

    \I__2636\ : InMux
    port map (
            O => \N__11711\,
            I => \N__11693\
        );

    \I__2635\ : Odrv4
    port map (
            O => \N__11708\,
            I => \DUT.rTransmitZ0\
        );

    \I__2634\ : Odrv4
    port map (
            O => \N__11705\,
            I => \DUT.rTransmitZ0\
        );

    \I__2633\ : Odrv4
    port map (
            O => \N__11702\,
            I => \DUT.rTransmitZ0\
        );

    \I__2632\ : Odrv4
    port map (
            O => \N__11699\,
            I => \DUT.rTransmitZ0\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__11696\,
            I => \DUT.rTransmitZ0\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__11693\,
            I => \DUT.rTransmitZ0\
        );

    \I__2629\ : CascadeMux
    port map (
            O => \N__11680\,
            I => \N__11671\
        );

    \I__2628\ : CascadeMux
    port map (
            O => \N__11679\,
            I => \N__11667\
        );

    \I__2627\ : CascadeMux
    port map (
            O => \N__11678\,
            I => \N__11662\
        );

    \I__2626\ : CascadeMux
    port map (
            O => \N__11677\,
            I => \N__11653\
        );

    \I__2625\ : CascadeMux
    port map (
            O => \N__11676\,
            I => \N__11648\
        );

    \I__2624\ : InMux
    port map (
            O => \N__11675\,
            I => \N__11641\
        );

    \I__2623\ : InMux
    port map (
            O => \N__11674\,
            I => \N__11641\
        );

    \I__2622\ : InMux
    port map (
            O => \N__11671\,
            I => \N__11641\
        );

    \I__2621\ : InMux
    port map (
            O => \N__11670\,
            I => \N__11636\
        );

    \I__2620\ : InMux
    port map (
            O => \N__11667\,
            I => \N__11636\
        );

    \I__2619\ : InMux
    port map (
            O => \N__11666\,
            I => \N__11625\
        );

    \I__2618\ : InMux
    port map (
            O => \N__11665\,
            I => \N__11625\
        );

    \I__2617\ : InMux
    port map (
            O => \N__11662\,
            I => \N__11625\
        );

    \I__2616\ : InMux
    port map (
            O => \N__11661\,
            I => \N__11625\
        );

    \I__2615\ : InMux
    port map (
            O => \N__11660\,
            I => \N__11625\
        );

    \I__2614\ : InMux
    port map (
            O => \N__11659\,
            I => \N__11614\
        );

    \I__2613\ : InMux
    port map (
            O => \N__11658\,
            I => \N__11614\
        );

    \I__2612\ : InMux
    port map (
            O => \N__11657\,
            I => \N__11614\
        );

    \I__2611\ : InMux
    port map (
            O => \N__11656\,
            I => \N__11614\
        );

    \I__2610\ : InMux
    port map (
            O => \N__11653\,
            I => \N__11614\
        );

    \I__2609\ : InMux
    port map (
            O => \N__11652\,
            I => \N__11607\
        );

    \I__2608\ : InMux
    port map (
            O => \N__11651\,
            I => \N__11607\
        );

    \I__2607\ : InMux
    port map (
            O => \N__11648\,
            I => \N__11607\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__11641\,
            I => \N__11604\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__11636\,
            I => \N__11595\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__11625\,
            I => \N__11595\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__11614\,
            I => \N__11595\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__11607\,
            I => \N__11592\
        );

    \I__2601\ : Span4Mux_v
    port map (
            O => \N__11604\,
            I => \N__11589\
        );

    \I__2600\ : InMux
    port map (
            O => \N__11603\,
            I => \N__11584\
        );

    \I__2599\ : InMux
    port map (
            O => \N__11602\,
            I => \N__11584\
        );

    \I__2598\ : Span4Mux_v
    port map (
            O => \N__11595\,
            I => \N__11581\
        );

    \I__2597\ : Span4Mux_h
    port map (
            O => \N__11592\,
            I => \N__11576\
        );

    \I__2596\ : Span4Mux_h
    port map (
            O => \N__11589\,
            I => \N__11576\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__11584\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__2594\ : Odrv4
    port map (
            O => \N__11581\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__2593\ : Odrv4
    port map (
            O => \N__11576\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__2592\ : InMux
    port map (
            O => \N__11569\,
            I => \N__11566\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__11566\,
            I => \DUT.fifo_tx_inst.un1_i11_2_i\
        );

    \I__2590\ : InMux
    port map (
            O => \N__11563\,
            I => \N__11554\
        );

    \I__2589\ : InMux
    port map (
            O => \N__11562\,
            I => \N__11554\
        );

    \I__2588\ : InMux
    port map (
            O => \N__11561\,
            I => \N__11554\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__11554\,
            I => \N__11551\
        );

    \I__2586\ : Span4Mux_h
    port map (
            O => \N__11551\,
            I => \N__11548\
        );

    \I__2585\ : Odrv4
    port map (
            O => \N__11548\,
            I => \DUT.fifo_tx_inst.rReadPtr11\
        );

    \I__2584\ : CascadeMux
    port map (
            O => \N__11545\,
            I => \DUT.fifo_tx_inst.un1_i11_2_i_cascade_\
        );

    \I__2583\ : InMux
    port map (
            O => \N__11542\,
            I => \N__11531\
        );

    \I__2582\ : InMux
    port map (
            O => \N__11541\,
            I => \N__11524\
        );

    \I__2581\ : InMux
    port map (
            O => \N__11540\,
            I => \N__11524\
        );

    \I__2580\ : InMux
    port map (
            O => \N__11539\,
            I => \N__11524\
        );

    \I__2579\ : InMux
    port map (
            O => \N__11538\,
            I => \N__11517\
        );

    \I__2578\ : InMux
    port map (
            O => \N__11537\,
            I => \N__11517\
        );

    \I__2577\ : InMux
    port map (
            O => \N__11536\,
            I => \N__11512\
        );

    \I__2576\ : InMux
    port map (
            O => \N__11535\,
            I => \N__11512\
        );

    \I__2575\ : CascadeMux
    port map (
            O => \N__11534\,
            I => \N__11508\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__11531\,
            I => \N__11504\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__11524\,
            I => \N__11501\
        );

    \I__2572\ : InMux
    port map (
            O => \N__11523\,
            I => \N__11496\
        );

    \I__2571\ : InMux
    port map (
            O => \N__11522\,
            I => \N__11496\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__11517\,
            I => \N__11491\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__11512\,
            I => \N__11491\
        );

    \I__2568\ : InMux
    port map (
            O => \N__11511\,
            I => \N__11488\
        );

    \I__2567\ : InMux
    port map (
            O => \N__11508\,
            I => \N__11483\
        );

    \I__2566\ : InMux
    port map (
            O => \N__11507\,
            I => \N__11483\
        );

    \I__2565\ : Span4Mux_h
    port map (
            O => \N__11504\,
            I => \N__11480\
        );

    \I__2564\ : Span4Mux_v
    port map (
            O => \N__11501\,
            I => \N__11475\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__11496\,
            I => \N__11475\
        );

    \I__2562\ : Span4Mux_h
    port map (
            O => \N__11491\,
            I => \N__11472\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__11488\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__11483\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__2559\ : Odrv4
    port map (
            O => \N__11480\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__2558\ : Odrv4
    port map (
            O => \N__11475\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__2557\ : Odrv4
    port map (
            O => \N__11472\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__2556\ : InMux
    port map (
            O => \N__11461\,
            I => \N__11456\
        );

    \I__2555\ : InMux
    port map (
            O => \N__11460\,
            I => \N__11453\
        );

    \I__2554\ : InMux
    port map (
            O => \N__11459\,
            I => \N__11450\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__11456\,
            I => \DUT.uart_inst0.N_74\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__11453\,
            I => \DUT.uart_inst0.N_74\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__11450\,
            I => \DUT.uart_inst0.N_74\
        );

    \I__2550\ : CascadeMux
    port map (
            O => \N__11443\,
            I => \N__11438\
        );

    \I__2549\ : CascadeMux
    port map (
            O => \N__11442\,
            I => \N__11429\
        );

    \I__2548\ : InMux
    port map (
            O => \N__11441\,
            I => \N__11424\
        );

    \I__2547\ : InMux
    port map (
            O => \N__11438\,
            I => \N__11419\
        );

    \I__2546\ : InMux
    port map (
            O => \N__11437\,
            I => \N__11412\
        );

    \I__2545\ : InMux
    port map (
            O => \N__11436\,
            I => \N__11412\
        );

    \I__2544\ : InMux
    port map (
            O => \N__11435\,
            I => \N__11412\
        );

    \I__2543\ : InMux
    port map (
            O => \N__11434\,
            I => \N__11409\
        );

    \I__2542\ : InMux
    port map (
            O => \N__11433\,
            I => \N__11399\
        );

    \I__2541\ : InMux
    port map (
            O => \N__11432\,
            I => \N__11399\
        );

    \I__2540\ : InMux
    port map (
            O => \N__11429\,
            I => \N__11399\
        );

    \I__2539\ : InMux
    port map (
            O => \N__11428\,
            I => \N__11396\
        );

    \I__2538\ : CascadeMux
    port map (
            O => \N__11427\,
            I => \N__11388\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__11424\,
            I => \N__11385\
        );

    \I__2536\ : InMux
    port map (
            O => \N__11423\,
            I => \N__11380\
        );

    \I__2535\ : InMux
    port map (
            O => \N__11422\,
            I => \N__11380\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__11419\,
            I => \N__11375\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__11412\,
            I => \N__11375\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__11409\,
            I => \N__11372\
        );

    \I__2531\ : InMux
    port map (
            O => \N__11408\,
            I => \N__11363\
        );

    \I__2530\ : InMux
    port map (
            O => \N__11407\,
            I => \N__11363\
        );

    \I__2529\ : InMux
    port map (
            O => \N__11406\,
            I => \N__11363\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__11399\,
            I => \N__11360\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__11396\,
            I => \N__11357\
        );

    \I__2526\ : InMux
    port map (
            O => \N__11395\,
            I => \N__11350\
        );

    \I__2525\ : InMux
    port map (
            O => \N__11394\,
            I => \N__11350\
        );

    \I__2524\ : InMux
    port map (
            O => \N__11393\,
            I => \N__11350\
        );

    \I__2523\ : InMux
    port map (
            O => \N__11392\,
            I => \N__11345\
        );

    \I__2522\ : InMux
    port map (
            O => \N__11391\,
            I => \N__11345\
        );

    \I__2521\ : InMux
    port map (
            O => \N__11388\,
            I => \N__11342\
        );

    \I__2520\ : Span12Mux_s10_v
    port map (
            O => \N__11385\,
            I => \N__11339\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__11380\,
            I => \N__11336\
        );

    \I__2518\ : Span4Mux_v
    port map (
            O => \N__11375\,
            I => \N__11331\
        );

    \I__2517\ : Span4Mux_h
    port map (
            O => \N__11372\,
            I => \N__11331\
        );

    \I__2516\ : InMux
    port map (
            O => \N__11371\,
            I => \N__11328\
        );

    \I__2515\ : InMux
    port map (
            O => \N__11370\,
            I => \N__11325\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__11363\,
            I => \N__11318\
        );

    \I__2513\ : Span4Mux_h
    port map (
            O => \N__11360\,
            I => \N__11318\
        );

    \I__2512\ : Span4Mux_h
    port map (
            O => \N__11357\,
            I => \N__11318\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__11350\,
            I => \N__11313\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__11345\,
            I => \N__11313\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__11342\,
            I => \DUT.tx_state_0\
        );

    \I__2508\ : Odrv12
    port map (
            O => \N__11339\,
            I => \DUT.tx_state_0\
        );

    \I__2507\ : Odrv4
    port map (
            O => \N__11336\,
            I => \DUT.tx_state_0\
        );

    \I__2506\ : Odrv4
    port map (
            O => \N__11331\,
            I => \DUT.tx_state_0\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__11328\,
            I => \DUT.tx_state_0\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__11325\,
            I => \DUT.tx_state_0\
        );

    \I__2503\ : Odrv4
    port map (
            O => \N__11318\,
            I => \DUT.tx_state_0\
        );

    \I__2502\ : Odrv12
    port map (
            O => \N__11313\,
            I => \DUT.tx_state_0\
        );

    \I__2501\ : InMux
    port map (
            O => \N__11296\,
            I => \N__11293\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__11293\,
            I => \DUT.uart_inst0.tx_countdown_7_1_2\
        );

    \I__2499\ : CascadeMux
    port map (
            O => \N__11290\,
            I => \N__11287\
        );

    \I__2498\ : InMux
    port map (
            O => \N__11287\,
            I => \N__11284\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__11284\,
            I => \DUT.uart_inst0.N_91\
        );

    \I__2496\ : InMux
    port map (
            O => \N__11281\,
            I => \N__11278\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__11278\,
            I => \rTxBusReady_rep1_i_ess\
        );

    \I__2494\ : InMux
    port map (
            O => \N__11275\,
            I => \N__11272\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__11272\,
            I => \N__11269\
        );

    \I__2492\ : Odrv12
    port map (
            O => \N__11269\,
            I => \rTxBusReady_rep3_i_ess\
        );

    \I__2491\ : InMux
    port map (
            O => \N__11266\,
            I => \N__11263\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__11263\,
            I => \N__11260\
        );

    \I__2489\ : Span4Mux_s3_v
    port map (
            O => \N__11260\,
            I => \N__11257\
        );

    \I__2488\ : Odrv4
    port map (
            O => \N__11257\,
            I => \rTxBusReady_rep0_i_ess\
        );

    \I__2487\ : InMux
    port map (
            O => \N__11254\,
            I => \N__11251\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__11251\,
            I => \N__11245\
        );

    \I__2485\ : InMux
    port map (
            O => \N__11250\,
            I => \N__11242\
        );

    \I__2484\ : CascadeMux
    port map (
            O => \N__11249\,
            I => \N__11236\
        );

    \I__2483\ : CascadeMux
    port map (
            O => \N__11248\,
            I => \N__11232\
        );

    \I__2482\ : Span4Mux_h
    port map (
            O => \N__11245\,
            I => \N__11227\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__11242\,
            I => \N__11227\
        );

    \I__2480\ : InMux
    port map (
            O => \N__11241\,
            I => \N__11224\
        );

    \I__2479\ : InMux
    port map (
            O => \N__11240\,
            I => \N__11215\
        );

    \I__2478\ : InMux
    port map (
            O => \N__11239\,
            I => \N__11215\
        );

    \I__2477\ : InMux
    port map (
            O => \N__11236\,
            I => \N__11215\
        );

    \I__2476\ : InMux
    port map (
            O => \N__11235\,
            I => \N__11215\
        );

    \I__2475\ : InMux
    port map (
            O => \N__11232\,
            I => \N__11212\
        );

    \I__2474\ : Span4Mux_v
    port map (
            O => \N__11227\,
            I => \N__11209\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__11224\,
            I => \N__11206\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__11215\,
            I => \N__11201\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__11212\,
            I => \N__11201\
        );

    \I__2470\ : Sp12to4
    port map (
            O => \N__11209\,
            I => \N__11198\
        );

    \I__2469\ : Span4Mux_h
    port map (
            O => \N__11206\,
            I => \N__11195\
        );

    \I__2468\ : Span12Mux_v
    port map (
            O => \N__11201\,
            I => \N__11188\
        );

    \I__2467\ : Span12Mux_s7_h
    port map (
            O => \N__11198\,
            I => \N__11188\
        );

    \I__2466\ : Sp12to4
    port map (
            O => \N__11195\,
            I => \N__11188\
        );

    \I__2465\ : Span12Mux_v
    port map (
            O => \N__11188\,
            I => \N__11185\
        );

    \I__2464\ : Odrv12
    port map (
            O => \N__11185\,
            I => \iTxE_n_c\
        );

    \I__2463\ : InMux
    port map (
            O => \N__11182\,
            I => \N__11178\
        );

    \I__2462\ : InMux
    port map (
            O => \N__11181\,
            I => \N__11175\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__11178\,
            I => \N__11172\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__11175\,
            I => \N__11167\
        );

    \I__2459\ : Span4Mux_h
    port map (
            O => \N__11172\,
            I => \N__11164\
        );

    \I__2458\ : InMux
    port map (
            O => \N__11171\,
            I => \N__11159\
        );

    \I__2457\ : InMux
    port map (
            O => \N__11170\,
            I => \N__11159\
        );

    \I__2456\ : Span12Mux_s9_v
    port map (
            O => \N__11167\,
            I => \N__11156\
        );

    \I__2455\ : Odrv4
    port map (
            O => \N__11164\,
            I => \fifo_inst.ftdi_output_inst.N_68_0\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__11159\,
            I => \fifo_inst.ftdi_output_inst.N_68_0\
        );

    \I__2453\ : Odrv12
    port map (
            O => \N__11156\,
            I => \fifo_inst.ftdi_output_inst.N_68_0\
        );

    \I__2452\ : InMux
    port map (
            O => \N__11149\,
            I => \N__11143\
        );

    \I__2451\ : InMux
    port map (
            O => \N__11148\,
            I => \N__11138\
        );

    \I__2450\ : InMux
    port map (
            O => \N__11147\,
            I => \N__11138\
        );

    \I__2449\ : InMux
    port map (
            O => \N__11146\,
            I => \N__11135\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__11143\,
            I => \N__11131\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__11138\,
            I => \N__11126\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__11135\,
            I => \N__11120\
        );

    \I__2445\ : SRMux
    port map (
            O => \N__11134\,
            I => \N__11074\
        );

    \I__2444\ : Glb2LocalMux
    port map (
            O => \N__11131\,
            I => \N__11074\
        );

    \I__2443\ : SRMux
    port map (
            O => \N__11130\,
            I => \N__11074\
        );

    \I__2442\ : SRMux
    port map (
            O => \N__11129\,
            I => \N__11074\
        );

    \I__2441\ : Glb2LocalMux
    port map (
            O => \N__11126\,
            I => \N__11074\
        );

    \I__2440\ : SRMux
    port map (
            O => \N__11125\,
            I => \N__11074\
        );

    \I__2439\ : SRMux
    port map (
            O => \N__11124\,
            I => \N__11074\
        );

    \I__2438\ : SRMux
    port map (
            O => \N__11123\,
            I => \N__11074\
        );

    \I__2437\ : Glb2LocalMux
    port map (
            O => \N__11120\,
            I => \N__11074\
        );

    \I__2436\ : SRMux
    port map (
            O => \N__11119\,
            I => \N__11074\
        );

    \I__2435\ : SRMux
    port map (
            O => \N__11118\,
            I => \N__11074\
        );

    \I__2434\ : SRMux
    port map (
            O => \N__11117\,
            I => \N__11074\
        );

    \I__2433\ : SRMux
    port map (
            O => \N__11116\,
            I => \N__11074\
        );

    \I__2432\ : SRMux
    port map (
            O => \N__11115\,
            I => \N__11074\
        );

    \I__2431\ : SRMux
    port map (
            O => \N__11114\,
            I => \N__11074\
        );

    \I__2430\ : SRMux
    port map (
            O => \N__11113\,
            I => \N__11074\
        );

    \I__2429\ : SRMux
    port map (
            O => \N__11112\,
            I => \N__11074\
        );

    \I__2428\ : SRMux
    port map (
            O => \N__11111\,
            I => \N__11074\
        );

    \I__2427\ : GlobalMux
    port map (
            O => \N__11074\,
            I => \N__11071\
        );

    \I__2426\ : gio2CtrlBuf
    port map (
            O => \N__11071\,
            I => \wPllLocked_i_g\
        );

    \I__2425\ : CascadeMux
    port map (
            O => \N__11068\,
            I => \fifo_inst.ftdi_output_inst.un1_oTx_n_1_sqmuxa_0_i_cascade_\
        );

    \I__2424\ : CEMux
    port map (
            O => \N__11065\,
            I => \N__11062\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__11062\,
            I => \fifo_inst.ftdi_output_inst.un1_oTx_n_1_sqmuxa_0_i_0\
        );

    \I__2422\ : InMux
    port map (
            O => \N__11059\,
            I => \N__11056\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__11056\,
            I => \N__11051\
        );

    \I__2420\ : InMux
    port map (
            O => \N__11055\,
            I => \N__11048\
        );

    \I__2419\ : InMux
    port map (
            O => \N__11054\,
            I => \N__11045\
        );

    \I__2418\ : Span4Mux_v
    port map (
            O => \N__11051\,
            I => \N__11031\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__11048\,
            I => \N__11031\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__11045\,
            I => \N__11031\
        );

    \I__2415\ : InMux
    port map (
            O => \N__11044\,
            I => \N__11028\
        );

    \I__2414\ : InMux
    port map (
            O => \N__11043\,
            I => \N__11019\
        );

    \I__2413\ : InMux
    port map (
            O => \N__11042\,
            I => \N__11019\
        );

    \I__2412\ : InMux
    port map (
            O => \N__11041\,
            I => \N__11019\
        );

    \I__2411\ : InMux
    port map (
            O => \N__11040\,
            I => \N__11019\
        );

    \I__2410\ : InMux
    port map (
            O => \N__11039\,
            I => \N__11016\
        );

    \I__2409\ : InMux
    port map (
            O => \N__11038\,
            I => \N__11013\
        );

    \I__2408\ : Span4Mux_v
    port map (
            O => \N__11031\,
            I => \N__11010\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__11028\,
            I => \N__11007\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__11019\,
            I => \N__11000\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__11016\,
            I => \N__11000\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__11013\,
            I => \N__11000\
        );

    \I__2403\ : Sp12to4
    port map (
            O => \N__11010\,
            I => \N__10997\
        );

    \I__2402\ : Span4Mux_h
    port map (
            O => \N__11007\,
            I => \N__10994\
        );

    \I__2401\ : Span12Mux_v
    port map (
            O => \N__11000\,
            I => \N__10991\
        );

    \I__2400\ : Span12Mux_h
    port map (
            O => \N__10997\,
            I => \N__10986\
        );

    \I__2399\ : Sp12to4
    port map (
            O => \N__10994\,
            I => \N__10986\
        );

    \I__2398\ : Span12Mux_v
    port map (
            O => \N__10991\,
            I => \N__10983\
        );

    \I__2397\ : Span12Mux_v
    port map (
            O => \N__10986\,
            I => \N__10980\
        );

    \I__2396\ : Odrv12
    port map (
            O => \N__10983\,
            I => \iRxF_n_c\
        );

    \I__2395\ : Odrv12
    port map (
            O => \N__10980\,
            I => \iRxF_n_c\
        );

    \I__2394\ : InMux
    port map (
            O => \N__10975\,
            I => \N__10966\
        );

    \I__2393\ : InMux
    port map (
            O => \N__10974\,
            I => \N__10957\
        );

    \I__2392\ : InMux
    port map (
            O => \N__10973\,
            I => \N__10957\
        );

    \I__2391\ : InMux
    port map (
            O => \N__10972\,
            I => \N__10957\
        );

    \I__2390\ : InMux
    port map (
            O => \N__10971\,
            I => \N__10957\
        );

    \I__2389\ : InMux
    port map (
            O => \N__10970\,
            I => \N__10953\
        );

    \I__2388\ : InMux
    port map (
            O => \N__10969\,
            I => \N__10950\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__10966\,
            I => \N__10947\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__10957\,
            I => \N__10943\
        );

    \I__2385\ : InMux
    port map (
            O => \N__10956\,
            I => \N__10940\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__10953\,
            I => \N__10934\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__10950\,
            I => \N__10934\
        );

    \I__2382\ : Span4Mux_h
    port map (
            O => \N__10947\,
            I => \N__10931\
        );

    \I__2381\ : InMux
    port map (
            O => \N__10946\,
            I => \N__10928\
        );

    \I__2380\ : Span4Mux_v
    port map (
            O => \N__10943\,
            I => \N__10923\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__10940\,
            I => \N__10923\
        );

    \I__2378\ : InMux
    port map (
            O => \N__10939\,
            I => \N__10920\
        );

    \I__2377\ : Span4Mux_h
    port map (
            O => \N__10934\,
            I => \N__10917\
        );

    \I__2376\ : Odrv4
    port map (
            O => \N__10931\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__10928\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0\
        );

    \I__2374\ : Odrv4
    port map (
            O => \N__10923\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__10920\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0\
        );

    \I__2372\ : Odrv4
    port map (
            O => \N__10917\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0\
        );

    \I__2371\ : InMux
    port map (
            O => \N__10906\,
            I => \N__10903\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__10903\,
            I => \fifo_inst.ftdi_output_inst.N_80\
        );

    \I__2369\ : CascadeMux
    port map (
            O => \N__10900\,
            I => \DUT.uart_inst0.N_77_cascade_\
        );

    \I__2368\ : InMux
    port map (
            O => \N__10897\,
            I => \N__10894\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__10894\,
            I => \DUT.uart_inst0.tx_state_RNI8CH01Z0Z_1\
        );

    \I__2366\ : CascadeMux
    port map (
            O => \N__10891\,
            I => \DUT.uart_inst0.tx_state_ns_i_i_o2_a0_3_0_cascade_\
        );

    \I__2365\ : CascadeMux
    port map (
            O => \N__10888\,
            I => \N__10884\
        );

    \I__2364\ : InMux
    port map (
            O => \N__10887\,
            I => \N__10880\
        );

    \I__2363\ : InMux
    port map (
            O => \N__10884\,
            I => \N__10875\
        );

    \I__2362\ : InMux
    port map (
            O => \N__10883\,
            I => \N__10875\
        );

    \I__2361\ : LocalMux
    port map (
            O => \N__10880\,
            I => \DUT.uart_inst0.N_69_i\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__10875\,
            I => \DUT.uart_inst0.N_69_i\
        );

    \I__2359\ : CascadeMux
    port map (
            O => \N__10870\,
            I => \DUT.uart_inst0.tx_countdown_30_3_cascade_\
        );

    \I__2358\ : InMux
    port map (
            O => \N__10867\,
            I => \N__10864\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__10864\,
            I => \N__10861\
        );

    \I__2356\ : Span4Mux_h
    port map (
            O => \N__10861\,
            I => \N__10856\
        );

    \I__2355\ : InMux
    port map (
            O => \N__10860\,
            I => \N__10853\
        );

    \I__2354\ : InMux
    port map (
            O => \N__10859\,
            I => \N__10849\
        );

    \I__2353\ : Span4Mux_v
    port map (
            O => \N__10856\,
            I => \N__10846\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__10853\,
            I => \N__10843\
        );

    \I__2351\ : InMux
    port map (
            O => \N__10852\,
            I => \N__10840\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__10849\,
            I => \N__10837\
        );

    \I__2349\ : Odrv4
    port map (
            O => \N__10846\,
            I => \DUT.uart_inst0.N_84\
        );

    \I__2348\ : Odrv4
    port map (
            O => \N__10843\,
            I => \DUT.uart_inst0.N_84\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__10840\,
            I => \DUT.uart_inst0.N_84\
        );

    \I__2346\ : Odrv4
    port map (
            O => \N__10837\,
            I => \DUT.uart_inst0.N_84\
        );

    \I__2345\ : InMux
    port map (
            O => \N__10828\,
            I => \N__10822\
        );

    \I__2344\ : InMux
    port map (
            O => \N__10827\,
            I => \N__10822\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__10822\,
            I => \DUT.uart_inst0.N_30_1\
        );

    \I__2342\ : IoInMux
    port map (
            O => \N__10819\,
            I => \N__10816\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__10816\,
            I => \N__10813\
        );

    \I__2340\ : Span4Mux_s0_v
    port map (
            O => \N__10813\,
            I => \N__10810\
        );

    \I__2339\ : Odrv4
    port map (
            O => \N__10810\,
            I => \N_1242_i\
        );

    \I__2338\ : IoInMux
    port map (
            O => \N__10807\,
            I => \N__10804\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__10804\,
            I => \N__10801\
        );

    \I__2336\ : Span4Mux_s2_v
    port map (
            O => \N__10801\,
            I => \N__10798\
        );

    \I__2335\ : Odrv4
    port map (
            O => \N__10798\,
            I => \N_1240_i\
        );

    \I__2334\ : InMux
    port map (
            O => \N__10795\,
            I => \N__10792\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__10792\,
            I => \N__10787\
        );

    \I__2332\ : InMux
    port map (
            O => \N__10791\,
            I => \N__10784\
        );

    \I__2331\ : InMux
    port map (
            O => \N__10790\,
            I => \N__10781\
        );

    \I__2330\ : Odrv12
    port map (
            O => \N__10787\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__10784\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__10781\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2\
        );

    \I__2327\ : CascadeMux
    port map (
            O => \N__10774\,
            I => \fifo_inst.ftdi_output_inst.N_78_cascade_\
        );

    \I__2326\ : InMux
    port map (
            O => \N__10771\,
            I => \N__10764\
        );

    \I__2325\ : InMux
    port map (
            O => \N__10770\,
            I => \N__10759\
        );

    \I__2324\ : InMux
    port map (
            O => \N__10769\,
            I => \N__10759\
        );

    \I__2323\ : InMux
    port map (
            O => \N__10768\,
            I => \N__10754\
        );

    \I__2322\ : InMux
    port map (
            O => \N__10767\,
            I => \N__10754\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__10764\,
            I => \DUT.uart_inst0.N_142\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__10759\,
            I => \DUT.uart_inst0.N_142\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__10754\,
            I => \DUT.uart_inst0.N_142\
        );

    \I__2318\ : InMux
    port map (
            O => \N__10747\,
            I => \N__10744\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__10744\,
            I => \DUT.uart_inst0.N_144\
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__10741\,
            I => \DUT.uart_inst0.N_74_cascade_\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__10738\,
            I => \N__10735\
        );

    \I__2314\ : InMux
    port map (
            O => \N__10735\,
            I => \N__10732\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__10732\,
            I => \DUT.uart_inst0.N_143\
        );

    \I__2312\ : CascadeMux
    port map (
            O => \N__10729\,
            I => \DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0_cascade_\
        );

    \I__2311\ : InMux
    port map (
            O => \N__10726\,
            I => \N__10722\
        );

    \I__2310\ : InMux
    port map (
            O => \N__10725\,
            I => \N__10718\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__10722\,
            I => \N__10715\
        );

    \I__2308\ : InMux
    port map (
            O => \N__10721\,
            I => \N__10712\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__10718\,
            I => \DUT.uart_inst0.N_75\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__10715\,
            I => \DUT.uart_inst0.N_75\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__10712\,
            I => \DUT.uart_inst0.N_75\
        );

    \I__2304\ : CascadeMux
    port map (
            O => \N__10705\,
            I => \DUT.uart_inst0.N_75_cascade_\
        );

    \I__2303\ : InMux
    port map (
            O => \N__10702\,
            I => \N__10699\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__10699\,
            I => \DUT.uart_inst0.tx_countdown_7s2_0_0\
        );

    \I__2301\ : InMux
    port map (
            O => \N__10696\,
            I => \N__10687\
        );

    \I__2300\ : InMux
    port map (
            O => \N__10695\,
            I => \N__10687\
        );

    \I__2299\ : InMux
    port map (
            O => \N__10694\,
            I => \N__10687\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__10687\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_2\
        );

    \I__2297\ : CascadeMux
    port map (
            O => \N__10684\,
            I => \N__10679\
        );

    \I__2296\ : CascadeMux
    port map (
            O => \N__10683\,
            I => \N__10676\
        );

    \I__2295\ : InMux
    port map (
            O => \N__10682\,
            I => \N__10666\
        );

    \I__2294\ : InMux
    port map (
            O => \N__10679\,
            I => \N__10666\
        );

    \I__2293\ : InMux
    port map (
            O => \N__10676\,
            I => \N__10666\
        );

    \I__2292\ : InMux
    port map (
            O => \N__10675\,
            I => \N__10666\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__10666\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_1\
        );

    \I__2290\ : InMux
    port map (
            O => \N__10663\,
            I => \N__10648\
        );

    \I__2289\ : InMux
    port map (
            O => \N__10662\,
            I => \N__10648\
        );

    \I__2288\ : InMux
    port map (
            O => \N__10661\,
            I => \N__10648\
        );

    \I__2287\ : InMux
    port map (
            O => \N__10660\,
            I => \N__10648\
        );

    \I__2286\ : InMux
    port map (
            O => \N__10659\,
            I => \N__10648\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__10648\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_0\
        );

    \I__2284\ : CascadeMux
    port map (
            O => \N__10645\,
            I => \DUT.uart_inst0.N_142_cascade_\
        );

    \I__2283\ : CascadeMux
    port map (
            O => \N__10642\,
            I => \N__10635\
        );

    \I__2282\ : InMux
    port map (
            O => \N__10641\,
            I => \N__10630\
        );

    \I__2281\ : CascadeMux
    port map (
            O => \N__10640\,
            I => \N__10627\
        );

    \I__2280\ : IoInMux
    port map (
            O => \N__10639\,
            I => \N__10622\
        );

    \I__2279\ : InMux
    port map (
            O => \N__10638\,
            I => \N__10619\
        );

    \I__2278\ : InMux
    port map (
            O => \N__10635\,
            I => \N__10616\
        );

    \I__2277\ : InMux
    port map (
            O => \N__10634\,
            I => \N__10613\
        );

    \I__2276\ : InMux
    port map (
            O => \N__10633\,
            I => \N__10610\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__10630\,
            I => \N__10607\
        );

    \I__2274\ : InMux
    port map (
            O => \N__10627\,
            I => \N__10604\
        );

    \I__2273\ : CascadeMux
    port map (
            O => \N__10626\,
            I => \N__10601\
        );

    \I__2272\ : InMux
    port map (
            O => \N__10625\,
            I => \N__10598\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__10622\,
            I => \N__10595\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__10619\,
            I => \N__10592\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__10616\,
            I => \N__10585\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__10613\,
            I => \N__10585\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__10610\,
            I => \N__10585\
        );

    \I__2266\ : Span4Mux_v
    port map (
            O => \N__10607\,
            I => \N__10582\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__10604\,
            I => \N__10579\
        );

    \I__2264\ : InMux
    port map (
            O => \N__10601\,
            I => \N__10576\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__10598\,
            I => \N__10573\
        );

    \I__2262\ : Span4Mux_s1_v
    port map (
            O => \N__10595\,
            I => \N__10570\
        );

    \I__2261\ : Span4Mux_v
    port map (
            O => \N__10592\,
            I => \N__10567\
        );

    \I__2260\ : Span4Mux_v
    port map (
            O => \N__10585\,
            I => \N__10564\
        );

    \I__2259\ : Span4Mux_h
    port map (
            O => \N__10582\,
            I => \N__10559\
        );

    \I__2258\ : Span4Mux_v
    port map (
            O => \N__10579\,
            I => \N__10559\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__10576\,
            I => \N__10556\
        );

    \I__2256\ : Span4Mux_v
    port map (
            O => \N__10573\,
            I => \N__10553\
        );

    \I__2255\ : Span4Mux_v
    port map (
            O => \N__10570\,
            I => \N__10546\
        );

    \I__2254\ : Span4Mux_h
    port map (
            O => \N__10567\,
            I => \N__10546\
        );

    \I__2253\ : Span4Mux_h
    port map (
            O => \N__10564\,
            I => \N__10546\
        );

    \I__2252\ : Span4Mux_h
    port map (
            O => \N__10559\,
            I => \N__10543\
        );

    \I__2251\ : Sp12to4
    port map (
            O => \N__10556\,
            I => \N__10540\
        );

    \I__2250\ : Span4Mux_h
    port map (
            O => \N__10553\,
            I => \N__10537\
        );

    \I__2249\ : Sp12to4
    port map (
            O => \N__10546\,
            I => \N__10532\
        );

    \I__2248\ : Sp12to4
    port map (
            O => \N__10543\,
            I => \N__10532\
        );

    \I__2247\ : Span12Mux_v
    port map (
            O => \N__10540\,
            I => \N__10529\
        );

    \I__2246\ : Sp12to4
    port map (
            O => \N__10537\,
            I => \N__10526\
        );

    \I__2245\ : Span12Mux_h
    port map (
            O => \N__10532\,
            I => \N__10523\
        );

    \I__2244\ : Span12Mux_h
    port map (
            O => \N__10529\,
            I => \N__10520\
        );

    \I__2243\ : Span12Mux_v
    port map (
            O => \N__10526\,
            I => \N__10517\
        );

    \I__2242\ : Span12Mux_v
    port map (
            O => \N__10523\,
            I => \N__10514\
        );

    \I__2241\ : Span12Mux_v
    port map (
            O => \N__10520\,
            I => \N__10509\
        );

    \I__2240\ : Span12Mux_h
    port map (
            O => \N__10517\,
            I => \N__10509\
        );

    \I__2239\ : Odrv12
    port map (
            O => \N__10514\,
            I => \wPllLocked\
        );

    \I__2238\ : Odrv12
    port map (
            O => \N__10509\,
            I => \wPllLocked\
        );

    \I__2237\ : CascadeMux
    port map (
            O => \N__10504\,
            I => \DUT.uart_inst0.N_84_cascade_\
        );

    \I__2236\ : CascadeMux
    port map (
            O => \N__10501\,
            I => \N__10498\
        );

    \I__2235\ : InMux
    port map (
            O => \N__10498\,
            I => \N__10486\
        );

    \I__2234\ : InMux
    port map (
            O => \N__10497\,
            I => \N__10486\
        );

    \I__2233\ : InMux
    port map (
            O => \N__10496\,
            I => \N__10486\
        );

    \I__2232\ : InMux
    port map (
            O => \N__10495\,
            I => \N__10486\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__10486\,
            I => \N__10483\
        );

    \I__2230\ : Odrv4
    port map (
            O => \N__10483\,
            I => \DUT.uart_inst0.N_22\
        );

    \I__2229\ : CascadeMux
    port map (
            O => \N__10480\,
            I => \DUT.uart_inst0.N_22_cascade_\
        );

    \I__2228\ : InMux
    port map (
            O => \N__10477\,
            I => \N__10474\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__10474\,
            I => \DUT.uart_inst0.un1_tx_bits_remaining_c3\
        );

    \I__2226\ : CascadeMux
    port map (
            O => \N__10471\,
            I => \N__10467\
        );

    \I__2225\ : InMux
    port map (
            O => \N__10470\,
            I => \N__10464\
        );

    \I__2224\ : InMux
    port map (
            O => \N__10467\,
            I => \N__10461\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__10464\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_3\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__10461\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_3\
        );

    \I__2221\ : InMux
    port map (
            O => \N__10456\,
            I => \N__10453\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__10453\,
            I => \N__10447\
        );

    \I__2219\ : InMux
    port map (
            O => \N__10452\,
            I => \N__10444\
        );

    \I__2218\ : InMux
    port map (
            O => \N__10451\,
            I => \N__10439\
        );

    \I__2217\ : InMux
    port map (
            O => \N__10450\,
            I => \N__10439\
        );

    \I__2216\ : Odrv12
    port map (
            O => \N__10447\,
            I => \rRxReadZ0\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__10444\,
            I => \rRxReadZ0\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__10439\,
            I => \rRxReadZ0\
        );

    \I__2213\ : InMux
    port map (
            O => \N__10432\,
            I => \N__10429\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__10429\,
            I => \N__10425\
        );

    \I__2211\ : InMux
    port map (
            O => \N__10428\,
            I => \N__10422\
        );

    \I__2210\ : Odrv12
    port map (
            O => \N__10425\,
            I => \DUT.fifo_rx_inst.N_206\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__10422\,
            I => \DUT.fifo_rx_inst.N_206\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__10417\,
            I => \N__10414\
        );

    \I__2207\ : InMux
    port map (
            O => \N__10414\,
            I => \N__10409\
        );

    \I__2206\ : CascadeMux
    port map (
            O => \N__10413\,
            I => \N__10405\
        );

    \I__2205\ : InMux
    port map (
            O => \N__10412\,
            I => \N__10400\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__10409\,
            I => \N__10397\
        );

    \I__2203\ : InMux
    port map (
            O => \N__10408\,
            I => \N__10392\
        );

    \I__2202\ : InMux
    port map (
            O => \N__10405\,
            I => \N__10392\
        );

    \I__2201\ : InMux
    port map (
            O => \N__10404\,
            I => \N__10389\
        );

    \I__2200\ : InMux
    port map (
            O => \N__10403\,
            I => \N__10386\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__10400\,
            I => \N__10377\
        );

    \I__2198\ : Span4Mux_v
    port map (
            O => \N__10397\,
            I => \N__10377\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__10392\,
            I => \N__10377\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__10389\,
            I => \N__10377\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__10386\,
            I => \N__10372\
        );

    \I__2194\ : Span4Mux_h
    port map (
            O => \N__10377\,
            I => \N__10372\
        );

    \I__2193\ : Odrv4
    port map (
            O => \N__10372\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_0\
        );

    \I__2192\ : InMux
    port map (
            O => \N__10369\,
            I => \N__10364\
        );

    \I__2191\ : InMux
    port map (
            O => \N__10368\,
            I => \N__10359\
        );

    \I__2190\ : InMux
    port map (
            O => \N__10367\,
            I => \N__10359\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__10364\,
            I => \N__10356\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__10359\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1\
        );

    \I__2187\ : Odrv12
    port map (
            O => \N__10356\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1\
        );

    \I__2186\ : IoInMux
    port map (
            O => \N__10351\,
            I => \N__10348\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__10348\,
            I => \N__10344\
        );

    \I__2184\ : CascadeMux
    port map (
            O => \N__10347\,
            I => \N__10337\
        );

    \I__2183\ : Span4Mux_s2_v
    port map (
            O => \N__10344\,
            I => \N__10330\
        );

    \I__2182\ : InMux
    port map (
            O => \N__10343\,
            I => \N__10323\
        );

    \I__2181\ : InMux
    port map (
            O => \N__10342\,
            I => \N__10323\
        );

    \I__2180\ : InMux
    port map (
            O => \N__10341\,
            I => \N__10323\
        );

    \I__2179\ : InMux
    port map (
            O => \N__10340\,
            I => \N__10316\
        );

    \I__2178\ : InMux
    port map (
            O => \N__10337\,
            I => \N__10316\
        );

    \I__2177\ : InMux
    port map (
            O => \N__10336\,
            I => \N__10309\
        );

    \I__2176\ : InMux
    port map (
            O => \N__10335\,
            I => \N__10309\
        );

    \I__2175\ : InMux
    port map (
            O => \N__10334\,
            I => \N__10309\
        );

    \I__2174\ : InMux
    port map (
            O => \N__10333\,
            I => \N__10306\
        );

    \I__2173\ : Sp12to4
    port map (
            O => \N__10330\,
            I => \N__10303\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__10323\,
            I => \N__10298\
        );

    \I__2171\ : InMux
    port map (
            O => \N__10322\,
            I => \N__10295\
        );

    \I__2170\ : InMux
    port map (
            O => \N__10321\,
            I => \N__10292\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__10316\,
            I => \N__10285\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__10309\,
            I => \N__10285\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__10306\,
            I => \N__10285\
        );

    \I__2166\ : Span12Mux_h
    port map (
            O => \N__10303\,
            I => \N__10282\
        );

    \I__2165\ : InMux
    port map (
            O => \N__10302\,
            I => \N__10279\
        );

    \I__2164\ : InMux
    port map (
            O => \N__10301\,
            I => \N__10276\
        );

    \I__2163\ : Span12Mux_h
    port map (
            O => \N__10298\,
            I => \N__10273\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__10295\,
            I => \N__10270\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__10292\,
            I => \N__10265\
        );

    \I__2160\ : Span4Mux_v
    port map (
            O => \N__10285\,
            I => \N__10265\
        );

    \I__2159\ : Odrv12
    port map (
            O => \N__10282\,
            I => \P1A2_c\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__10279\,
            I => \P1A2_c\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__10276\,
            I => \P1A2_c\
        );

    \I__2156\ : Odrv12
    port map (
            O => \N__10273\,
            I => \P1A2_c\
        );

    \I__2155\ : Odrv12
    port map (
            O => \N__10270\,
            I => \P1A2_c\
        );

    \I__2154\ : Odrv4
    port map (
            O => \N__10265\,
            I => \P1A2_c\
        );

    \I__2153\ : CascadeMux
    port map (
            O => \N__10252\,
            I => \N__10248\
        );

    \I__2152\ : InMux
    port map (
            O => \N__10251\,
            I => \N__10245\
        );

    \I__2151\ : InMux
    port map (
            O => \N__10248\,
            I => \N__10242\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__10245\,
            I => \N__10239\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__10242\,
            I => \N__10234\
        );

    \I__2148\ : Span4Mux_v
    port map (
            O => \N__10239\,
            I => \N__10234\
        );

    \I__2147\ : Span4Mux_h
    port map (
            O => \N__10234\,
            I => \N__10230\
        );

    \I__2146\ : InMux
    port map (
            O => \N__10233\,
            I => \N__10227\
        );

    \I__2145\ : Odrv4
    port map (
            O => \N__10230\,
            I => \rFifoCount_RNIHH0D1_0\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__10227\,
            I => \rFifoCount_RNIHH0D1_0\
        );

    \I__2143\ : InMux
    port map (
            O => \N__10222\,
            I => \N__10219\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__10219\,
            I => \N__10214\
        );

    \I__2141\ : InMux
    port map (
            O => \N__10218\,
            I => \N__10211\
        );

    \I__2140\ : InMux
    port map (
            O => \N__10217\,
            I => \N__10208\
        );

    \I__2139\ : Span4Mux_h
    port map (
            O => \N__10214\,
            I => \N__10201\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__10211\,
            I => \N__10201\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__10208\,
            I => \N__10201\
        );

    \I__2136\ : Span4Mux_v
    port map (
            O => \N__10201\,
            I => \N__10198\
        );

    \I__2135\ : Odrv4
    port map (
            O => \N__10198\,
            I => \rTxWriteZ0\
        );

    \I__2134\ : IoInMux
    port map (
            O => \N__10195\,
            I => \N__10192\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__10192\,
            I => \N__10189\
        );

    \I__2132\ : IoSpan4Mux
    port map (
            O => \N__10189\,
            I => \N__10186\
        );

    \I__2131\ : Span4Mux_s3_v
    port map (
            O => \N__10186\,
            I => \N__10183\
        );

    \I__2130\ : Span4Mux_h
    port map (
            O => \N__10183\,
            I => \N__10179\
        );

    \I__2129\ : IoInMux
    port map (
            O => \N__10182\,
            I => \N__10176\
        );

    \I__2128\ : Span4Mux_h
    port map (
            O => \N__10179\,
            I => \N__10172\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__10176\,
            I => \N__10169\
        );

    \I__2126\ : InMux
    port map (
            O => \N__10175\,
            I => \N__10166\
        );

    \I__2125\ : Odrv4
    port map (
            O => \N__10172\,
            I => \P1A3_c\
        );

    \I__2124\ : Odrv12
    port map (
            O => \N__10169\,
            I => \P1A3_c\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__10166\,
            I => \P1A3_c\
        );

    \I__2122\ : InMux
    port map (
            O => \N__10159\,
            I => \N__10155\
        );

    \I__2121\ : InMux
    port map (
            O => \N__10158\,
            I => \N__10152\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__10155\,
            I => \N__10148\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__10152\,
            I => \N__10145\
        );

    \I__2118\ : InMux
    port map (
            O => \N__10151\,
            I => \N__10142\
        );

    \I__2117\ : Span4Mux_h
    port map (
            O => \N__10148\,
            I => \N__10134\
        );

    \I__2116\ : Span4Mux_v
    port map (
            O => \N__10145\,
            I => \N__10134\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__10142\,
            I => \N__10134\
        );

    \I__2114\ : InMux
    port map (
            O => \N__10141\,
            I => \N__10131\
        );

    \I__2113\ : Odrv4
    port map (
            O => \N__10134\,
            I => \rTxByteZ0Z_2\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__10131\,
            I => \rTxByteZ0Z_2\
        );

    \I__2111\ : InMux
    port map (
            O => \N__10126\,
            I => \N__10123\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__10123\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_2\
        );

    \I__2109\ : InMux
    port map (
            O => \N__10120\,
            I => \N__10117\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__10117\,
            I => \N__10113\
        );

    \I__2107\ : InMux
    port map (
            O => \N__10116\,
            I => \N__10109\
        );

    \I__2106\ : Span4Mux_v
    port map (
            O => \N__10113\,
            I => \N__10106\
        );

    \I__2105\ : InMux
    port map (
            O => \N__10112\,
            I => \N__10103\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__10109\,
            I => \N__10095\
        );

    \I__2103\ : Sp12to4
    port map (
            O => \N__10106\,
            I => \N__10095\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__10103\,
            I => \N__10095\
        );

    \I__2101\ : InMux
    port map (
            O => \N__10102\,
            I => \N__10092\
        );

    \I__2100\ : Odrv12
    port map (
            O => \N__10095\,
            I => \rTxByteZ0Z_7\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__10092\,
            I => \rTxByteZ0Z_7\
        );

    \I__2098\ : InMux
    port map (
            O => \N__10087\,
            I => \N__10084\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__10084\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_7\
        );

    \I__2096\ : CEMux
    port map (
            O => \N__10081\,
            I => \N__10075\
        );

    \I__2095\ : CEMux
    port map (
            O => \N__10080\,
            I => \N__10072\
        );

    \I__2094\ : CEMux
    port map (
            O => \N__10079\,
            I => \N__10068\
        );

    \I__2093\ : CEMux
    port map (
            O => \N__10078\,
            I => \N__10065\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__10075\,
            I => \N__10062\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__10072\,
            I => \N__10058\
        );

    \I__2090\ : CEMux
    port map (
            O => \N__10071\,
            I => \N__10055\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__10068\,
            I => \N__10052\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__10065\,
            I => \N__10049\
        );

    \I__2087\ : Span4Mux_v
    port map (
            O => \N__10062\,
            I => \N__10046\
        );

    \I__2086\ : CEMux
    port map (
            O => \N__10061\,
            I => \N__10043\
        );

    \I__2085\ : Span4Mux_v
    port map (
            O => \N__10058\,
            I => \N__10038\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__10055\,
            I => \N__10038\
        );

    \I__2083\ : Span4Mux_v
    port map (
            O => \N__10052\,
            I => \N__10033\
        );

    \I__2082\ : Span4Mux_h
    port map (
            O => \N__10049\,
            I => \N__10033\
        );

    \I__2081\ : Sp12to4
    port map (
            O => \N__10046\,
            I => \N__10028\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__10043\,
            I => \N__10028\
        );

    \I__2079\ : Span4Mux_h
    port map (
            O => \N__10038\,
            I => \N__10024\
        );

    \I__2078\ : Sp12to4
    port map (
            O => \N__10033\,
            I => \N__10019\
        );

    \I__2077\ : Span12Mux_s11_h
    port map (
            O => \N__10028\,
            I => \N__10019\
        );

    \I__2076\ : InMux
    port map (
            O => \N__10027\,
            I => \N__10016\
        );

    \I__2075\ : Odrv4
    port map (
            O => \N__10024\,
            I => \DUT.fifo_tx_inst.rFifoData_awe0\
        );

    \I__2074\ : Odrv12
    port map (
            O => \N__10019\,
            I => \DUT.fifo_tx_inst.rFifoData_awe0\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__10016\,
            I => \DUT.fifo_tx_inst.rFifoData_awe0\
        );

    \I__2072\ : InMux
    port map (
            O => \N__10009\,
            I => \N__10006\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__10006\,
            I => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0\
        );

    \I__2070\ : CascadeMux
    port map (
            O => \N__10003\,
            I => \N__9998\
        );

    \I__2069\ : CascadeMux
    port map (
            O => \N__10002\,
            I => \N__9995\
        );

    \I__2068\ : InMux
    port map (
            O => \N__10001\,
            I => \N__9990\
        );

    \I__2067\ : InMux
    port map (
            O => \N__9998\,
            I => \N__9987\
        );

    \I__2066\ : InMux
    port map (
            O => \N__9995\,
            I => \N__9980\
        );

    \I__2065\ : InMux
    port map (
            O => \N__9994\,
            I => \N__9980\
        );

    \I__2064\ : InMux
    port map (
            O => \N__9993\,
            I => \N__9980\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__9990\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_0\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__9987\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_0\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__9980\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_0\
        );

    \I__2060\ : CascadeMux
    port map (
            O => \N__9973\,
            I => \N__9970\
        );

    \I__2059\ : InMux
    port map (
            O => \N__9970\,
            I => \N__9967\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__9967\,
            I => \DUT.fifo_tx_inst.rFifoCount_RNISSQ21Z0Z_1\
        );

    \I__2057\ : InMux
    port map (
            O => \N__9964\,
            I => \N__9958\
        );

    \I__2056\ : InMux
    port map (
            O => \N__9963\,
            I => \N__9953\
        );

    \I__2055\ : InMux
    port map (
            O => \N__9962\,
            I => \N__9953\
        );

    \I__2054\ : InMux
    port map (
            O => \N__9961\,
            I => \N__9950\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__9958\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_1\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__9953\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_1\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__9950\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_1\
        );

    \I__2050\ : InMux
    port map (
            O => \N__9943\,
            I => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0\
        );

    \I__2049\ : InMux
    port map (
            O => \N__9940\,
            I => \N__9935\
        );

    \I__2048\ : InMux
    port map (
            O => \N__9939\,
            I => \N__9932\
        );

    \I__2047\ : InMux
    port map (
            O => \N__9938\,
            I => \N__9929\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__9935\,
            I => \DUT.fifo_tx_inst.N_83\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__9932\,
            I => \DUT.fifo_tx_inst.N_83\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__9929\,
            I => \DUT.fifo_tx_inst.N_83\
        );

    \I__2043\ : InMux
    port map (
            O => \N__9922\,
            I => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1\
        );

    \I__2042\ : InMux
    port map (
            O => \N__9919\,
            I => \N__9916\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__9916\,
            I => \N__9911\
        );

    \I__2040\ : CascadeMux
    port map (
            O => \N__9915\,
            I => \N__9907\
        );

    \I__2039\ : InMux
    port map (
            O => \N__9914\,
            I => \N__9903\
        );

    \I__2038\ : Span4Mux_h
    port map (
            O => \N__9911\,
            I => \N__9900\
        );

    \I__2037\ : InMux
    port map (
            O => \N__9910\,
            I => \N__9897\
        );

    \I__2036\ : InMux
    port map (
            O => \N__9907\,
            I => \N__9892\
        );

    \I__2035\ : InMux
    port map (
            O => \N__9906\,
            I => \N__9892\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__9903\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_2\
        );

    \I__2033\ : Odrv4
    port map (
            O => \N__9900\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_2\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__9897\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_2\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__9892\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_2\
        );

    \I__2030\ : CascadeMux
    port map (
            O => \N__9883\,
            I => \N__9878\
        );

    \I__2029\ : InMux
    port map (
            O => \N__9882\,
            I => \N__9871\
        );

    \I__2028\ : InMux
    port map (
            O => \N__9881\,
            I => \N__9871\
        );

    \I__2027\ : InMux
    port map (
            O => \N__9878\,
            I => \N__9871\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__9871\,
            I => \N__9866\
        );

    \I__2025\ : InMux
    port map (
            O => \N__9870\,
            I => \N__9863\
        );

    \I__2024\ : CascadeMux
    port map (
            O => \N__9869\,
            I => \N__9857\
        );

    \I__2023\ : Span4Mux_v
    port map (
            O => \N__9866\,
            I => \N__9852\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__9863\,
            I => \N__9849\
        );

    \I__2021\ : InMux
    port map (
            O => \N__9862\,
            I => \N__9844\
        );

    \I__2020\ : InMux
    port map (
            O => \N__9861\,
            I => \N__9844\
        );

    \I__2019\ : InMux
    port map (
            O => \N__9860\,
            I => \N__9839\
        );

    \I__2018\ : InMux
    port map (
            O => \N__9857\,
            I => \N__9839\
        );

    \I__2017\ : CascadeMux
    port map (
            O => \N__9856\,
            I => \N__9836\
        );

    \I__2016\ : InMux
    port map (
            O => \N__9855\,
            I => \N__9833\
        );

    \I__2015\ : Span4Mux_h
    port map (
            O => \N__9852\,
            I => \N__9824\
        );

    \I__2014\ : Span4Mux_s2_v
    port map (
            O => \N__9849\,
            I => \N__9824\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__9844\,
            I => \N__9824\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__9839\,
            I => \N__9824\
        );

    \I__2011\ : InMux
    port map (
            O => \N__9836\,
            I => \N__9821\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__9833\,
            I => \N__9818\
        );

    \I__2009\ : Span4Mux_h
    port map (
            O => \N__9824\,
            I => \N__9813\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__9821\,
            I => \N__9813\
        );

    \I__2007\ : Span12Mux_h
    port map (
            O => \N__9818\,
            I => \N__9810\
        );

    \I__2006\ : IoSpan4Mux
    port map (
            O => \N__9813\,
            I => \N__9807\
        );

    \I__2005\ : Odrv12
    port map (
            O => \N__9810\,
            I => \P1A1_c\
        );

    \I__2004\ : Odrv4
    port map (
            O => \N__9807\,
            I => \P1A1_c\
        );

    \I__2003\ : InMux
    port map (
            O => \N__9802\,
            I => \N__9797\
        );

    \I__2002\ : InMux
    port map (
            O => \N__9801\,
            I => \N__9794\
        );

    \I__2001\ : InMux
    port map (
            O => \N__9800\,
            I => \N__9791\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__9797\,
            I => \DUT.uart_inst0.recv_stateZ0Z_3\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__9794\,
            I => \DUT.uart_inst0.recv_stateZ0Z_3\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__9791\,
            I => \DUT.uart_inst0.recv_stateZ0Z_3\
        );

    \I__1997\ : InMux
    port map (
            O => \N__9784\,
            I => \N__9781\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__9781\,
            I => \N__9778\
        );

    \I__1995\ : Span4Mux_h
    port map (
            O => \N__9778\,
            I => \N__9775\
        );

    \I__1994\ : Odrv4
    port map (
            O => \N__9775\,
            I => \DUT.uart_inst0.g0_1\
        );

    \I__1993\ : InMux
    port map (
            O => \N__9772\,
            I => \N__9765\
        );

    \I__1992\ : InMux
    port map (
            O => \N__9771\,
            I => \N__9765\
        );

    \I__1991\ : InMux
    port map (
            O => \N__9770\,
            I => \N__9762\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__9765\,
            I => \N__9756\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__9762\,
            I => \N__9753\
        );

    \I__1988\ : InMux
    port map (
            O => \N__9761\,
            I => \N__9748\
        );

    \I__1987\ : InMux
    port map (
            O => \N__9760\,
            I => \N__9748\
        );

    \I__1986\ : InMux
    port map (
            O => \N__9759\,
            I => \N__9743\
        );

    \I__1985\ : Span4Mux_s2_v
    port map (
            O => \N__9756\,
            I => \N__9738\
        );

    \I__1984\ : Span4Mux_h
    port map (
            O => \N__9753\,
            I => \N__9738\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__9748\,
            I => \N__9735\
        );

    \I__1982\ : InMux
    port map (
            O => \N__9747\,
            I => \N__9730\
        );

    \I__1981\ : InMux
    port map (
            O => \N__9746\,
            I => \N__9730\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__9743\,
            I => \DUT.uart_inst0.recv_stateZ0Z_5\
        );

    \I__1979\ : Odrv4
    port map (
            O => \N__9738\,
            I => \DUT.uart_inst0.recv_stateZ0Z_5\
        );

    \I__1978\ : Odrv4
    port map (
            O => \N__9735\,
            I => \DUT.uart_inst0.recv_stateZ0Z_5\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__9730\,
            I => \DUT.uart_inst0.recv_stateZ0Z_5\
        );

    \I__1976\ : InMux
    port map (
            O => \N__9721\,
            I => \N__9717\
        );

    \I__1975\ : CascadeMux
    port map (
            O => \N__9720\,
            I => \N__9708\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__9717\,
            I => \N__9702\
        );

    \I__1973\ : InMux
    port map (
            O => \N__9716\,
            I => \N__9697\
        );

    \I__1972\ : InMux
    port map (
            O => \N__9715\,
            I => \N__9697\
        );

    \I__1971\ : InMux
    port map (
            O => \N__9714\,
            I => \N__9694\
        );

    \I__1970\ : InMux
    port map (
            O => \N__9713\,
            I => \N__9689\
        );

    \I__1969\ : InMux
    port map (
            O => \N__9712\,
            I => \N__9689\
        );

    \I__1968\ : InMux
    port map (
            O => \N__9711\,
            I => \N__9682\
        );

    \I__1967\ : InMux
    port map (
            O => \N__9708\,
            I => \N__9682\
        );

    \I__1966\ : InMux
    port map (
            O => \N__9707\,
            I => \N__9682\
        );

    \I__1965\ : InMux
    port map (
            O => \N__9706\,
            I => \N__9677\
        );

    \I__1964\ : InMux
    port map (
            O => \N__9705\,
            I => \N__9677\
        );

    \I__1963\ : Odrv4
    port map (
            O => \N__9702\,
            I => \DUT.uart_inst0.rx_countdown_3_4\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__9697\,
            I => \DUT.uart_inst0.rx_countdown_3_4\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__9694\,
            I => \DUT.uart_inst0.rx_countdown_3_4\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__9689\,
            I => \DUT.uart_inst0.rx_countdown_3_4\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__9682\,
            I => \DUT.uart_inst0.rx_countdown_3_4\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__9677\,
            I => \DUT.uart_inst0.rx_countdown_3_4\
        );

    \I__1957\ : CascadeMux
    port map (
            O => \N__9664\,
            I => \N__9661\
        );

    \I__1956\ : InMux
    port map (
            O => \N__9661\,
            I => \N__9658\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__9658\,
            I => \N__9655\
        );

    \I__1954\ : Odrv4
    port map (
            O => \N__9655\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_4\
        );

    \I__1953\ : InMux
    port map (
            O => \N__9652\,
            I => \N__9647\
        );

    \I__1952\ : InMux
    port map (
            O => \N__9651\,
            I => \N__9644\
        );

    \I__1951\ : InMux
    port map (
            O => \N__9650\,
            I => \N__9641\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__9647\,
            I => \N__9634\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__9644\,
            I => \N__9634\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__9641\,
            I => \N__9631\
        );

    \I__1947\ : InMux
    port map (
            O => \N__9640\,
            I => \N__9620\
        );

    \I__1946\ : InMux
    port map (
            O => \N__9639\,
            I => \N__9620\
        );

    \I__1945\ : Span4Mux_s2_v
    port map (
            O => \N__9634\,
            I => \N__9617\
        );

    \I__1944\ : Span4Mux_v
    port map (
            O => \N__9631\,
            I => \N__9614\
        );

    \I__1943\ : InMux
    port map (
            O => \N__9630\,
            I => \N__9607\
        );

    \I__1942\ : InMux
    port map (
            O => \N__9629\,
            I => \N__9607\
        );

    \I__1941\ : InMux
    port map (
            O => \N__9628\,
            I => \N__9607\
        );

    \I__1940\ : InMux
    port map (
            O => \N__9627\,
            I => \N__9602\
        );

    \I__1939\ : InMux
    port map (
            O => \N__9626\,
            I => \N__9602\
        );

    \I__1938\ : InMux
    port map (
            O => \N__9625\,
            I => \N__9599\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__9620\,
            I => \DUT.uart_inst0.rx_countdown_3_5\
        );

    \I__1936\ : Odrv4
    port map (
            O => \N__9617\,
            I => \DUT.uart_inst0.rx_countdown_3_5\
        );

    \I__1935\ : Odrv4
    port map (
            O => \N__9614\,
            I => \DUT.uart_inst0.rx_countdown_3_5\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__9607\,
            I => \DUT.uart_inst0.rx_countdown_3_5\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__9602\,
            I => \DUT.uart_inst0.rx_countdown_3_5\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__9599\,
            I => \DUT.uart_inst0.rx_countdown_3_5\
        );

    \I__1931\ : InMux
    port map (
            O => \N__9586\,
            I => \N__9583\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__9583\,
            I => \N__9580\
        );

    \I__1929\ : Odrv4
    port map (
            O => \N__9580\,
            I => \DUT.uart_inst0.recv_state_RNO_2Z0Z_1\
        );

    \I__1928\ : InMux
    port map (
            O => \N__9577\,
            I => \N__9572\
        );

    \I__1927\ : InMux
    port map (
            O => \N__9576\,
            I => \N__9568\
        );

    \I__1926\ : InMux
    port map (
            O => \N__9575\,
            I => \N__9565\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__9572\,
            I => \N__9562\
        );

    \I__1924\ : CascadeMux
    port map (
            O => \N__9571\,
            I => \N__9553\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__9568\,
            I => \N__9548\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__9565\,
            I => \N__9543\
        );

    \I__1921\ : Span4Mux_h
    port map (
            O => \N__9562\,
            I => \N__9543\
        );

    \I__1920\ : InMux
    port map (
            O => \N__9561\,
            I => \N__9536\
        );

    \I__1919\ : InMux
    port map (
            O => \N__9560\,
            I => \N__9536\
        );

    \I__1918\ : InMux
    port map (
            O => \N__9559\,
            I => \N__9536\
        );

    \I__1917\ : InMux
    port map (
            O => \N__9558\,
            I => \N__9531\
        );

    \I__1916\ : InMux
    port map (
            O => \N__9557\,
            I => \N__9531\
        );

    \I__1915\ : InMux
    port map (
            O => \N__9556\,
            I => \N__9526\
        );

    \I__1914\ : InMux
    port map (
            O => \N__9553\,
            I => \N__9526\
        );

    \I__1913\ : InMux
    port map (
            O => \N__9552\,
            I => \N__9523\
        );

    \I__1912\ : InMux
    port map (
            O => \N__9551\,
            I => \N__9520\
        );

    \I__1911\ : Odrv4
    port map (
            O => \N__9548\,
            I => \DUT.uart_inst0.rx_countdown_3_0\
        );

    \I__1910\ : Odrv4
    port map (
            O => \N__9543\,
            I => \DUT.uart_inst0.rx_countdown_3_0\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__9536\,
            I => \DUT.uart_inst0.rx_countdown_3_0\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__9531\,
            I => \DUT.uart_inst0.rx_countdown_3_0\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__9526\,
            I => \DUT.uart_inst0.rx_countdown_3_0\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__9523\,
            I => \DUT.uart_inst0.rx_countdown_3_0\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__9520\,
            I => \DUT.uart_inst0.rx_countdown_3_0\
        );

    \I__1904\ : InMux
    port map (
            O => \N__9505\,
            I => \N__9500\
        );

    \I__1903\ : CascadeMux
    port map (
            O => \N__9504\,
            I => \N__9494\
        );

    \I__1902\ : CascadeMux
    port map (
            O => \N__9503\,
            I => \N__9491\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__9500\,
            I => \N__9488\
        );

    \I__1900\ : CascadeMux
    port map (
            O => \N__9499\,
            I => \N__9483\
        );

    \I__1899\ : CascadeMux
    port map (
            O => \N__9498\,
            I => \N__9480\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__9497\,
            I => \N__9476\
        );

    \I__1897\ : InMux
    port map (
            O => \N__9494\,
            I => \N__9471\
        );

    \I__1896\ : InMux
    port map (
            O => \N__9491\,
            I => \N__9471\
        );

    \I__1895\ : Span4Mux_h
    port map (
            O => \N__9488\,
            I => \N__9468\
        );

    \I__1894\ : InMux
    port map (
            O => \N__9487\,
            I => \N__9465\
        );

    \I__1893\ : InMux
    port map (
            O => \N__9486\,
            I => \N__9462\
        );

    \I__1892\ : InMux
    port map (
            O => \N__9483\,
            I => \N__9459\
        );

    \I__1891\ : InMux
    port map (
            O => \N__9480\,
            I => \N__9452\
        );

    \I__1890\ : InMux
    port map (
            O => \N__9479\,
            I => \N__9452\
        );

    \I__1889\ : InMux
    port map (
            O => \N__9476\,
            I => \N__9452\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__9471\,
            I => \DUT.uart_inst0.rx_countdown_3_2\
        );

    \I__1887\ : Odrv4
    port map (
            O => \N__9468\,
            I => \DUT.uart_inst0.rx_countdown_3_2\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__9465\,
            I => \DUT.uart_inst0.rx_countdown_3_2\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__9462\,
            I => \DUT.uart_inst0.rx_countdown_3_2\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__9459\,
            I => \DUT.uart_inst0.rx_countdown_3_2\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__9452\,
            I => \DUT.uart_inst0.rx_countdown_3_2\
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__9439\,
            I => \DUT.uart_inst0.G_10_i_a4_0_4_cascade_\
        );

    \I__1881\ : InMux
    port map (
            O => \N__9436\,
            I => \N__9432\
        );

    \I__1880\ : InMux
    port map (
            O => \N__9435\,
            I => \N__9425\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__9432\,
            I => \N__9422\
        );

    \I__1878\ : CascadeMux
    port map (
            O => \N__9431\,
            I => \N__9413\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__9430\,
            I => \N__9410\
        );

    \I__1876\ : InMux
    port map (
            O => \N__9429\,
            I => \N__9405\
        );

    \I__1875\ : InMux
    port map (
            O => \N__9428\,
            I => \N__9405\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__9425\,
            I => \N__9400\
        );

    \I__1873\ : Span4Mux_h
    port map (
            O => \N__9422\,
            I => \N__9400\
        );

    \I__1872\ : InMux
    port map (
            O => \N__9421\,
            I => \N__9397\
        );

    \I__1871\ : InMux
    port map (
            O => \N__9420\,
            I => \N__9388\
        );

    \I__1870\ : InMux
    port map (
            O => \N__9419\,
            I => \N__9388\
        );

    \I__1869\ : InMux
    port map (
            O => \N__9418\,
            I => \N__9388\
        );

    \I__1868\ : InMux
    port map (
            O => \N__9417\,
            I => \N__9388\
        );

    \I__1867\ : InMux
    port map (
            O => \N__9416\,
            I => \N__9385\
        );

    \I__1866\ : InMux
    port map (
            O => \N__9413\,
            I => \N__9380\
        );

    \I__1865\ : InMux
    port map (
            O => \N__9410\,
            I => \N__9380\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__9405\,
            I => \DUT.uart_inst0.rx_countdown_3_3\
        );

    \I__1863\ : Odrv4
    port map (
            O => \N__9400\,
            I => \DUT.uart_inst0.rx_countdown_3_3\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__9397\,
            I => \DUT.uart_inst0.rx_countdown_3_3\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__9388\,
            I => \DUT.uart_inst0.rx_countdown_3_3\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__9385\,
            I => \DUT.uart_inst0.rx_countdown_3_3\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__9380\,
            I => \DUT.uart_inst0.rx_countdown_3_3\
        );

    \I__1858\ : CascadeMux
    port map (
            O => \N__9367\,
            I => \DUT.uart_inst0.N_4_i_0_1_cascade_\
        );

    \I__1857\ : InMux
    port map (
            O => \N__9364\,
            I => \N__9355\
        );

    \I__1856\ : InMux
    port map (
            O => \N__9363\,
            I => \N__9355\
        );

    \I__1855\ : InMux
    port map (
            O => \N__9362\,
            I => \N__9355\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__9355\,
            I => \N__9343\
        );

    \I__1853\ : InMux
    port map (
            O => \N__9354\,
            I => \N__9332\
        );

    \I__1852\ : InMux
    port map (
            O => \N__9353\,
            I => \N__9332\
        );

    \I__1851\ : InMux
    port map (
            O => \N__9352\,
            I => \N__9332\
        );

    \I__1850\ : InMux
    port map (
            O => \N__9351\,
            I => \N__9332\
        );

    \I__1849\ : InMux
    port map (
            O => \N__9350\,
            I => \N__9332\
        );

    \I__1848\ : InMux
    port map (
            O => \N__9349\,
            I => \N__9327\
        );

    \I__1847\ : InMux
    port map (
            O => \N__9348\,
            I => \N__9327\
        );

    \I__1846\ : CascadeMux
    port map (
            O => \N__9347\,
            I => \N__9324\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__9346\,
            I => \N__9321\
        );

    \I__1844\ : Span4Mux_s2_v
    port map (
            O => \N__9343\,
            I => \N__9305\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__9332\,
            I => \N__9300\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__9327\,
            I => \N__9300\
        );

    \I__1841\ : InMux
    port map (
            O => \N__9324\,
            I => \N__9287\
        );

    \I__1840\ : InMux
    port map (
            O => \N__9321\,
            I => \N__9287\
        );

    \I__1839\ : InMux
    port map (
            O => \N__9320\,
            I => \N__9287\
        );

    \I__1838\ : InMux
    port map (
            O => \N__9319\,
            I => \N__9287\
        );

    \I__1837\ : InMux
    port map (
            O => \N__9318\,
            I => \N__9287\
        );

    \I__1836\ : InMux
    port map (
            O => \N__9317\,
            I => \N__9287\
        );

    \I__1835\ : InMux
    port map (
            O => \N__9316\,
            I => \N__9284\
        );

    \I__1834\ : InMux
    port map (
            O => \N__9315\,
            I => \N__9281\
        );

    \I__1833\ : InMux
    port map (
            O => \N__9314\,
            I => \N__9278\
        );

    \I__1832\ : InMux
    port map (
            O => \N__9313\,
            I => \N__9271\
        );

    \I__1831\ : InMux
    port map (
            O => \N__9312\,
            I => \N__9271\
        );

    \I__1830\ : InMux
    port map (
            O => \N__9311\,
            I => \N__9271\
        );

    \I__1829\ : InMux
    port map (
            O => \N__9310\,
            I => \N__9264\
        );

    \I__1828\ : InMux
    port map (
            O => \N__9309\,
            I => \N__9264\
        );

    \I__1827\ : InMux
    port map (
            O => \N__9308\,
            I => \N__9264\
        );

    \I__1826\ : Span4Mux_h
    port map (
            O => \N__9305\,
            I => \N__9259\
        );

    \I__1825\ : Span4Mux_s2_v
    port map (
            O => \N__9300\,
            I => \N__9259\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__9287\,
            I => \N__9254\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__9284\,
            I => \N__9254\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__9281\,
            I => \DUT.uart_inst0.N_149\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__9278\,
            I => \DUT.uart_inst0.N_149\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__9271\,
            I => \DUT.uart_inst0.N_149\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__9264\,
            I => \DUT.uart_inst0.N_149\
        );

    \I__1818\ : Odrv4
    port map (
            O => \N__9259\,
            I => \DUT.uart_inst0.N_149\
        );

    \I__1817\ : Odrv4
    port map (
            O => \N__9254\,
            I => \DUT.uart_inst0.N_149\
        );

    \I__1816\ : InMux
    port map (
            O => \N__9241\,
            I => \N__9238\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__9238\,
            I => \N__9231\
        );

    \I__1814\ : InMux
    port map (
            O => \N__9237\,
            I => \N__9224\
        );

    \I__1813\ : InMux
    port map (
            O => \N__9236\,
            I => \N__9224\
        );

    \I__1812\ : InMux
    port map (
            O => \N__9235\,
            I => \N__9224\
        );

    \I__1811\ : InMux
    port map (
            O => \N__9234\,
            I => \N__9216\
        );

    \I__1810\ : Span4Mux_h
    port map (
            O => \N__9231\,
            I => \N__9213\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__9224\,
            I => \N__9210\
        );

    \I__1808\ : InMux
    port map (
            O => \N__9223\,
            I => \N__9205\
        );

    \I__1807\ : InMux
    port map (
            O => \N__9222\,
            I => \N__9205\
        );

    \I__1806\ : InMux
    port map (
            O => \N__9221\,
            I => \N__9198\
        );

    \I__1805\ : InMux
    port map (
            O => \N__9220\,
            I => \N__9198\
        );

    \I__1804\ : InMux
    port map (
            O => \N__9219\,
            I => \N__9198\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__9216\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__1802\ : Odrv4
    port map (
            O => \N__9213\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__1801\ : Odrv4
    port map (
            O => \N__9210\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__9205\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__9198\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__1798\ : InMux
    port map (
            O => \N__9187\,
            I => \N__9184\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__9184\,
            I => \DUT.rFifoDatarx_4\
        );

    \I__1796\ : CascadeMux
    port map (
            O => \N__9181\,
            I => \N__9178\
        );

    \I__1795\ : InMux
    port map (
            O => \N__9178\,
            I => \N__9175\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__9175\,
            I => \DUT.uart_inst0.tx_dataZ0Z_5\
        );

    \I__1793\ : CascadeMux
    port map (
            O => \N__9172\,
            I => \N__9169\
        );

    \I__1792\ : InMux
    port map (
            O => \N__9169\,
            I => \N__9166\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__9166\,
            I => \N__9163\
        );

    \I__1790\ : Odrv12
    port map (
            O => \N__9163\,
            I => \DUT.uart_inst0.tx_dataZ0Z_4\
        );

    \I__1789\ : InMux
    port map (
            O => \N__9160\,
            I => \N__9157\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__9157\,
            I => \DUT.rFifoDatarx_7\
        );

    \I__1787\ : CascadeMux
    port map (
            O => \N__9154\,
            I => \N__9150\
        );

    \I__1786\ : InMux
    port map (
            O => \N__9153\,
            I => \N__9139\
        );

    \I__1785\ : InMux
    port map (
            O => \N__9150\,
            I => \N__9139\
        );

    \I__1784\ : InMux
    port map (
            O => \N__9149\,
            I => \N__9139\
        );

    \I__1783\ : InMux
    port map (
            O => \N__9148\,
            I => \N__9139\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__9139\,
            I => \N__9132\
        );

    \I__1781\ : InMux
    port map (
            O => \N__9138\,
            I => \N__9123\
        );

    \I__1780\ : InMux
    port map (
            O => \N__9137\,
            I => \N__9123\
        );

    \I__1779\ : InMux
    port map (
            O => \N__9136\,
            I => \N__9123\
        );

    \I__1778\ : InMux
    port map (
            O => \N__9135\,
            I => \N__9123\
        );

    \I__1777\ : Odrv4
    port map (
            O => \N__9132\,
            I => \DUT.uart_inst0.N_145\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__9123\,
            I => \DUT.uart_inst0.N_145\
        );

    \I__1775\ : CascadeMux
    port map (
            O => \N__9118\,
            I => \N__9115\
        );

    \I__1774\ : InMux
    port map (
            O => \N__9115\,
            I => \N__9112\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__9112\,
            I => \DUT.uart_inst0.tx_dataZ0Z_7\
        );

    \I__1772\ : CEMux
    port map (
            O => \N__9109\,
            I => \N__9106\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__9106\,
            I => \N__9103\
        );

    \I__1770\ : Span4Mux_v
    port map (
            O => \N__9103\,
            I => \N__9099\
        );

    \I__1769\ : CEMux
    port map (
            O => \N__9102\,
            I => \N__9096\
        );

    \I__1768\ : Span4Mux_h
    port map (
            O => \N__9099\,
            I => \N__9093\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__9096\,
            I => \N__9090\
        );

    \I__1766\ : Odrv4
    port map (
            O => \N__9093\,
            I => \DUT.uart_inst0.N_22_i\
        );

    \I__1765\ : Odrv12
    port map (
            O => \N__9090\,
            I => \DUT.uart_inst0.N_22_i\
        );

    \I__1764\ : CascadeMux
    port map (
            O => \N__9085\,
            I => \DUT.fifo_tx_inst.N_83_cascade_\
        );

    \I__1763\ : InMux
    port map (
            O => \N__9082\,
            I => \N__9078\
        );

    \I__1762\ : CascadeMux
    port map (
            O => \N__9081\,
            I => \N__9075\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__9078\,
            I => \N__9072\
        );

    \I__1760\ : InMux
    port map (
            O => \N__9075\,
            I => \N__9069\
        );

    \I__1759\ : Odrv12
    port map (
            O => \N__9072\,
            I => \DUT.uart_inst0.tx_dataZ0Z_0\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__9069\,
            I => \DUT.uart_inst0.tx_dataZ0Z_0\
        );

    \I__1757\ : CascadeMux
    port map (
            O => \N__9064\,
            I => \N__9061\
        );

    \I__1756\ : InMux
    port map (
            O => \N__9061\,
            I => \N__9057\
        );

    \I__1755\ : IoInMux
    port map (
            O => \N__9060\,
            I => \N__9054\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__9057\,
            I => \N__9050\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__9054\,
            I => \N__9047\
        );

    \I__1752\ : InMux
    port map (
            O => \N__9053\,
            I => \N__9043\
        );

    \I__1751\ : Span4Mux_h
    port map (
            O => \N__9050\,
            I => \N__9040\
        );

    \I__1750\ : Span4Mux_s0_v
    port map (
            O => \N__9047\,
            I => \N__9037\
        );

    \I__1749\ : CascadeMux
    port map (
            O => \N__9046\,
            I => \N__9034\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__9043\,
            I => \N__9031\
        );

    \I__1747\ : Span4Mux_v
    port map (
            O => \N__9040\,
            I => \N__9028\
        );

    \I__1746\ : Span4Mux_h
    port map (
            O => \N__9037\,
            I => \N__9025\
        );

    \I__1745\ : InMux
    port map (
            O => \N__9034\,
            I => \N__9022\
        );

    \I__1744\ : Span12Mux_s11_h
    port map (
            O => \N__9031\,
            I => \N__9019\
        );

    \I__1743\ : Span4Mux_v
    port map (
            O => \N__9028\,
            I => \N__9016\
        );

    \I__1742\ : Odrv4
    port map (
            O => \N__9025\,
            I => \P1A7_c\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__9022\,
            I => \P1A7_c\
        );

    \I__1740\ : Odrv12
    port map (
            O => \N__9019\,
            I => \P1A7_c\
        );

    \I__1739\ : Odrv4
    port map (
            O => \N__9016\,
            I => \P1A7_c\
        );

    \I__1738\ : CascadeMux
    port map (
            O => \N__9007\,
            I => \N__9004\
        );

    \I__1737\ : InMux
    port map (
            O => \N__9004\,
            I => \N__9001\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__9001\,
            I => \N__8998\
        );

    \I__1735\ : Odrv4
    port map (
            O => \N__8998\,
            I => \DUT.uart_inst0.N_98\
        );

    \I__1734\ : InMux
    port map (
            O => \N__8995\,
            I => \N__8992\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__8992\,
            I => \fifo_inst.ftdi_output_inst.rFifoStatec_0\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__8989\,
            I => \N__8986\
        );

    \I__1731\ : InMux
    port map (
            O => \N__8986\,
            I => \N__8978\
        );

    \I__1730\ : InMux
    port map (
            O => \N__8985\,
            I => \N__8969\
        );

    \I__1729\ : InMux
    port map (
            O => \N__8984\,
            I => \N__8969\
        );

    \I__1728\ : InMux
    port map (
            O => \N__8983\,
            I => \N__8969\
        );

    \I__1727\ : InMux
    port map (
            O => \N__8982\,
            I => \N__8969\
        );

    \I__1726\ : InMux
    port map (
            O => \N__8981\,
            I => \N__8966\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__8978\,
            I => \DUT.fifo_tx_inst.N_79\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__8969\,
            I => \DUT.fifo_tx_inst.N_79\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__8966\,
            I => \DUT.fifo_tx_inst.N_79\
        );

    \I__1722\ : InMux
    port map (
            O => \N__8959\,
            I => \N__8956\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__8956\,
            I => \DUT.uart_inst0.tx_dataZ0Z_2\
        );

    \I__1720\ : InMux
    port map (
            O => \N__8953\,
            I => \N__8950\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__8950\,
            I => \DUT.rFifoDatarx_0_3\
        );

    \I__1718\ : InMux
    port map (
            O => \N__8947\,
            I => \N__8944\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__8944\,
            I => \N__8941\
        );

    \I__1716\ : Odrv4
    port map (
            O => \N__8941\,
            I => \DUT.uart_inst0.tx_dataZ0Z_3\
        );

    \I__1715\ : InMux
    port map (
            O => \N__8938\,
            I => \N__8935\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__8935\,
            I => \N__8932\
        );

    \I__1713\ : Span4Mux_h
    port map (
            O => \N__8932\,
            I => \N__8929\
        );

    \I__1712\ : Odrv4
    port map (
            O => \N__8929\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_7\
        );

    \I__1711\ : InMux
    port map (
            O => \N__8926\,
            I => \N__8923\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__8923\,
            I => \N__8920\
        );

    \I__1709\ : Odrv4
    port map (
            O => \N__8920\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_7\
        );

    \I__1708\ : CascadeMux
    port map (
            O => \N__8917\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_\
        );

    \I__1707\ : InMux
    port map (
            O => \N__8914\,
            I => \N__8911\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__8911\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_7\
        );

    \I__1705\ : InMux
    port map (
            O => \N__8908\,
            I => \N__8905\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__8905\,
            I => \DUT.uart_inst0.tx_out_6_iv_0_a3_0_1\
        );

    \I__1703\ : InMux
    port map (
            O => \N__8902\,
            I => \N__8899\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__8899\,
            I => \DUT.uart_inst0.N_101\
        );

    \I__1701\ : InMux
    port map (
            O => \N__8896\,
            I => \N__8893\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8893\,
            I => \DUT.rFifoDatarx_5\
        );

    \I__1699\ : InMux
    port map (
            O => \N__8890\,
            I => \N__8887\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__8887\,
            I => \DUT.rFifoDatarx_0_6\
        );

    \I__1697\ : CascadeMux
    port map (
            O => \N__8884\,
            I => \N__8881\
        );

    \I__1696\ : InMux
    port map (
            O => \N__8881\,
            I => \N__8878\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__8878\,
            I => \DUT.uart_inst0.tx_dataZ0Z_6\
        );

    \I__1694\ : InMux
    port map (
            O => \N__8875\,
            I => \N__8872\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__8872\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_2\
        );

    \I__1692\ : CascadeMux
    port map (
            O => \N__8869\,
            I => \N__8866\
        );

    \I__1691\ : InMux
    port map (
            O => \N__8866\,
            I => \N__8863\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__8863\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_2\
        );

    \I__1689\ : InMux
    port map (
            O => \N__8860\,
            I => \N__8857\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__8857\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_1\
        );

    \I__1687\ : CascadeMux
    port map (
            O => \N__8854\,
            I => \N__8851\
        );

    \I__1686\ : InMux
    port map (
            O => \N__8851\,
            I => \N__8848\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__8848\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_1\
        );

    \I__1684\ : InMux
    port map (
            O => \N__8845\,
            I => \N__8842\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__8842\,
            I => \N__8839\
        );

    \I__1682\ : Odrv4
    port map (
            O => \N__8839\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1\
        );

    \I__1681\ : InMux
    port map (
            O => \N__8836\,
            I => \N__8833\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__8833\,
            I => \N__8830\
        );

    \I__1679\ : Span4Mux_h
    port map (
            O => \N__8830\,
            I => \N__8827\
        );

    \I__1678\ : Odrv4
    port map (
            O => \N__8827\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_2\
        );

    \I__1677\ : InMux
    port map (
            O => \N__8824\,
            I => \N__8821\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__8821\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2\
        );

    \I__1675\ : InMux
    port map (
            O => \N__8818\,
            I => \N__8815\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__8815\,
            I => \N__8812\
        );

    \I__1673\ : Span4Mux_h
    port map (
            O => \N__8812\,
            I => \N__8809\
        );

    \I__1672\ : Odrv4
    port map (
            O => \N__8809\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_3\
        );

    \I__1671\ : CascadeMux
    port map (
            O => \N__8806\,
            I => \N__8803\
        );

    \I__1670\ : InMux
    port map (
            O => \N__8803\,
            I => \N__8800\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__8800\,
            I => \N__8797\
        );

    \I__1668\ : Span4Mux_v
    port map (
            O => \N__8797\,
            I => \N__8794\
        );

    \I__1667\ : Odrv4
    port map (
            O => \N__8794\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_3\
        );

    \I__1666\ : InMux
    port map (
            O => \N__8791\,
            I => \N__8788\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__8788\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_3\
        );

    \I__1664\ : CascadeMux
    port map (
            O => \N__8785\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_\
        );

    \I__1663\ : InMux
    port map (
            O => \N__8782\,
            I => \N__8779\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__8779\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_3\
        );

    \I__1661\ : InMux
    port map (
            O => \N__8776\,
            I => \N__8773\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__8773\,
            I => \N__8770\
        );

    \I__1659\ : Span4Mux_h
    port map (
            O => \N__8770\,
            I => \N__8767\
        );

    \I__1658\ : Odrv4
    port map (
            O => \N__8767\,
            I => \DUT.rFifoDatarx_0_0\
        );

    \I__1657\ : InMux
    port map (
            O => \N__8764\,
            I => \N__8761\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__8761\,
            I => \N__8758\
        );

    \I__1655\ : Span4Mux_s2_v
    port map (
            O => \N__8758\,
            I => \N__8755\
        );

    \I__1654\ : Span4Mux_v
    port map (
            O => \N__8755\,
            I => \N__8752\
        );

    \I__1653\ : Odrv4
    port map (
            O => \N__8752\,
            I => \DUT.uart_inst0.tx_out_6_iv_0_1\
        );

    \I__1652\ : InMux
    port map (
            O => \N__8749\,
            I => \N__8746\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__8746\,
            I => \DUT.rFifoDatarx_1\
        );

    \I__1650\ : CascadeMux
    port map (
            O => \N__8743\,
            I => \N__8740\
        );

    \I__1649\ : InMux
    port map (
            O => \N__8740\,
            I => \N__8737\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__8737\,
            I => \DUT.uart_inst0.tx_dataZ0Z_1\
        );

    \I__1647\ : InMux
    port map (
            O => \N__8734\,
            I => \N__8731\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__8731\,
            I => \DUT.rFifoDatarx_2\
        );

    \I__1645\ : InMux
    port map (
            O => \N__8728\,
            I => \N__8725\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__8725\,
            I => \N__8722\
        );

    \I__1643\ : Odrv4
    port map (
            O => \N__8722\,
            I => \DUT.uart_inst0.N_31_0\
        );

    \I__1642\ : InMux
    port map (
            O => \N__8719\,
            I => \N__8716\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__8716\,
            I => \DUT.uart_inst0.N_203\
        );

    \I__1640\ : InMux
    port map (
            O => \N__8713\,
            I => \N__8710\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__8710\,
            I => \DUT.uart_inst0.recv_state_ns_0_i_0_0_a3_0_0_3\
        );

    \I__1638\ : InMux
    port map (
            O => \N__8707\,
            I => \N__8703\
        );

    \I__1637\ : InMux
    port map (
            O => \N__8706\,
            I => \N__8698\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__8703\,
            I => \N__8695\
        );

    \I__1635\ : InMux
    port map (
            O => \N__8702\,
            I => \N__8692\
        );

    \I__1634\ : InMux
    port map (
            O => \N__8701\,
            I => \N__8689\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__8698\,
            I => \N__8686\
        );

    \I__1632\ : Span4Mux_h
    port map (
            O => \N__8695\,
            I => \N__8683\
        );

    \I__1631\ : LocalMux
    port map (
            O => \N__8692\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_2\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__8689\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_2\
        );

    \I__1629\ : Odrv4
    port map (
            O => \N__8686\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_2\
        );

    \I__1628\ : Odrv4
    port map (
            O => \N__8683\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_2\
        );

    \I__1627\ : InMux
    port map (
            O => \N__8674\,
            I => \N__8669\
        );

    \I__1626\ : InMux
    port map (
            O => \N__8673\,
            I => \N__8666\
        );

    \I__1625\ : CascadeMux
    port map (
            O => \N__8672\,
            I => \N__8663\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__8669\,
            I => \N__8655\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__8666\,
            I => \N__8655\
        );

    \I__1622\ : InMux
    port map (
            O => \N__8663\,
            I => \N__8652\
        );

    \I__1621\ : InMux
    port map (
            O => \N__8662\,
            I => \N__8645\
        );

    \I__1620\ : InMux
    port map (
            O => \N__8661\,
            I => \N__8645\
        );

    \I__1619\ : InMux
    port map (
            O => \N__8660\,
            I => \N__8645\
        );

    \I__1618\ : Span4Mux_v
    port map (
            O => \N__8655\,
            I => \N__8642\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__8652\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_1\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__8645\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_1\
        );

    \I__1615\ : Odrv4
    port map (
            O => \N__8642\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_1\
        );

    \I__1614\ : CascadeMux
    port map (
            O => \N__8635\,
            I => \N__8632\
        );

    \I__1613\ : InMux
    port map (
            O => \N__8632\,
            I => \N__8628\
        );

    \I__1612\ : InMux
    port map (
            O => \N__8631\,
            I => \N__8625\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__8628\,
            I => \N__8622\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__8625\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_3\
        );

    \I__1609\ : Odrv4
    port map (
            O => \N__8622\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_3\
        );

    \I__1608\ : CascadeMux
    port map (
            O => \N__8617\,
            I => \N__8614\
        );

    \I__1607\ : InMux
    port map (
            O => \N__8614\,
            I => \N__8610\
        );

    \I__1606\ : CascadeMux
    port map (
            O => \N__8613\,
            I => \N__8606\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__8610\,
            I => \N__8601\
        );

    \I__1604\ : InMux
    port map (
            O => \N__8609\,
            I => \N__8598\
        );

    \I__1603\ : InMux
    port map (
            O => \N__8606\,
            I => \N__8591\
        );

    \I__1602\ : InMux
    port map (
            O => \N__8605\,
            I => \N__8591\
        );

    \I__1601\ : InMux
    port map (
            O => \N__8604\,
            I => \N__8591\
        );

    \I__1600\ : Span4Mux_s3_v
    port map (
            O => \N__8601\,
            I => \N__8586\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__8598\,
            I => \N__8586\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__8591\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_0\
        );

    \I__1597\ : Odrv4
    port map (
            O => \N__8586\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_0\
        );

    \I__1596\ : InMux
    port map (
            O => \N__8581\,
            I => \N__8578\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__8578\,
            I => \DUT.uart_inst0.N_215_4\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__8575\,
            I => \DUT.uart_inst0.N_215_4_cascade_\
        );

    \I__1593\ : CascadeMux
    port map (
            O => \N__8572\,
            I => \DUT.uart_inst0.recv_state_srsts_1_2_cascade_\
        );

    \I__1592\ : InMux
    port map (
            O => \N__8569\,
            I => \N__8565\
        );

    \I__1591\ : InMux
    port map (
            O => \N__8568\,
            I => \N__8562\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__8565\,
            I => \DUT.uart_inst0.N_193\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__8562\,
            I => \DUT.uart_inst0.N_193\
        );

    \I__1588\ : InMux
    port map (
            O => \N__8557\,
            I => \N__8548\
        );

    \I__1587\ : InMux
    port map (
            O => \N__8556\,
            I => \N__8543\
        );

    \I__1586\ : InMux
    port map (
            O => \N__8555\,
            I => \N__8543\
        );

    \I__1585\ : InMux
    port map (
            O => \N__8554\,
            I => \N__8540\
        );

    \I__1584\ : InMux
    port map (
            O => \N__8553\,
            I => \N__8533\
        );

    \I__1583\ : InMux
    port map (
            O => \N__8552\,
            I => \N__8533\
        );

    \I__1582\ : InMux
    port map (
            O => \N__8551\,
            I => \N__8533\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__8548\,
            I => \DUT.uart_inst0.recv_stateZ0Z_2\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__8543\,
            I => \DUT.uart_inst0.recv_stateZ0Z_2\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__8540\,
            I => \DUT.uart_inst0.recv_stateZ0Z_2\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__8533\,
            I => \DUT.uart_inst0.recv_stateZ0Z_2\
        );

    \I__1577\ : InMux
    port map (
            O => \N__8524\,
            I => \N__8521\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__8521\,
            I => \N__8518\
        );

    \I__1575\ : Odrv4
    port map (
            O => \N__8518\,
            I => \DUT.uart_inst0.g0_0\
        );

    \I__1574\ : InMux
    port map (
            O => \N__8515\,
            I => \N__8511\
        );

    \I__1573\ : InMux
    port map (
            O => \N__8514\,
            I => \N__8507\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__8511\,
            I => \N__8503\
        );

    \I__1571\ : InMux
    port map (
            O => \N__8510\,
            I => \N__8500\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__8507\,
            I => \N__8497\
        );

    \I__1569\ : InMux
    port map (
            O => \N__8506\,
            I => \N__8494\
        );

    \I__1568\ : Span4Mux_v
    port map (
            O => \N__8503\,
            I => \N__8491\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__8500\,
            I => \N__8488\
        );

    \I__1566\ : Span4Mux_h
    port map (
            O => \N__8497\,
            I => \N__8483\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__8494\,
            I => \N__8483\
        );

    \I__1564\ : Span4Mux_v
    port map (
            O => \N__8491\,
            I => \N__8479\
        );

    \I__1563\ : Span4Mux_v
    port map (
            O => \N__8488\,
            I => \N__8476\
        );

    \I__1562\ : Span4Mux_v
    port map (
            O => \N__8483\,
            I => \N__8473\
        );

    \I__1561\ : InMux
    port map (
            O => \N__8482\,
            I => \N__8470\
        );

    \I__1560\ : Odrv4
    port map (
            O => \N__8479\,
            I => \DUT.wRxByte_3\
        );

    \I__1559\ : Odrv4
    port map (
            O => \N__8476\,
            I => \DUT.wRxByte_3\
        );

    \I__1558\ : Odrv4
    port map (
            O => \N__8473\,
            I => \DUT.wRxByte_3\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__8470\,
            I => \DUT.wRxByte_3\
        );

    \I__1556\ : InMux
    port map (
            O => \N__8461\,
            I => \N__8456\
        );

    \I__1555\ : InMux
    port map (
            O => \N__8460\,
            I => \N__8453\
        );

    \I__1554\ : InMux
    port map (
            O => \N__8459\,
            I => \N__8450\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__8456\,
            I => \N__8446\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__8453\,
            I => \N__8441\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__8450\,
            I => \N__8441\
        );

    \I__1550\ : InMux
    port map (
            O => \N__8449\,
            I => \N__8438\
        );

    \I__1549\ : Span4Mux_h
    port map (
            O => \N__8446\,
            I => \N__8431\
        );

    \I__1548\ : Span4Mux_v
    port map (
            O => \N__8441\,
            I => \N__8431\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__8438\,
            I => \N__8431\
        );

    \I__1546\ : Span4Mux_v
    port map (
            O => \N__8431\,
            I => \N__8427\
        );

    \I__1545\ : InMux
    port map (
            O => \N__8430\,
            I => \N__8424\
        );

    \I__1544\ : Odrv4
    port map (
            O => \N__8427\,
            I => \DUT.wRxByte_2\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__8424\,
            I => \DUT.wRxByte_2\
        );

    \I__1542\ : CEMux
    port map (
            O => \N__8419\,
            I => \N__8415\
        );

    \I__1541\ : CEMux
    port map (
            O => \N__8418\,
            I => \N__8412\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__8415\,
            I => \N__8409\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__8412\,
            I => \N__8406\
        );

    \I__1538\ : Span4Mux_h
    port map (
            O => \N__8409\,
            I => \N__8403\
        );

    \I__1537\ : Span4Mux_h
    port map (
            O => \N__8406\,
            I => \N__8400\
        );

    \I__1536\ : Odrv4
    port map (
            O => \N__8403\,
            I => \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa\
        );

    \I__1535\ : Odrv4
    port map (
            O => \N__8400\,
            I => \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa\
        );

    \I__1534\ : InMux
    port map (
            O => \N__8395\,
            I => \N__8392\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__8392\,
            I => \DUT.uart_inst0.g0_0_3\
        );

    \I__1532\ : InMux
    port map (
            O => \N__8389\,
            I => \N__8386\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__8386\,
            I => \DUT.uart_inst0.g1\
        );

    \I__1530\ : CascadeMux
    port map (
            O => \N__8383\,
            I => \N__8380\
        );

    \I__1529\ : InMux
    port map (
            O => \N__8380\,
            I => \N__8377\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__8377\,
            I => \DUT.uart_inst0.g0_0_0\
        );

    \I__1527\ : InMux
    port map (
            O => \N__8374\,
            I => \N__8371\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__8371\,
            I => \N__8368\
        );

    \I__1525\ : Span4Mux_v
    port map (
            O => \N__8368\,
            I => \N__8365\
        );

    \I__1524\ : Odrv4
    port map (
            O => \N__8365\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_2\
        );

    \I__1523\ : InMux
    port map (
            O => \N__8362\,
            I => \N__8358\
        );

    \I__1522\ : InMux
    port map (
            O => \N__8361\,
            I => \N__8355\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__8358\,
            I => \DUT.uart_inst0.rx_clk_divider_1_17\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__8355\,
            I => \DUT.uart_inst0.rx_clk_divider_1_17\
        );

    \I__1519\ : InMux
    port map (
            O => \N__8350\,
            I => \N__8347\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__8347\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_17\
        );

    \I__1517\ : InMux
    port map (
            O => \N__8344\,
            I => \N__8340\
        );

    \I__1516\ : InMux
    port map (
            O => \N__8343\,
            I => \N__8337\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__8340\,
            I => \DUT.uart_inst0.rx_clk_divider_1_10\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__8337\,
            I => \DUT.uart_inst0.rx_clk_divider_1_10\
        );

    \I__1513\ : InMux
    port map (
            O => \N__8332\,
            I => \N__8329\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__8329\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_10\
        );

    \I__1511\ : InMux
    port map (
            O => \N__8326\,
            I => \N__8322\
        );

    \I__1510\ : InMux
    port map (
            O => \N__8325\,
            I => \N__8319\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__8322\,
            I => \DUT.uart_inst0.rx_clk_divider_1_13\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__8319\,
            I => \DUT.uart_inst0.rx_clk_divider_1_13\
        );

    \I__1507\ : InMux
    port map (
            O => \N__8314\,
            I => \N__8311\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__8311\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_13\
        );

    \I__1505\ : InMux
    port map (
            O => \N__8308\,
            I => \N__8305\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__8305\,
            I => \N__8302\
        );

    \I__1503\ : Span4Mux_h
    port map (
            O => \N__8302\,
            I => \N__8299\
        );

    \I__1502\ : Odrv4
    port map (
            O => \N__8299\,
            I => \DUT.uart_inst0.N_199_0\
        );

    \I__1501\ : IoInMux
    port map (
            O => \N__8296\,
            I => \N__8293\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__8293\,
            I => \N__8290\
        );

    \I__1499\ : IoSpan4Mux
    port map (
            O => \N__8290\,
            I => \N__8287\
        );

    \I__1498\ : Odrv4
    port map (
            O => \N__8287\,
            I => \N_1239_i\
        );

    \I__1497\ : CascadeMux
    port map (
            O => \N__8284\,
            I => \N__8281\
        );

    \I__1496\ : InMux
    port map (
            O => \N__8281\,
            I => \N__8276\
        );

    \I__1495\ : InMux
    port map (
            O => \N__8280\,
            I => \N__8273\
        );

    \I__1494\ : InMux
    port map (
            O => \N__8279\,
            I => \N__8270\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__8276\,
            I => \N__8265\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__8273\,
            I => \N__8265\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__8270\,
            I => \DUT.uart_inst0.recv_stateZ0Z_0\
        );

    \I__1490\ : Odrv12
    port map (
            O => \N__8265\,
            I => \DUT.uart_inst0.recv_stateZ0Z_0\
        );

    \I__1489\ : CascadeMux
    port map (
            O => \N__8260\,
            I => \N__8257\
        );

    \I__1488\ : InMux
    port map (
            O => \N__8257\,
            I => \N__8253\
        );

    \I__1487\ : InMux
    port map (
            O => \N__8256\,
            I => \N__8250\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__8253\,
            I => \N__8247\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__8250\,
            I => \N__8244\
        );

    \I__1484\ : Span4Mux_h
    port map (
            O => \N__8247\,
            I => \N__8241\
        );

    \I__1483\ : Odrv4
    port map (
            O => \N__8244\,
            I => \DUT.uart_inst0.rx_clk_divider_5_i_a2_12_1_5\
        );

    \I__1482\ : Odrv4
    port map (
            O => \N__8241\,
            I => \DUT.uart_inst0.rx_clk_divider_5_i_a2_12_1_5\
        );

    \I__1481\ : InMux
    port map (
            O => \N__8236\,
            I => \N__8231\
        );

    \I__1480\ : InMux
    port map (
            O => \N__8235\,
            I => \N__8226\
        );

    \I__1479\ : InMux
    port map (
            O => \N__8234\,
            I => \N__8226\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__8231\,
            I => \DUT.uart_inst0.rx_clk_divider_1_16\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__8226\,
            I => \DUT.uart_inst0.rx_clk_divider_1_16\
        );

    \I__1476\ : CascadeMux
    port map (
            O => \N__8221\,
            I => \N__8217\
        );

    \I__1475\ : InMux
    port map (
            O => \N__8220\,
            I => \N__8214\
        );

    \I__1474\ : InMux
    port map (
            O => \N__8217\,
            I => \N__8211\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__8214\,
            I => \N__8208\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__8211\,
            I => \N__8205\
        );

    \I__1471\ : Span4Mux_h
    port map (
            O => \N__8208\,
            I => \N__8202\
        );

    \I__1470\ : Odrv4
    port map (
            O => \N__8205\,
            I => \DUT.uart_inst0.rx_clk_divider_5_i_a2_12_4_5\
        );

    \I__1469\ : Odrv4
    port map (
            O => \N__8202\,
            I => \DUT.uart_inst0.rx_clk_divider_5_i_a2_12_4_5\
        );

    \I__1468\ : InMux
    port map (
            O => \N__8197\,
            I => \N__8192\
        );

    \I__1467\ : InMux
    port map (
            O => \N__8196\,
            I => \N__8187\
        );

    \I__1466\ : InMux
    port map (
            O => \N__8195\,
            I => \N__8187\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__8192\,
            I => \DUT.uart_inst0.rx_clk_divider_1_14\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__8187\,
            I => \DUT.uart_inst0.rx_clk_divider_1_14\
        );

    \I__1463\ : InMux
    port map (
            O => \N__8182\,
            I => \N__8176\
        );

    \I__1462\ : InMux
    port map (
            O => \N__8181\,
            I => \N__8176\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__8176\,
            I => \N__8173\
        );

    \I__1460\ : Span4Mux_s2_v
    port map (
            O => \N__8173\,
            I => \N__8170\
        );

    \I__1459\ : Odrv4
    port map (
            O => \N__8170\,
            I => \DUT.uart_inst0.rx_clk_divider_5_i_a2_12_5\
        );

    \I__1458\ : CascadeMux
    port map (
            O => \N__8167\,
            I => \N__8163\
        );

    \I__1457\ : CascadeMux
    port map (
            O => \N__8166\,
            I => \N__8160\
        );

    \I__1456\ : InMux
    port map (
            O => \N__8163\,
            I => \N__8155\
        );

    \I__1455\ : InMux
    port map (
            O => \N__8160\,
            I => \N__8155\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__8155\,
            I => \DUT.uart_inst0.rx_clk_divider_1_9\
        );

    \I__1453\ : InMux
    port map (
            O => \N__8152\,
            I => \N__8149\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__8149\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_9\
        );

    \I__1451\ : InMux
    port map (
            O => \N__8146\,
            I => \N__8140\
        );

    \I__1450\ : InMux
    port map (
            O => \N__8145\,
            I => \N__8140\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__8140\,
            I => \DUT.uart_inst0.rx_clk_divider_1_11\
        );

    \I__1448\ : InMux
    port map (
            O => \N__8137\,
            I => \N__8134\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__8134\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_11\
        );

    \I__1446\ : InMux
    port map (
            O => \N__8131\,
            I => \N__8125\
        );

    \I__1445\ : InMux
    port map (
            O => \N__8130\,
            I => \N__8125\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__8125\,
            I => \DUT.uart_inst0.rx_clk_divider_1_12\
        );

    \I__1443\ : InMux
    port map (
            O => \N__8122\,
            I => \N__8119\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__8119\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_12\
        );

    \I__1441\ : CascadeMux
    port map (
            O => \N__8116\,
            I => \N__8111\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__8115\,
            I => \N__8108\
        );

    \I__1439\ : InMux
    port map (
            O => \N__8114\,
            I => \N__8103\
        );

    \I__1438\ : InMux
    port map (
            O => \N__8111\,
            I => \N__8103\
        );

    \I__1437\ : InMux
    port map (
            O => \N__8108\,
            I => \N__8100\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__8103\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_1\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__8100\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_1\
        );

    \I__1434\ : InMux
    port map (
            O => \N__8095\,
            I => \N__8092\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__8092\,
            I => \N__8088\
        );

    \I__1432\ : InMux
    port map (
            O => \N__8091\,
            I => \N__8085\
        );

    \I__1431\ : Odrv4
    port map (
            O => \N__8088\,
            I => \DUT.uart_inst0.rx_clk_divider_1_7\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__8085\,
            I => \DUT.uart_inst0.rx_clk_divider_1_7\
        );

    \I__1429\ : InMux
    port map (
            O => \N__8080\,
            I => \N__8074\
        );

    \I__1428\ : InMux
    port map (
            O => \N__8079\,
            I => \N__8074\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__8074\,
            I => \DUT.uart_inst0.rx_clk_divider_1_1\
        );

    \I__1426\ : CascadeMux
    port map (
            O => \N__8071\,
            I => \N__8068\
        );

    \I__1425\ : InMux
    port map (
            O => \N__8068\,
            I => \N__8065\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__8065\,
            I => \DUT.uart_inst0.rx_clk_dividerZ1Z_1\
        );

    \I__1423\ : InMux
    port map (
            O => \N__8062\,
            I => \N__8059\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__8059\,
            I => \N__8056\
        );

    \I__1421\ : Span4Mux_h
    port map (
            O => \N__8056\,
            I => \N__8053\
        );

    \I__1420\ : Odrv4
    port map (
            O => \N__8053\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_5\
        );

    \I__1419\ : InMux
    port map (
            O => \N__8050\,
            I => \N__8047\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__8047\,
            I => \N__8043\
        );

    \I__1417\ : InMux
    port map (
            O => \N__8046\,
            I => \N__8040\
        );

    \I__1416\ : Span4Mux_s2_v
    port map (
            O => \N__8043\,
            I => \N__8036\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__8040\,
            I => \N__8033\
        );

    \I__1414\ : CascadeMux
    port map (
            O => \N__8039\,
            I => \N__8023\
        );

    \I__1413\ : Span4Mux_h
    port map (
            O => \N__8036\,
            I => \N__8017\
        );

    \I__1412\ : Span4Mux_s2_v
    port map (
            O => \N__8033\,
            I => \N__8017\
        );

    \I__1411\ : InMux
    port map (
            O => \N__8032\,
            I => \N__8012\
        );

    \I__1410\ : InMux
    port map (
            O => \N__8031\,
            I => \N__8012\
        );

    \I__1409\ : InMux
    port map (
            O => \N__8030\,
            I => \N__8005\
        );

    \I__1408\ : InMux
    port map (
            O => \N__8029\,
            I => \N__8005\
        );

    \I__1407\ : InMux
    port map (
            O => \N__8028\,
            I => \N__8005\
        );

    \I__1406\ : InMux
    port map (
            O => \N__8027\,
            I => \N__8002\
        );

    \I__1405\ : InMux
    port map (
            O => \N__8026\,
            I => \N__7995\
        );

    \I__1404\ : InMux
    port map (
            O => \N__8023\,
            I => \N__7995\
        );

    \I__1403\ : InMux
    port map (
            O => \N__8022\,
            I => \N__7995\
        );

    \I__1402\ : Odrv4
    port map (
            O => \N__8017\,
            I => \DUT.uart_inst0.rx_countdown_3_1\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__8012\,
            I => \DUT.uart_inst0.rx_countdown_3_1\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__8005\,
            I => \DUT.uart_inst0.rx_countdown_3_1\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__8002\,
            I => \DUT.uart_inst0.rx_countdown_3_1\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__7995\,
            I => \DUT.uart_inst0.rx_countdown_3_1\
        );

    \I__1397\ : InMux
    port map (
            O => \N__7984\,
            I => \N__7981\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__7981\,
            I => \N__7978\
        );

    \I__1395\ : Span4Mux_h
    port map (
            O => \N__7978\,
            I => \N__7975\
        );

    \I__1394\ : Odrv4
    port map (
            O => \N__7975\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_1\
        );

    \I__1393\ : InMux
    port map (
            O => \N__7972\,
            I => \N__7969\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__7969\,
            I => \N__7965\
        );

    \I__1391\ : InMux
    port map (
            O => \N__7968\,
            I => \N__7962\
        );

    \I__1390\ : Odrv4
    port map (
            O => \N__7965\,
            I => \DUT.uart_inst0.rx_clk_divider_1_2\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__7962\,
            I => \DUT.uart_inst0.rx_clk_divider_1_2\
        );

    \I__1388\ : CascadeMux
    port map (
            O => \N__7957\,
            I => \N__7954\
        );

    \I__1387\ : InMux
    port map (
            O => \N__7954\,
            I => \N__7951\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__7951\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_2\
        );

    \I__1385\ : CEMux
    port map (
            O => \N__7948\,
            I => \N__7945\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__7945\,
            I => \N__7942\
        );

    \I__1383\ : Span4Mux_h
    port map (
            O => \N__7942\,
            I => \N__7938\
        );

    \I__1382\ : InMux
    port map (
            O => \N__7941\,
            I => \N__7935\
        );

    \I__1381\ : Odrv4
    port map (
            O => \N__7938\,
            I => \DUT.fifo_tx_inst.rFifoData_awe2\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__7935\,
            I => \DUT.fifo_tx_inst.rFifoData_awe2\
        );

    \I__1379\ : InMux
    port map (
            O => \N__7930\,
            I => \N__7926\
        );

    \I__1378\ : InMux
    port map (
            O => \N__7929\,
            I => \N__7923\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__7926\,
            I => \N__7920\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__7923\,
            I => \DUT.fifo_tx_inst.rFifoDataro_2\
        );

    \I__1375\ : Odrv4
    port map (
            O => \N__7920\,
            I => \DUT.fifo_tx_inst.rFifoDataro_2\
        );

    \I__1374\ : InMux
    port map (
            O => \N__7915\,
            I => \N__7908\
        );

    \I__1373\ : InMux
    port map (
            O => \N__7914\,
            I => \N__7908\
        );

    \I__1372\ : InMux
    port map (
            O => \N__7913\,
            I => \N__7905\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__7908\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__7905\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4\
        );

    \I__1369\ : CascadeMux
    port map (
            O => \N__7900\,
            I => \N__7897\
        );

    \I__1368\ : InMux
    port map (
            O => \N__7897\,
            I => \N__7890\
        );

    \I__1367\ : InMux
    port map (
            O => \N__7896\,
            I => \N__7890\
        );

    \I__1366\ : InMux
    port map (
            O => \N__7895\,
            I => \N__7887\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__7890\,
            I => \fifo_inst.ftdi_output_inst.rWrDelayZ0\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__7887\,
            I => \fifo_inst.ftdi_output_inst.rWrDelayZ0\
        );

    \I__1363\ : InMux
    port map (
            O => \N__7882\,
            I => \N__7876\
        );

    \I__1362\ : InMux
    port map (
            O => \N__7881\,
            I => \N__7876\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__7876\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_3\
        );

    \I__1360\ : IoInMux
    port map (
            O => \N__7873\,
            I => \N__7870\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__7870\,
            I => \N__7866\
        );

    \I__1358\ : IoInMux
    port map (
            O => \N__7869\,
            I => \N__7863\
        );

    \I__1357\ : Span4Mux_s3_v
    port map (
            O => \N__7866\,
            I => \N__7860\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__7863\,
            I => \N__7857\
        );

    \I__1355\ : Span4Mux_v
    port map (
            O => \N__7860\,
            I => \N__7854\
        );

    \I__1354\ : Span12Mux_s7_v
    port map (
            O => \N__7857\,
            I => \N__7851\
        );

    \I__1353\ : Span4Mux_h
    port map (
            O => \N__7854\,
            I => \N__7848\
        );

    \I__1352\ : Span12Mux_v
    port map (
            O => \N__7851\,
            I => \N__7844\
        );

    \I__1351\ : Span4Mux_h
    port map (
            O => \N__7848\,
            I => \N__7841\
        );

    \I__1350\ : InMux
    port map (
            O => \N__7847\,
            I => \N__7838\
        );

    \I__1349\ : Odrv12
    port map (
            O => \N__7844\,
            I => \P1A4_c\
        );

    \I__1348\ : Odrv4
    port map (
            O => \N__7841\,
            I => \P1A4_c\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__7838\,
            I => \P1A4_c\
        );

    \I__1346\ : IoInMux
    port map (
            O => \N__7831\,
            I => \N__7826\
        );

    \I__1345\ : IoInMux
    port map (
            O => \N__7830\,
            I => \N__7823\
        );

    \I__1344\ : IoInMux
    port map (
            O => \N__7829\,
            I => \N__7820\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__7826\,
            I => \N__7814\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__7823\,
            I => \N__7814\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__7820\,
            I => \N__7811\
        );

    \I__1340\ : IoInMux
    port map (
            O => \N__7819\,
            I => \N__7808\
        );

    \I__1339\ : Span4Mux_s3_v
    port map (
            O => \N__7814\,
            I => \N__7805\
        );

    \I__1338\ : IoSpan4Mux
    port map (
            O => \N__7811\,
            I => \N__7802\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__7808\,
            I => \N__7799\
        );

    \I__1336\ : Span4Mux_h
    port map (
            O => \N__7805\,
            I => \N__7796\
        );

    \I__1335\ : Span4Mux_s2_v
    port map (
            O => \N__7802\,
            I => \N__7791\
        );

    \I__1334\ : Span4Mux_s2_v
    port map (
            O => \N__7799\,
            I => \N__7791\
        );

    \I__1333\ : Sp12to4
    port map (
            O => \N__7796\,
            I => \N__7788\
        );

    \I__1332\ : Span4Mux_v
    port map (
            O => \N__7791\,
            I => \N__7785\
        );

    \I__1331\ : Span12Mux_v
    port map (
            O => \N__7788\,
            I => \N__7781\
        );

    \I__1330\ : Span4Mux_v
    port map (
            O => \N__7785\,
            I => \N__7778\
        );

    \I__1329\ : InMux
    port map (
            O => \N__7784\,
            I => \N__7775\
        );

    \I__1328\ : Odrv12
    port map (
            O => \N__7781\,
            I => \rTxBusReady\
        );

    \I__1327\ : Odrv4
    port map (
            O => \N__7778\,
            I => \rTxBusReady\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__7775\,
            I => \rTxBusReady\
        );

    \I__1325\ : InMux
    port map (
            O => \N__7768\,
            I => \N__7762\
        );

    \I__1324\ : InMux
    port map (
            O => \N__7767\,
            I => \N__7762\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__7762\,
            I => \DUT.uart_inst0.rx_clk_divider_1_8\
        );

    \I__1322\ : InMux
    port map (
            O => \N__7759\,
            I => \N__7756\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__7756\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_8\
        );

    \I__1320\ : InMux
    port map (
            O => \N__7753\,
            I => \N__7750\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__7750\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_6\
        );

    \I__1318\ : CascadeMux
    port map (
            O => \N__7747\,
            I => \N__7744\
        );

    \I__1317\ : InMux
    port map (
            O => \N__7744\,
            I => \N__7741\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__7741\,
            I => \N__7738\
        );

    \I__1315\ : Span4Mux_h
    port map (
            O => \N__7738\,
            I => \N__7735\
        );

    \I__1314\ : Span4Mux_h
    port map (
            O => \N__7735\,
            I => \N__7732\
        );

    \I__1313\ : Odrv4
    port map (
            O => \N__7732\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_6\
        );

    \I__1312\ : InMux
    port map (
            O => \N__7729\,
            I => \N__7725\
        );

    \I__1311\ : InMux
    port map (
            O => \N__7728\,
            I => \N__7722\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__7725\,
            I => \DUT.fifo_tx_inst.rFifoDataro_3\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__7722\,
            I => \DUT.fifo_tx_inst.rFifoDataro_3\
        );

    \I__1308\ : InMux
    port map (
            O => \N__7717\,
            I => \N__7713\
        );

    \I__1307\ : InMux
    port map (
            O => \N__7716\,
            I => \N__7710\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__7713\,
            I => \DUT.fifo_tx_inst.rFifoDataro_0\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__7710\,
            I => \DUT.fifo_tx_inst.rFifoDataro_0\
        );

    \I__1304\ : CascadeMux
    port map (
            O => \N__7705\,
            I => \N__7701\
        );

    \I__1303\ : InMux
    port map (
            O => \N__7704\,
            I => \N__7698\
        );

    \I__1302\ : InMux
    port map (
            O => \N__7701\,
            I => \N__7695\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__7698\,
            I => \DUT.fifo_tx_inst.rFifoDataro_1\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__7695\,
            I => \DUT.fifo_tx_inst.rFifoDataro_1\
        );

    \I__1299\ : InMux
    port map (
            O => \N__7690\,
            I => \N__7687\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__7687\,
            I => \DUT.rFifoDataror_0_0_0\
        );

    \I__1297\ : CascadeMux
    port map (
            O => \N__7684\,
            I => \DUT.rFifoDataror_1_0_cascade_\
        );

    \I__1296\ : InMux
    port map (
            O => \N__7681\,
            I => \N__7678\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__7678\,
            I => \N__7675\
        );

    \I__1294\ : Odrv4
    port map (
            O => \N__7675\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_6\
        );

    \I__1293\ : CascadeMux
    port map (
            O => \N__7672\,
            I => \N__7669\
        );

    \I__1292\ : InMux
    port map (
            O => \N__7669\,
            I => \N__7666\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__7666\,
            I => \N__7663\
        );

    \I__1290\ : Odrv12
    port map (
            O => \N__7663\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_6\
        );

    \I__1289\ : InMux
    port map (
            O => \N__7660\,
            I => \N__7657\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__7657\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6\
        );

    \I__1287\ : CascadeMux
    port map (
            O => \N__7654\,
            I => \N__7649\
        );

    \I__1286\ : CascadeMux
    port map (
            O => \N__7653\,
            I => \N__7643\
        );

    \I__1285\ : InMux
    port map (
            O => \N__7652\,
            I => \N__7640\
        );

    \I__1284\ : InMux
    port map (
            O => \N__7649\,
            I => \N__7631\
        );

    \I__1283\ : InMux
    port map (
            O => \N__7648\,
            I => \N__7631\
        );

    \I__1282\ : InMux
    port map (
            O => \N__7647\,
            I => \N__7631\
        );

    \I__1281\ : InMux
    port map (
            O => \N__7646\,
            I => \N__7631\
        );

    \I__1280\ : InMux
    port map (
            O => \N__7643\,
            I => \N__7628\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__7640\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_0\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__7631\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_0\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__7628\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_0\
        );

    \I__1276\ : CascadeMux
    port map (
            O => \N__7621\,
            I => \DUT.fifo_tx_inst.N_79_cascade_\
        );

    \I__1275\ : CascadeMux
    port map (
            O => \N__7618\,
            I => \N__7613\
        );

    \I__1274\ : InMux
    port map (
            O => \N__7617\,
            I => \N__7608\
        );

    \I__1273\ : InMux
    port map (
            O => \N__7616\,
            I => \N__7605\
        );

    \I__1272\ : InMux
    port map (
            O => \N__7613\,
            I => \N__7598\
        );

    \I__1271\ : InMux
    port map (
            O => \N__7612\,
            I => \N__7598\
        );

    \I__1270\ : InMux
    port map (
            O => \N__7611\,
            I => \N__7598\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__7608\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_1\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__7605\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_1\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__7598\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_1\
        );

    \I__1266\ : InMux
    port map (
            O => \N__7591\,
            I => \N__7587\
        );

    \I__1265\ : InMux
    port map (
            O => \N__7590\,
            I => \N__7584\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__7587\,
            I => \N__7579\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__7584\,
            I => \N__7576\
        );

    \I__1262\ : InMux
    port map (
            O => \N__7583\,
            I => \N__7573\
        );

    \I__1261\ : InMux
    port map (
            O => \N__7582\,
            I => \N__7570\
        );

    \I__1260\ : Span4Mux_v
    port map (
            O => \N__7579\,
            I => \N__7563\
        );

    \I__1259\ : Span4Mux_h
    port map (
            O => \N__7576\,
            I => \N__7563\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__7573\,
            I => \N__7563\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__7570\,
            I => \N__7560\
        );

    \I__1256\ : Odrv4
    port map (
            O => \N__7563\,
            I => \rTxByteZ0Z_6\
        );

    \I__1255\ : Odrv4
    port map (
            O => \N__7560\,
            I => \rTxByteZ0Z_6\
        );

    \I__1254\ : InMux
    port map (
            O => \N__7555\,
            I => \N__7552\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__7552\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_4\
        );

    \I__1252\ : InMux
    port map (
            O => \N__7549\,
            I => \N__7546\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__7546\,
            I => \N__7543\
        );

    \I__1250\ : Odrv4
    port map (
            O => \N__7543\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_4\
        );

    \I__1249\ : CascadeMux
    port map (
            O => \N__7540\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_\
        );

    \I__1248\ : InMux
    port map (
            O => \N__7537\,
            I => \N__7534\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__7534\,
            I => \N__7531\
        );

    \I__1246\ : Odrv4
    port map (
            O => \N__7531\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_4\
        );

    \I__1245\ : InMux
    port map (
            O => \N__7528\,
            I => \N__7523\
        );

    \I__1244\ : InMux
    port map (
            O => \N__7527\,
            I => \N__7520\
        );

    \I__1243\ : InMux
    port map (
            O => \N__7526\,
            I => \N__7517\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__7523\,
            I => \N__7513\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__7520\,
            I => \N__7510\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__7517\,
            I => \N__7507\
        );

    \I__1239\ : InMux
    port map (
            O => \N__7516\,
            I => \N__7504\
        );

    \I__1238\ : Span4Mux_v
    port map (
            O => \N__7513\,
            I => \N__7495\
        );

    \I__1237\ : Span4Mux_v
    port map (
            O => \N__7510\,
            I => \N__7495\
        );

    \I__1236\ : Span4Mux_h
    port map (
            O => \N__7507\,
            I => \N__7495\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__7504\,
            I => \N__7495\
        );

    \I__1234\ : Odrv4
    port map (
            O => \N__7495\,
            I => \rTxByteZ0Z_4\
        );

    \I__1233\ : CascadeMux
    port map (
            O => \N__7492\,
            I => \N__7489\
        );

    \I__1232\ : InMux
    port map (
            O => \N__7489\,
            I => \N__7486\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__7486\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_4\
        );

    \I__1230\ : InMux
    port map (
            O => \N__7483\,
            I => \N__7480\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__7480\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_5\
        );

    \I__1228\ : InMux
    port map (
            O => \N__7477\,
            I => \N__7474\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__7474\,
            I => \N__7471\
        );

    \I__1226\ : Odrv4
    port map (
            O => \N__7471\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_5\
        );

    \I__1225\ : InMux
    port map (
            O => \N__7468\,
            I => \N__7465\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__7465\,
            I => \N__7462\
        );

    \I__1223\ : Odrv4
    port map (
            O => \N__7462\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_5\
        );

    \I__1222\ : CascadeMux
    port map (
            O => \N__7459\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_\
        );

    \I__1221\ : InMux
    port map (
            O => \N__7456\,
            I => \N__7452\
        );

    \I__1220\ : InMux
    port map (
            O => \N__7455\,
            I => \N__7449\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__7452\,
            I => \N__7445\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__7449\,
            I => \N__7442\
        );

    \I__1217\ : InMux
    port map (
            O => \N__7448\,
            I => \N__7439\
        );

    \I__1216\ : Span4Mux_v
    port map (
            O => \N__7445\,
            I => \N__7433\
        );

    \I__1215\ : Span4Mux_v
    port map (
            O => \N__7442\,
            I => \N__7433\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__7439\,
            I => \N__7430\
        );

    \I__1213\ : InMux
    port map (
            O => \N__7438\,
            I => \N__7427\
        );

    \I__1212\ : Odrv4
    port map (
            O => \N__7433\,
            I => \rTxByteZ0Z_5\
        );

    \I__1211\ : Odrv4
    port map (
            O => \N__7430\,
            I => \rTxByteZ0Z_5\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__7427\,
            I => \rTxByteZ0Z_5\
        );

    \I__1209\ : InMux
    port map (
            O => \N__7420\,
            I => \N__7417\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__7417\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_5\
        );

    \I__1207\ : CEMux
    port map (
            O => \N__7414\,
            I => \N__7409\
        );

    \I__1206\ : CEMux
    port map (
            O => \N__7413\,
            I => \N__7406\
        );

    \I__1205\ : CEMux
    port map (
            O => \N__7412\,
            I => \N__7403\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__7409\,
            I => \N__7400\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__7406\,
            I => \N__7397\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__7403\,
            I => \N__7394\
        );

    \I__1201\ : Span4Mux_h
    port map (
            O => \N__7400\,
            I => \N__7390\
        );

    \I__1200\ : Span4Mux_v
    port map (
            O => \N__7397\,
            I => \N__7387\
        );

    \I__1199\ : Span4Mux_h
    port map (
            O => \N__7394\,
            I => \N__7384\
        );

    \I__1198\ : InMux
    port map (
            O => \N__7393\,
            I => \N__7381\
        );

    \I__1197\ : Odrv4
    port map (
            O => \N__7390\,
            I => \DUT.fifo_tx_inst.rFifoData_awe3\
        );

    \I__1196\ : Odrv4
    port map (
            O => \N__7387\,
            I => \DUT.fifo_tx_inst.rFifoData_awe3\
        );

    \I__1195\ : Odrv4
    port map (
            O => \N__7384\,
            I => \DUT.fifo_tx_inst.rFifoData_awe3\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__7381\,
            I => \DUT.fifo_tx_inst.rFifoData_awe3\
        );

    \I__1193\ : InMux
    port map (
            O => \N__7372\,
            I => \N__7367\
        );

    \I__1192\ : InMux
    port map (
            O => \N__7371\,
            I => \N__7364\
        );

    \I__1191\ : InMux
    port map (
            O => \N__7370\,
            I => \N__7361\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__7367\,
            I => \N__7357\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__7364\,
            I => \N__7354\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__7361\,
            I => \N__7351\
        );

    \I__1187\ : InMux
    port map (
            O => \N__7360\,
            I => \N__7348\
        );

    \I__1186\ : Span4Mux_v
    port map (
            O => \N__7357\,
            I => \N__7339\
        );

    \I__1185\ : Span4Mux_v
    port map (
            O => \N__7354\,
            I => \N__7339\
        );

    \I__1184\ : Span4Mux_h
    port map (
            O => \N__7351\,
            I => \N__7339\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__7348\,
            I => \N__7339\
        );

    \I__1182\ : Odrv4
    port map (
            O => \N__7339\,
            I => \rTxByteZ0Z_0\
        );

    \I__1181\ : InMux
    port map (
            O => \N__7336\,
            I => \N__7333\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__7333\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_0\
        );

    \I__1179\ : InMux
    port map (
            O => \N__7330\,
            I => \N__7326\
        );

    \I__1178\ : InMux
    port map (
            O => \N__7329\,
            I => \N__7323\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__7326\,
            I => \N__7319\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__7323\,
            I => \N__7316\
        );

    \I__1175\ : InMux
    port map (
            O => \N__7322\,
            I => \N__7313\
        );

    \I__1174\ : Span4Mux_h
    port map (
            O => \N__7319\,
            I => \N__7309\
        );

    \I__1173\ : Span4Mux_v
    port map (
            O => \N__7316\,
            I => \N__7304\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__7313\,
            I => \N__7304\
        );

    \I__1171\ : InMux
    port map (
            O => \N__7312\,
            I => \N__7301\
        );

    \I__1170\ : Odrv4
    port map (
            O => \N__7309\,
            I => \rTxByteZ0Z_1\
        );

    \I__1169\ : Odrv4
    port map (
            O => \N__7304\,
            I => \rTxByteZ0Z_1\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__7301\,
            I => \rTxByteZ0Z_1\
        );

    \I__1167\ : InMux
    port map (
            O => \N__7294\,
            I => \N__7291\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__7291\,
            I => \N__7286\
        );

    \I__1165\ : InMux
    port map (
            O => \N__7290\,
            I => \N__7283\
        );

    \I__1164\ : InMux
    port map (
            O => \N__7289\,
            I => \N__7280\
        );

    \I__1163\ : Span4Mux_h
    port map (
            O => \N__7286\,
            I => \N__7276\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__7283\,
            I => \N__7273\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__7280\,
            I => \N__7270\
        );

    \I__1160\ : InMux
    port map (
            O => \N__7279\,
            I => \N__7267\
        );

    \I__1159\ : Odrv4
    port map (
            O => \N__7276\,
            I => \rTxByteZ0Z_3\
        );

    \I__1158\ : Odrv4
    port map (
            O => \N__7273\,
            I => \rTxByteZ0Z_3\
        );

    \I__1157\ : Odrv4
    port map (
            O => \N__7270\,
            I => \rTxByteZ0Z_3\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__7267\,
            I => \rTxByteZ0Z_3\
        );

    \I__1155\ : InMux
    port map (
            O => \N__7258\,
            I => \N__7255\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__7255\,
            I => \DUT.uart_inst0.G_11_i_a4_0_4\
        );

    \I__1153\ : InMux
    port map (
            O => \N__7252\,
            I => \N__7249\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__7249\,
            I => \DUT.uart_inst0.N_4_i_1\
        );

    \I__1151\ : InMux
    port map (
            O => \N__7246\,
            I => \N__7242\
        );

    \I__1150\ : InMux
    port map (
            O => \N__7245\,
            I => \N__7238\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__7242\,
            I => \N__7234\
        );

    \I__1148\ : InMux
    port map (
            O => \N__7241\,
            I => \N__7231\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__7238\,
            I => \N__7228\
        );

    \I__1146\ : InMux
    port map (
            O => \N__7237\,
            I => \N__7225\
        );

    \I__1145\ : Span4Mux_v
    port map (
            O => \N__7234\,
            I => \N__7220\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__7231\,
            I => \N__7220\
        );

    \I__1143\ : Span4Mux_h
    port map (
            O => \N__7228\,
            I => \N__7215\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__7225\,
            I => \N__7215\
        );

    \I__1141\ : Span4Mux_h
    port map (
            O => \N__7220\,
            I => \N__7211\
        );

    \I__1140\ : Span4Mux_v
    port map (
            O => \N__7215\,
            I => \N__7208\
        );

    \I__1139\ : InMux
    port map (
            O => \N__7214\,
            I => \N__7205\
        );

    \I__1138\ : Odrv4
    port map (
            O => \N__7211\,
            I => \DUT.wRxByte_1\
        );

    \I__1137\ : Odrv4
    port map (
            O => \N__7208\,
            I => \DUT.wRxByte_1\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__7205\,
            I => \DUT.wRxByte_1\
        );

    \I__1135\ : InMux
    port map (
            O => \N__7198\,
            I => \N__7195\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__7195\,
            I => \N__7189\
        );

    \I__1133\ : InMux
    port map (
            O => \N__7194\,
            I => \N__7186\
        );

    \I__1132\ : InMux
    port map (
            O => \N__7193\,
            I => \N__7183\
        );

    \I__1131\ : InMux
    port map (
            O => \N__7192\,
            I => \N__7180\
        );

    \I__1130\ : Span4Mux_v
    port map (
            O => \N__7189\,
            I => \N__7173\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__7186\,
            I => \N__7173\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__7183\,
            I => \N__7173\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__7180\,
            I => \N__7170\
        );

    \I__1126\ : Span4Mux_v
    port map (
            O => \N__7173\,
            I => \N__7167\
        );

    \I__1125\ : Span4Mux_h
    port map (
            O => \N__7170\,
            I => \N__7164\
        );

    \I__1124\ : Odrv4
    port map (
            O => \N__7167\,
            I => \DUT.wRxByte_0\
        );

    \I__1123\ : Odrv4
    port map (
            O => \N__7164\,
            I => \DUT.wRxByte_0\
        );

    \I__1122\ : InMux
    port map (
            O => \N__7159\,
            I => \N__7155\
        );

    \I__1121\ : InMux
    port map (
            O => \N__7158\,
            I => \N__7152\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__7155\,
            I => \N__7145\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__7152\,
            I => \N__7145\
        );

    \I__1118\ : InMux
    port map (
            O => \N__7151\,
            I => \N__7142\
        );

    \I__1117\ : InMux
    port map (
            O => \N__7150\,
            I => \N__7139\
        );

    \I__1116\ : Span4Mux_v
    port map (
            O => \N__7145\,
            I => \N__7134\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__7142\,
            I => \N__7134\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__7139\,
            I => \N__7131\
        );

    \I__1113\ : Span4Mux_v
    port map (
            O => \N__7134\,
            I => \N__7127\
        );

    \I__1112\ : Span4Mux_v
    port map (
            O => \N__7131\,
            I => \N__7124\
        );

    \I__1111\ : InMux
    port map (
            O => \N__7130\,
            I => \N__7121\
        );

    \I__1110\ : Odrv4
    port map (
            O => \N__7127\,
            I => \DUT.wRxByte_4\
        );

    \I__1109\ : Odrv4
    port map (
            O => \N__7124\,
            I => \DUT.wRxByte_4\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__7121\,
            I => \DUT.wRxByte_4\
        );

    \I__1107\ : InMux
    port map (
            O => \N__7114\,
            I => \N__7110\
        );

    \I__1106\ : InMux
    port map (
            O => \N__7113\,
            I => \N__7107\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__7110\,
            I => \N__7100\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__7107\,
            I => \N__7100\
        );

    \I__1103\ : InMux
    port map (
            O => \N__7106\,
            I => \N__7097\
        );

    \I__1102\ : InMux
    port map (
            O => \N__7105\,
            I => \N__7094\
        );

    \I__1101\ : Span4Mux_v
    port map (
            O => \N__7100\,
            I => \N__7089\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__7097\,
            I => \N__7089\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__7094\,
            I => \N__7086\
        );

    \I__1098\ : Span4Mux_v
    port map (
            O => \N__7089\,
            I => \N__7082\
        );

    \I__1097\ : Span4Mux_v
    port map (
            O => \N__7086\,
            I => \N__7079\
        );

    \I__1096\ : InMux
    port map (
            O => \N__7085\,
            I => \N__7076\
        );

    \I__1095\ : Odrv4
    port map (
            O => \N__7082\,
            I => \DUT.wRxByte_5\
        );

    \I__1094\ : Odrv4
    port map (
            O => \N__7079\,
            I => \DUT.wRxByte_5\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__7076\,
            I => \DUT.wRxByte_5\
        );

    \I__1092\ : InMux
    port map (
            O => \N__7069\,
            I => \N__7065\
        );

    \I__1091\ : InMux
    port map (
            O => \N__7068\,
            I => \N__7062\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__7065\,
            I => \N__7058\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__7062\,
            I => \N__7055\
        );

    \I__1088\ : InMux
    port map (
            O => \N__7061\,
            I => \N__7052\
        );

    \I__1087\ : Span4Mux_v
    port map (
            O => \N__7058\,
            I => \N__7044\
        );

    \I__1086\ : Span4Mux_h
    port map (
            O => \N__7055\,
            I => \N__7044\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__7052\,
            I => \N__7044\
        );

    \I__1084\ : InMux
    port map (
            O => \N__7051\,
            I => \N__7041\
        );

    \I__1083\ : Span4Mux_v
    port map (
            O => \N__7044\,
            I => \N__7037\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__7041\,
            I => \N__7034\
        );

    \I__1081\ : InMux
    port map (
            O => \N__7040\,
            I => \N__7031\
        );

    \I__1080\ : Odrv4
    port map (
            O => \N__7037\,
            I => \DUT.wRxByte_6\
        );

    \I__1079\ : Odrv4
    port map (
            O => \N__7034\,
            I => \DUT.wRxByte_6\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__7031\,
            I => \DUT.wRxByte_6\
        );

    \I__1077\ : InMux
    port map (
            O => \N__7024\,
            I => \N__7019\
        );

    \I__1076\ : InMux
    port map (
            O => \N__7023\,
            I => \N__7016\
        );

    \I__1075\ : InMux
    port map (
            O => \N__7022\,
            I => \N__7013\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__7019\,
            I => \N__7007\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__7016\,
            I => \N__7007\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__7013\,
            I => \N__7004\
        );

    \I__1071\ : InMux
    port map (
            O => \N__7012\,
            I => \N__7001\
        );

    \I__1070\ : Span4Mux_v
    port map (
            O => \N__7007\,
            I => \N__6997\
        );

    \I__1069\ : Span4Mux_h
    port map (
            O => \N__7004\,
            I => \N__6992\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__7001\,
            I => \N__6992\
        );

    \I__1067\ : InMux
    port map (
            O => \N__7000\,
            I => \N__6989\
        );

    \I__1066\ : Odrv4
    port map (
            O => \N__6997\,
            I => \DUT.wRxByte_7\
        );

    \I__1065\ : Odrv4
    port map (
            O => \N__6992\,
            I => \DUT.wRxByte_7\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__6989\,
            I => \DUT.wRxByte_7\
        );

    \I__1063\ : InMux
    port map (
            O => \N__6982\,
            I => \N__6979\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__6979\,
            I => \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa_0_a2_0_a2_0_a3_1\
        );

    \I__1061\ : CascadeMux
    port map (
            O => \N__6976\,
            I => \DUT.uart_inst0.rx_countdown_8_i_0_o2_1_2_2_cascade_\
        );

    \I__1060\ : InMux
    port map (
            O => \N__6973\,
            I => \N__6967\
        );

    \I__1059\ : InMux
    port map (
            O => \N__6972\,
            I => \N__6967\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__6967\,
            I => \DUT.uart_inst0.recv_state_ns_0_i_0_0_o2_0_3\
        );

    \I__1057\ : CascadeMux
    port map (
            O => \N__6964\,
            I => \DUT.uart_inst0.G_9_1_cascade_\
        );

    \I__1056\ : InMux
    port map (
            O => \N__6961\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_11\
        );

    \I__1055\ : InMux
    port map (
            O => \N__6958\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_12\
        );

    \I__1054\ : CascadeMux
    port map (
            O => \N__6955\,
            I => \N__6952\
        );

    \I__1053\ : InMux
    port map (
            O => \N__6952\,
            I => \N__6949\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__6949\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_14\
        );

    \I__1051\ : InMux
    port map (
            O => \N__6946\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_13\
        );

    \I__1050\ : InMux
    port map (
            O => \N__6943\,
            I => \N__6940\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__6940\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_15\
        );

    \I__1048\ : InMux
    port map (
            O => \N__6937\,
            I => \N__6933\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6936\,
            I => \N__6930\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__6933\,
            I => \DUT.uart_inst0.rx_clk_divider_1_15\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__6930\,
            I => \DUT.uart_inst0.rx_clk_divider_1_15\
        );

    \I__1044\ : InMux
    port map (
            O => \N__6925\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_14\
        );

    \I__1043\ : InMux
    port map (
            O => \N__6922\,
            I => \N__6919\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__6919\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_16\
        );

    \I__1041\ : InMux
    port map (
            O => \N__6916\,
            I => \bfn_15_3_0_\
        );

    \I__1040\ : InMux
    port map (
            O => \N__6913\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_16\
        );

    \I__1039\ : CascadeMux
    port map (
            O => \N__6910\,
            I => \DUT.uart_inst0.recv_state_RNO_2Z0Z_4_cascade_\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6907\,
            I => \N__6904\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__6904\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_4\
        );

    \I__1036\ : InMux
    port map (
            O => \N__6901\,
            I => \N__6897\
        );

    \I__1035\ : InMux
    port map (
            O => \N__6900\,
            I => \N__6894\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__6897\,
            I => \DUT.uart_inst0.rx_clk_divider_1_4\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__6894\,
            I => \DUT.uart_inst0.rx_clk_divider_1_4\
        );

    \I__1032\ : InMux
    port map (
            O => \N__6889\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_3\
        );

    \I__1031\ : CascadeMux
    port map (
            O => \N__6886\,
            I => \N__6883\
        );

    \I__1030\ : InMux
    port map (
            O => \N__6883\,
            I => \N__6880\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__6880\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_5\
        );

    \I__1028\ : InMux
    port map (
            O => \N__6877\,
            I => \N__6868\
        );

    \I__1027\ : InMux
    port map (
            O => \N__6876\,
            I => \N__6868\
        );

    \I__1026\ : InMux
    port map (
            O => \N__6875\,
            I => \N__6868\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__6868\,
            I => \DUT.uart_inst0.rx_clk_divider_1_5\
        );

    \I__1024\ : InMux
    port map (
            O => \N__6865\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_4\
        );

    \I__1023\ : InMux
    port map (
            O => \N__6862\,
            I => \N__6859\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__6859\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_6\
        );

    \I__1021\ : CascadeMux
    port map (
            O => \N__6856\,
            I => \N__6851\
        );

    \I__1020\ : CascadeMux
    port map (
            O => \N__6855\,
            I => \N__6848\
        );

    \I__1019\ : InMux
    port map (
            O => \N__6854\,
            I => \N__6845\
        );

    \I__1018\ : InMux
    port map (
            O => \N__6851\,
            I => \N__6840\
        );

    \I__1017\ : InMux
    port map (
            O => \N__6848\,
            I => \N__6840\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__6845\,
            I => \DUT.uart_inst0.rx_clk_divider_1_6\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__6840\,
            I => \DUT.uart_inst0.rx_clk_divider_1_6\
        );

    \I__1014\ : InMux
    port map (
            O => \N__6835\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_5\
        );

    \I__1013\ : InMux
    port map (
            O => \N__6832\,
            I => \N__6829\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__6829\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_7\
        );

    \I__1011\ : InMux
    port map (
            O => \N__6826\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_6\
        );

    \I__1010\ : InMux
    port map (
            O => \N__6823\,
            I => \bfn_15_2_0_\
        );

    \I__1009\ : InMux
    port map (
            O => \N__6820\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_8\
        );

    \I__1008\ : InMux
    port map (
            O => \N__6817\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_9\
        );

    \I__1007\ : InMux
    port map (
            O => \N__6814\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_10\
        );

    \I__1006\ : CascadeMux
    port map (
            O => \N__6811\,
            I => \N__6807\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6810\,
            I => \N__6803\
        );

    \I__1004\ : InMux
    port map (
            O => \N__6807\,
            I => \N__6797\
        );

    \I__1003\ : InMux
    port map (
            O => \N__6806\,
            I => \N__6797\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__6803\,
            I => \N__6794\
        );

    \I__1001\ : InMux
    port map (
            O => \N__6802\,
            I => \N__6791\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__6797\,
            I => \DUT.fifo_rx_inst.N_194\
        );

    \I__999\ : Odrv4
    port map (
            O => \N__6794\,
            I => \DUT.fifo_rx_inst.N_194\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__6791\,
            I => \DUT.fifo_rx_inst.N_194\
        );

    \I__997\ : InMux
    port map (
            O => \N__6784\,
            I => \N__6779\
        );

    \I__996\ : CascadeMux
    port map (
            O => \N__6783\,
            I => \N__6773\
        );

    \I__995\ : InMux
    port map (
            O => \N__6782\,
            I => \N__6770\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__6779\,
            I => \N__6767\
        );

    \I__993\ : InMux
    port map (
            O => \N__6778\,
            I => \N__6764\
        );

    \I__992\ : InMux
    port map (
            O => \N__6777\,
            I => \N__6757\
        );

    \I__991\ : InMux
    port map (
            O => \N__6776\,
            I => \N__6757\
        );

    \I__990\ : InMux
    port map (
            O => \N__6773\,
            I => \N__6757\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__6770\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_0\
        );

    \I__988\ : Odrv4
    port map (
            O => \N__6767\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_0\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__6764\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_0\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__6757\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_0\
        );

    \I__985\ : InMux
    port map (
            O => \N__6748\,
            I => \N__6745\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__6745\,
            I => \N__6738\
        );

    \I__983\ : InMux
    port map (
            O => \N__6744\,
            I => \N__6735\
        );

    \I__982\ : InMux
    port map (
            O => \N__6743\,
            I => \N__6728\
        );

    \I__981\ : InMux
    port map (
            O => \N__6742\,
            I => \N__6728\
        );

    \I__980\ : InMux
    port map (
            O => \N__6741\,
            I => \N__6728\
        );

    \I__979\ : Odrv4
    port map (
            O => \N__6738\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_1\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__6735\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_1\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__6728\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_1\
        );

    \I__976\ : InMux
    port map (
            O => \N__6721\,
            I => \N__6718\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__6718\,
            I => \N__6715\
        );

    \I__974\ : Span4Mux_v
    port map (
            O => \N__6715\,
            I => \N__6712\
        );

    \I__973\ : Odrv4
    port map (
            O => \N__6712\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_5\
        );

    \I__972\ : InMux
    port map (
            O => \N__6709\,
            I => \N__6706\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__6706\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_3\
        );

    \I__970\ : InMux
    port map (
            O => \N__6703\,
            I => \N__6700\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__6700\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_4\
        );

    \I__968\ : CEMux
    port map (
            O => \N__6697\,
            I => \N__6694\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__6694\,
            I => \N__6691\
        );

    \I__966\ : Span4Mux_v
    port map (
            O => \N__6691\,
            I => \N__6686\
        );

    \I__965\ : CEMux
    port map (
            O => \N__6690\,
            I => \N__6683\
        );

    \I__964\ : InMux
    port map (
            O => \N__6689\,
            I => \N__6679\
        );

    \I__963\ : Span4Mux_h
    port map (
            O => \N__6686\,
            I => \N__6674\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__6683\,
            I => \N__6674\
        );

    \I__961\ : CEMux
    port map (
            O => \N__6682\,
            I => \N__6671\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__6679\,
            I => \N__6668\
        );

    \I__959\ : Span4Mux_h
    port map (
            O => \N__6674\,
            I => \N__6665\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__6671\,
            I => \N__6660\
        );

    \I__957\ : Span4Mux_h
    port map (
            O => \N__6668\,
            I => \N__6660\
        );

    \I__956\ : Odrv4
    port map (
            O => \N__6665\,
            I => \DUT.fifo_rx_inst.rFifoData_awe1\
        );

    \I__955\ : Odrv4
    port map (
            O => \N__6660\,
            I => \DUT.fifo_rx_inst.rFifoData_awe1\
        );

    \I__954\ : InMux
    port map (
            O => \N__6655\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_0\
        );

    \I__953\ : InMux
    port map (
            O => \N__6652\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_1\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__6649\,
            I => \N__6646\
        );

    \I__951\ : InMux
    port map (
            O => \N__6646\,
            I => \N__6643\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__6643\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_3\
        );

    \I__949\ : InMux
    port map (
            O => \N__6640\,
            I => \N__6636\
        );

    \I__948\ : InMux
    port map (
            O => \N__6639\,
            I => \N__6633\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__6636\,
            I => \N__6630\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__6633\,
            I => \DUT.uart_inst0.rx_clk_divider_1_3\
        );

    \I__945\ : Odrv4
    port map (
            O => \N__6630\,
            I => \DUT.uart_inst0.rx_clk_divider_1_3\
        );

    \I__944\ : InMux
    port map (
            O => \N__6625\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_2\
        );

    \I__943\ : CEMux
    port map (
            O => \N__6622\,
            I => \N__6619\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__6619\,
            I => \N__6614\
        );

    \I__941\ : CEMux
    port map (
            O => \N__6618\,
            I => \N__6610\
        );

    \I__940\ : CEMux
    port map (
            O => \N__6617\,
            I => \N__6607\
        );

    \I__939\ : Span4Mux_h
    port map (
            O => \N__6614\,
            I => \N__6604\
        );

    \I__938\ : CEMux
    port map (
            O => \N__6613\,
            I => \N__6601\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__6610\,
            I => \N__6598\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__6607\,
            I => \N__6595\
        );

    \I__935\ : Span4Mux_h
    port map (
            O => \N__6604\,
            I => \N__6591\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__6601\,
            I => \N__6588\
        );

    \I__933\ : Span4Mux_v
    port map (
            O => \N__6598\,
            I => \N__6583\
        );

    \I__932\ : Span4Mux_v
    port map (
            O => \N__6595\,
            I => \N__6583\
        );

    \I__931\ : InMux
    port map (
            O => \N__6594\,
            I => \N__6580\
        );

    \I__930\ : Odrv4
    port map (
            O => \N__6591\,
            I => \DUT.fifo_rx_inst.rFifoData_awe2\
        );

    \I__929\ : Odrv12
    port map (
            O => \N__6588\,
            I => \DUT.fifo_rx_inst.rFifoData_awe2\
        );

    \I__928\ : Odrv4
    port map (
            O => \N__6583\,
            I => \DUT.fifo_rx_inst.rFifoData_awe2\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__6580\,
            I => \DUT.fifo_rx_inst.rFifoData_awe2\
        );

    \I__926\ : InMux
    port map (
            O => \N__6571\,
            I => \N__6567\
        );

    \I__925\ : InMux
    port map (
            O => \N__6570\,
            I => \N__6564\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__6567\,
            I => \DUT.fifo_rx_inst.rFifoDataro_2\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__6564\,
            I => \DUT.fifo_rx_inst.rFifoDataro_2\
        );

    \I__922\ : CEMux
    port map (
            O => \N__6559\,
            I => \N__6556\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__6556\,
            I => \N__6553\
        );

    \I__920\ : Span4Mux_h
    port map (
            O => \N__6553\,
            I => \N__6549\
        );

    \I__919\ : InMux
    port map (
            O => \N__6552\,
            I => \N__6546\
        );

    \I__918\ : Odrv4
    port map (
            O => \N__6549\,
            I => \DUT.fifo_tx_inst.rFifoData_awe1\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__6546\,
            I => \DUT.fifo_tx_inst.rFifoData_awe1\
        );

    \I__916\ : CascadeMux
    port map (
            O => \N__6541\,
            I => \DUT.fifo_tx_inst.rFifoData_awe3_cascade_\
        );

    \I__915\ : InMux
    port map (
            O => \N__6538\,
            I => \N__6535\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__6535\,
            I => \DUT.fifo_tx_inst.un1_i11_i\
        );

    \I__913\ : CascadeMux
    port map (
            O => \N__6532\,
            I => \DUT.fifo_tx_inst.un1_i11_i_cascade_\
        );

    \I__912\ : InMux
    port map (
            O => \N__6529\,
            I => \N__6526\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__6526\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_1\
        );

    \I__910\ : CascadeMux
    port map (
            O => \N__6523\,
            I => \N__6520\
        );

    \I__909\ : InMux
    port map (
            O => \N__6520\,
            I => \N__6517\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__6517\,
            I => \N__6514\
        );

    \I__907\ : Odrv4
    port map (
            O => \N__6514\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_6\
        );

    \I__906\ : InMux
    port map (
            O => \N__6511\,
            I => \N__6508\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__6508\,
            I => \N__6505\
        );

    \I__904\ : Odrv4
    port map (
            O => \N__6505\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_7\
        );

    \I__903\ : CEMux
    port map (
            O => \N__6502\,
            I => \N__6497\
        );

    \I__902\ : InMux
    port map (
            O => \N__6501\,
            I => \N__6494\
        );

    \I__901\ : InMux
    port map (
            O => \N__6500\,
            I => \N__6491\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__6497\,
            I => \DUT.fifo_rx_inst.rFifoData_awe3\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__6494\,
            I => \DUT.fifo_rx_inst.rFifoData_awe3\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__6491\,
            I => \DUT.fifo_rx_inst.rFifoData_awe3\
        );

    \I__897\ : InMux
    port map (
            O => \N__6484\,
            I => \N__6480\
        );

    \I__896\ : InMux
    port map (
            O => \N__6483\,
            I => \N__6477\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__6480\,
            I => \DUT.fifo_rx_inst.rFifoDataro_3\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__6477\,
            I => \DUT.fifo_rx_inst.rFifoDataro_3\
        );

    \I__893\ : InMux
    port map (
            O => \N__6472\,
            I => \N__6469\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__6469\,
            I => \N__6465\
        );

    \I__891\ : InMux
    port map (
            O => \N__6468\,
            I => \N__6462\
        );

    \I__890\ : Span4Mux_s2_v
    port map (
            O => \N__6465\,
            I => \N__6459\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__6462\,
            I => \DUT.uart_inst0.recv_stateZ0Z_4\
        );

    \I__888\ : Odrv4
    port map (
            O => \N__6459\,
            I => \DUT.uart_inst0.recv_stateZ0Z_4\
        );

    \I__887\ : CEMux
    port map (
            O => \N__6454\,
            I => \N__6451\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__6451\,
            I => \N__6447\
        );

    \I__885\ : CEMux
    port map (
            O => \N__6450\,
            I => \N__6444\
        );

    \I__884\ : Span4Mux_h
    port map (
            O => \N__6447\,
            I => \N__6441\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__6444\,
            I => \N__6438\
        );

    \I__882\ : Odrv4
    port map (
            O => \N__6441\,
            I => \fifo_inst.ftdi_output_inst.rFifoState_0_1\
        );

    \I__881\ : Odrv4
    port map (
            O => \N__6438\,
            I => \fifo_inst.ftdi_output_inst.rFifoState_0_1\
        );

    \I__880\ : InMux
    port map (
            O => \N__6433\,
            I => \N__6430\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__6430\,
            I => \N__6427\
        );

    \I__878\ : Odrv12
    port map (
            O => \N__6427\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_0\
        );

    \I__877\ : CascadeMux
    port map (
            O => \N__6424\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_\
        );

    \I__876\ : CascadeMux
    port map (
            O => \N__6421\,
            I => \N__6418\
        );

    \I__875\ : InMux
    port map (
            O => \N__6418\,
            I => \N__6415\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__6415\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_0\
        );

    \I__873\ : InMux
    port map (
            O => \N__6412\,
            I => \N__6409\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__6409\,
            I => \N__6406\
        );

    \I__871\ : Span4Mux_h
    port map (
            O => \N__6406\,
            I => \N__6403\
        );

    \I__870\ : Odrv4
    port map (
            O => \N__6403\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_1\
        );

    \I__869\ : InMux
    port map (
            O => \N__6400\,
            I => \N__6397\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__6397\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_0\
        );

    \I__867\ : InMux
    port map (
            O => \N__6394\,
            I => \N__6391\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__6391\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_1\
        );

    \I__865\ : InMux
    port map (
            O => \N__6388\,
            I => \N__6382\
        );

    \I__864\ : InMux
    port map (
            O => \N__6387\,
            I => \N__6382\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__6382\,
            I => \N__6379\
        );

    \I__862\ : Odrv4
    port map (
            O => \N__6379\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_0\
        );

    \I__861\ : CascadeMux
    port map (
            O => \N__6376\,
            I => \N__6372\
        );

    \I__860\ : CascadeMux
    port map (
            O => \N__6375\,
            I => \N__6369\
        );

    \I__859\ : InMux
    port map (
            O => \N__6372\,
            I => \N__6362\
        );

    \I__858\ : InMux
    port map (
            O => \N__6369\,
            I => \N__6362\
        );

    \I__857\ : InMux
    port map (
            O => \N__6368\,
            I => \N__6354\
        );

    \I__856\ : InMux
    port map (
            O => \N__6367\,
            I => \N__6351\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__6362\,
            I => \N__6348\
        );

    \I__854\ : InMux
    port map (
            O => \N__6361\,
            I => \N__6337\
        );

    \I__853\ : InMux
    port map (
            O => \N__6360\,
            I => \N__6337\
        );

    \I__852\ : InMux
    port map (
            O => \N__6359\,
            I => \N__6337\
        );

    \I__851\ : InMux
    port map (
            O => \N__6358\,
            I => \N__6337\
        );

    \I__850\ : InMux
    port map (
            O => \N__6357\,
            I => \N__6337\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__6354\,
            I => \DUT.uart_inst0.rx_clk_divider_1_i_3\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__6351\,
            I => \DUT.uart_inst0.rx_clk_divider_1_i_3\
        );

    \I__847\ : Odrv4
    port map (
            O => \N__6348\,
            I => \DUT.uart_inst0.rx_clk_divider_1_i_3\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__6337\,
            I => \DUT.uart_inst0.rx_clk_divider_1_i_3\
        );

    \I__845\ : CascadeMux
    port map (
            O => \N__6328\,
            I => \N__6321\
        );

    \I__844\ : CascadeMux
    port map (
            O => \N__6327\,
            I => \N__6318\
        );

    \I__843\ : InMux
    port map (
            O => \N__6326\,
            I => \N__6313\
        );

    \I__842\ : InMux
    port map (
            O => \N__6325\,
            I => \N__6308\
        );

    \I__841\ : InMux
    port map (
            O => \N__6324\,
            I => \N__6308\
        );

    \I__840\ : InMux
    port map (
            O => \N__6321\,
            I => \N__6299\
        );

    \I__839\ : InMux
    port map (
            O => \N__6318\,
            I => \N__6299\
        );

    \I__838\ : InMux
    port map (
            O => \N__6317\,
            I => \N__6299\
        );

    \I__837\ : InMux
    port map (
            O => \N__6316\,
            I => \N__6299\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__6313\,
            I => \DUT.uart_inst0.N_275\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__6308\,
            I => \DUT.uart_inst0.N_275\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__6299\,
            I => \DUT.uart_inst0.N_275\
        );

    \I__833\ : CascadeMux
    port map (
            O => \N__6292\,
            I => \DUT.uart_inst0.N_196_cascade_\
        );

    \I__832\ : CascadeMux
    port map (
            O => \N__6289\,
            I => \DUT.uart_inst0.N_33_cascade_\
        );

    \I__831\ : CEMux
    port map (
            O => \N__6286\,
            I => \N__6283\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__6283\,
            I => \N__6280\
        );

    \I__829\ : Span4Mux_s3_v
    port map (
            O => \N__6280\,
            I => \N__6277\
        );

    \I__828\ : Odrv4
    port map (
            O => \N__6277\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_3_0_c_RNIP8IZ0Z482\
        );

    \I__827\ : InMux
    port map (
            O => \N__6274\,
            I => \N__6271\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__6271\,
            I => \DUT.uart_inst0.rx_bits_remaining_RNO_0Z0Z_1\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__6268\,
            I => \N__6264\
        );

    \I__824\ : InMux
    port map (
            O => \N__6267\,
            I => \N__6261\
        );

    \I__823\ : InMux
    port map (
            O => \N__6264\,
            I => \N__6258\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__6261\,
            I => \DUT.uart_inst0.g0_8_1\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__6258\,
            I => \DUT.uart_inst0.g0_8_1\
        );

    \I__820\ : CEMux
    port map (
            O => \N__6253\,
            I => \N__6250\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__6250\,
            I => \P1A2_c_0_0\
        );

    \I__818\ : CascadeMux
    port map (
            O => \N__6247\,
            I => \DUT.uart_inst0.rx_clk_divider_5_i_a2_11_5_cascade_\
        );

    \I__817\ : InMux
    port map (
            O => \N__6244\,
            I => \N__6241\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__6241\,
            I => \DUT.uart_inst0.N_221\
        );

    \I__815\ : CascadeMux
    port map (
            O => \N__6238\,
            I => \N__6235\
        );

    \I__814\ : InMux
    port map (
            O => \N__6235\,
            I => \N__6232\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__6232\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_0_0_c_RNOZ0\
        );

    \I__812\ : CascadeMux
    port map (
            O => \N__6229\,
            I => \N__6226\
        );

    \I__811\ : InMux
    port map (
            O => \N__6226\,
            I => \N__6223\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__6223\,
            I => \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_0Z0Z_0\
        );

    \I__809\ : InMux
    port map (
            O => \N__6220\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_0\
        );

    \I__808\ : CascadeMux
    port map (
            O => \N__6217\,
            I => \N__6214\
        );

    \I__807\ : InMux
    port map (
            O => \N__6214\,
            I => \N__6211\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__6211\,
            I => \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_1Z0Z_0\
        );

    \I__805\ : InMux
    port map (
            O => \N__6208\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_1\
        );

    \I__804\ : InMux
    port map (
            O => \N__6205\,
            I => \N__6202\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__6202\,
            I => \N__6199\
        );

    \I__802\ : Odrv4
    port map (
            O => \N__6199\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__801\ : CascadeMux
    port map (
            O => \N__6196\,
            I => \N__6193\
        );

    \I__800\ : InMux
    port map (
            O => \N__6193\,
            I => \N__6190\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__6190\,
            I => \DUT.uart_inst0.rx_clk_divider_RNIP8N2BZ0Z_0\
        );

    \I__798\ : InMux
    port map (
            O => \N__6187\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_2\
        );

    \I__797\ : InMux
    port map (
            O => \N__6184\,
            I => \N__6181\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__6181\,
            I => \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_2Z0Z_0\
        );

    \I__795\ : InMux
    port map (
            O => \N__6178\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_3\
        );

    \I__794\ : InMux
    port map (
            O => \N__6175\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_4\
        );

    \I__793\ : CascadeMux
    port map (
            O => \N__6172\,
            I => \DUT.uart_inst0.rx_countdown_3_5_cascade_\
        );

    \I__792\ : InMux
    port map (
            O => \N__6169\,
            I => \N__6166\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__6166\,
            I => \DUT.uart_inst0.g3_4\
        );

    \I__790\ : InMux
    port map (
            O => \N__6163\,
            I => \N__6160\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__6160\,
            I => \DUT.uart_inst0.rx_clk_divider_5_i_a2_1_3\
        );

    \I__788\ : CascadeMux
    port map (
            O => \N__6157\,
            I => \DUT.uart_inst0.N_222_cascade_\
        );

    \I__787\ : CascadeMux
    port map (
            O => \N__6154\,
            I => \DUT.uart_inst0.rx_clk_divider_5_i_a2_11_0_5_cascade_\
        );

    \I__786\ : InMux
    port map (
            O => \N__6151\,
            I => \N__6147\
        );

    \I__785\ : InMux
    port map (
            O => \N__6150\,
            I => \N__6144\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__6147\,
            I => \DUT.uart_inst0.rx_clk_divider_5_i_a2_11_5\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__6144\,
            I => \DUT.uart_inst0.rx_clk_divider_5_i_a2_11_5\
        );

    \I__782\ : InMux
    port map (
            O => \N__6139\,
            I => \N__6136\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__6136\,
            I => \N__6133\
        );

    \I__780\ : Odrv4
    port map (
            O => \N__6133\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_2\
        );

    \I__779\ : InMux
    port map (
            O => \N__6130\,
            I => \N__6127\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__6127\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_3\
        );

    \I__777\ : InMux
    port map (
            O => \N__6124\,
            I => \N__6121\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__6121\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_4\
        );

    \I__775\ : CEMux
    port map (
            O => \N__6118\,
            I => \N__6115\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__6115\,
            I => \N__6110\
        );

    \I__773\ : CEMux
    port map (
            O => \N__6114\,
            I => \N__6107\
        );

    \I__772\ : CEMux
    port map (
            O => \N__6113\,
            I => \N__6104\
        );

    \I__771\ : Span4Mux_h
    port map (
            O => \N__6110\,
            I => \N__6097\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__6107\,
            I => \N__6097\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__6104\,
            I => \N__6094\
        );

    \I__768\ : CEMux
    port map (
            O => \N__6103\,
            I => \N__6091\
        );

    \I__767\ : InMux
    port map (
            O => \N__6102\,
            I => \N__6088\
        );

    \I__766\ : Span4Mux_h
    port map (
            O => \N__6097\,
            I => \N__6085\
        );

    \I__765\ : Sp12to4
    port map (
            O => \N__6094\,
            I => \N__6078\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__6091\,
            I => \N__6078\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__6088\,
            I => \N__6078\
        );

    \I__762\ : Odrv4
    port map (
            O => \N__6085\,
            I => \DUT.fifo_rx_inst.rFifoData_awe0\
        );

    \I__761\ : Odrv12
    port map (
            O => \N__6078\,
            I => \DUT.fifo_rx_inst.rFifoData_awe0\
        );

    \I__760\ : InMux
    port map (
            O => \N__6073\,
            I => \N__6070\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__6070\,
            I => \N__6067\
        );

    \I__758\ : Odrv4
    port map (
            O => \N__6067\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_2\
        );

    \I__757\ : InMux
    port map (
            O => \N__6064\,
            I => \N__6061\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__6061\,
            I => \N__6058\
        );

    \I__755\ : Odrv4
    port map (
            O => \N__6058\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_5\
        );

    \I__754\ : CascadeMux
    port map (
            O => \N__6055\,
            I => \DUT.fifo_rx_inst.N_194_cascade_\
        );

    \I__753\ : InMux
    port map (
            O => \N__6052\,
            I => \N__6049\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__6049\,
            I => \N__6046\
        );

    \I__751\ : Odrv4
    port map (
            O => \N__6046\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_2\
        );

    \I__750\ : InMux
    port map (
            O => \N__6043\,
            I => \N__6040\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__6040\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_2\
        );

    \I__748\ : CascadeMux
    port map (
            O => \N__6037\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2_cascade_\
        );

    \I__747\ : InMux
    port map (
            O => \N__6034\,
            I => \N__6031\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__6031\,
            I => \N__6028\
        );

    \I__745\ : Odrv4
    port map (
            O => \N__6028\,
            I => \DUT.rFifoDatarx_0_2\
        );

    \I__744\ : CascadeMux
    port map (
            O => \N__6025\,
            I => \DUT.rFifoDataror_0_0_cascade_\
        );

    \I__743\ : InMux
    port map (
            O => \N__6022\,
            I => \N__6019\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__6019\,
            I => \DUT.rFifoDataror_1\
        );

    \I__741\ : InMux
    port map (
            O => \N__6016\,
            I => \N__6002\
        );

    \I__740\ : InMux
    port map (
            O => \N__6015\,
            I => \N__6002\
        );

    \I__739\ : InMux
    port map (
            O => \N__6014\,
            I => \N__6002\
        );

    \I__738\ : InMux
    port map (
            O => \N__6013\,
            I => \N__5991\
        );

    \I__737\ : InMux
    port map (
            O => \N__6012\,
            I => \N__5991\
        );

    \I__736\ : InMux
    port map (
            O => \N__6011\,
            I => \N__5991\
        );

    \I__735\ : InMux
    port map (
            O => \N__6010\,
            I => \N__5991\
        );

    \I__734\ : InMux
    port map (
            O => \N__6009\,
            I => \N__5991\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__6002\,
            I => \N__5986\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__5991\,
            I => \N__5986\
        );

    \I__731\ : Odrv4
    port map (
            O => \N__5986\,
            I => \DUT.uart_inst0.N_257\
        );

    \I__730\ : InMux
    port map (
            O => \N__5983\,
            I => \N__5980\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__5980\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_3\
        );

    \I__728\ : InMux
    port map (
            O => \N__5977\,
            I => \N__5974\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__5974\,
            I => \N__5971\
        );

    \I__726\ : Odrv4
    port map (
            O => \N__5971\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_3\
        );

    \I__725\ : CascadeMux
    port map (
            O => \N__5968\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_\
        );

    \I__724\ : InMux
    port map (
            O => \N__5965\,
            I => \N__5962\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__5962\,
            I => \N__5959\
        );

    \I__722\ : Odrv4
    port map (
            O => \N__5959\,
            I => \DUT.rFifoDatarx_3\
        );

    \I__721\ : CascadeMux
    port map (
            O => \N__5956\,
            I => \N__5950\
        );

    \I__720\ : InMux
    port map (
            O => \N__5955\,
            I => \N__5938\
        );

    \I__719\ : InMux
    port map (
            O => \N__5954\,
            I => \N__5933\
        );

    \I__718\ : InMux
    port map (
            O => \N__5953\,
            I => \N__5933\
        );

    \I__717\ : InMux
    port map (
            O => \N__5950\,
            I => \N__5930\
        );

    \I__716\ : InMux
    port map (
            O => \N__5949\,
            I => \N__5925\
        );

    \I__715\ : InMux
    port map (
            O => \N__5948\,
            I => \N__5925\
        );

    \I__714\ : InMux
    port map (
            O => \N__5947\,
            I => \N__5920\
        );

    \I__713\ : InMux
    port map (
            O => \N__5946\,
            I => \N__5920\
        );

    \I__712\ : InMux
    port map (
            O => \N__5945\,
            I => \N__5915\
        );

    \I__711\ : InMux
    port map (
            O => \N__5944\,
            I => \N__5915\
        );

    \I__710\ : InMux
    port map (
            O => \N__5943\,
            I => \N__5908\
        );

    \I__709\ : InMux
    port map (
            O => \N__5942\,
            I => \N__5908\
        );

    \I__708\ : InMux
    port map (
            O => \N__5941\,
            I => \N__5908\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__5938\,
            I => \N__5903\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__5933\,
            I => \N__5903\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__5930\,
            I => \N__5900\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__5925\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__5920\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__5915\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__5908\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__700\ : Odrv4
    port map (
            O => \N__5903\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__699\ : Odrv4
    port map (
            O => \N__5900\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__698\ : CascadeMux
    port map (
            O => \N__5887\,
            I => \N__5882\
        );

    \I__697\ : CascadeMux
    port map (
            O => \N__5886\,
            I => \N__5871\
        );

    \I__696\ : CascadeMux
    port map (
            O => \N__5885\,
            I => \N__5866\
        );

    \I__695\ : InMux
    port map (
            O => \N__5882\,
            I => \N__5862\
        );

    \I__694\ : CascadeMux
    port map (
            O => \N__5881\,
            I => \N__5858\
        );

    \I__693\ : CascadeMux
    port map (
            O => \N__5880\,
            I => \N__5855\
        );

    \I__692\ : CascadeMux
    port map (
            O => \N__5879\,
            I => \N__5848\
        );

    \I__691\ : CascadeMux
    port map (
            O => \N__5878\,
            I => \N__5844\
        );

    \I__690\ : CascadeMux
    port map (
            O => \N__5877\,
            I => \N__5841\
        );

    \I__689\ : CascadeMux
    port map (
            O => \N__5876\,
            I => \N__5838\
        );

    \I__688\ : InMux
    port map (
            O => \N__5875\,
            I => \N__5831\
        );

    \I__687\ : InMux
    port map (
            O => \N__5874\,
            I => \N__5831\
        );

    \I__686\ : InMux
    port map (
            O => \N__5871\,
            I => \N__5831\
        );

    \I__685\ : InMux
    port map (
            O => \N__5870\,
            I => \N__5822\
        );

    \I__684\ : InMux
    port map (
            O => \N__5869\,
            I => \N__5822\
        );

    \I__683\ : InMux
    port map (
            O => \N__5866\,
            I => \N__5822\
        );

    \I__682\ : InMux
    port map (
            O => \N__5865\,
            I => \N__5822\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__5862\,
            I => \N__5819\
        );

    \I__680\ : InMux
    port map (
            O => \N__5861\,
            I => \N__5814\
        );

    \I__679\ : InMux
    port map (
            O => \N__5858\,
            I => \N__5814\
        );

    \I__678\ : InMux
    port map (
            O => \N__5855\,
            I => \N__5811\
        );

    \I__677\ : InMux
    port map (
            O => \N__5854\,
            I => \N__5800\
        );

    \I__676\ : InMux
    port map (
            O => \N__5853\,
            I => \N__5800\
        );

    \I__675\ : InMux
    port map (
            O => \N__5852\,
            I => \N__5800\
        );

    \I__674\ : InMux
    port map (
            O => \N__5851\,
            I => \N__5800\
        );

    \I__673\ : InMux
    port map (
            O => \N__5848\,
            I => \N__5800\
        );

    \I__672\ : InMux
    port map (
            O => \N__5847\,
            I => \N__5793\
        );

    \I__671\ : InMux
    port map (
            O => \N__5844\,
            I => \N__5793\
        );

    \I__670\ : InMux
    port map (
            O => \N__5841\,
            I => \N__5793\
        );

    \I__669\ : InMux
    port map (
            O => \N__5838\,
            I => \N__5790\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__5831\,
            I => \N__5787\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__5822\,
            I => \N__5784\
        );

    \I__666\ : Odrv4
    port map (
            O => \N__5819\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__5814\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__5811\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__5800\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__5793\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__5790\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__660\ : Odrv4
    port map (
            O => \N__5787\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__659\ : Odrv4
    port map (
            O => \N__5784\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__658\ : InMux
    port map (
            O => \N__5767\,
            I => \N__5764\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__5764\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4\
        );

    \I__656\ : InMux
    port map (
            O => \N__5761\,
            I => \N__5758\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__5758\,
            I => \wRxFifoData_3\
        );

    \I__654\ : InMux
    port map (
            O => \N__5755\,
            I => \N__5752\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__5752\,
            I => \N__5749\
        );

    \I__652\ : Span4Mux_h
    port map (
            O => \N__5749\,
            I => \N__5746\
        );

    \I__651\ : Odrv4
    port map (
            O => \N__5746\,
            I => \DUT.rFifoDatarx_0_5\
        );

    \I__650\ : CascadeMux
    port map (
            O => \N__5743\,
            I => \N__5740\
        );

    \I__649\ : InMux
    port map (
            O => \N__5740\,
            I => \N__5737\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__5737\,
            I => \wRxFifoData_5\
        );

    \I__647\ : InMux
    port map (
            O => \N__5734\,
            I => \N__5731\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__5731\,
            I => \DUT.rFifoDatarx_0_7\
        );

    \I__645\ : CascadeMux
    port map (
            O => \N__5728\,
            I => \N__5725\
        );

    \I__644\ : InMux
    port map (
            O => \N__5725\,
            I => \N__5722\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__5722\,
            I => \wRxFifoData_7\
        );

    \I__642\ : CEMux
    port map (
            O => \N__5719\,
            I => \N__5715\
        );

    \I__641\ : CEMux
    port map (
            O => \N__5718\,
            I => \N__5712\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__5715\,
            I => \N__5709\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__5712\,
            I => \N__5706\
        );

    \I__638\ : Odrv4
    port map (
            O => \N__5709\,
            I => \un1_oRxFlag_0_i_0\
        );

    \I__637\ : Odrv4
    port map (
            O => \N__5706\,
            I => \un1_oRxFlag_0_i_0\
        );

    \I__636\ : CascadeMux
    port map (
            O => \N__5701\,
            I => \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1_cascade_\
        );

    \I__635\ : InMux
    port map (
            O => \N__5698\,
            I => \N__5695\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__5695\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_1\
        );

    \I__633\ : InMux
    port map (
            O => \N__5692\,
            I => \N__5689\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__5689\,
            I => \N__5686\
        );

    \I__631\ : Odrv4
    port map (
            O => \N__5686\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1\
        );

    \I__630\ : InMux
    port map (
            O => \N__5683\,
            I => \N__5680\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__5680\,
            I => \DUT.rFifoDatarx_0_1\
        );

    \I__628\ : InMux
    port map (
            O => \N__5677\,
            I => \N__5674\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__5674\,
            I => \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1\
        );

    \I__626\ : InMux
    port map (
            O => \N__5671\,
            I => \N__5665\
        );

    \I__625\ : InMux
    port map (
            O => \N__5670\,
            I => \N__5665\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__5665\,
            I => \N__5658\
        );

    \I__623\ : InMux
    port map (
            O => \N__5664\,
            I => \N__5653\
        );

    \I__622\ : InMux
    port map (
            O => \N__5663\,
            I => \N__5653\
        );

    \I__621\ : InMux
    port map (
            O => \N__5662\,
            I => \N__5650\
        );

    \I__620\ : InMux
    port map (
            O => \N__5661\,
            I => \N__5647\
        );

    \I__619\ : Span4Mux_v
    port map (
            O => \N__5658\,
            I => \N__5642\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__5653\,
            I => \N__5642\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__5650\,
            I => \DUT.wRcvd\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__5647\,
            I => \DUT.wRcvd\
        );

    \I__615\ : Odrv4
    port map (
            O => \N__5642\,
            I => \DUT.wRcvd\
        );

    \I__614\ : InMux
    port map (
            O => \N__5635\,
            I => \N__5629\
        );

    \I__613\ : InMux
    port map (
            O => \N__5634\,
            I => \N__5629\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__5629\,
            I => \N__5625\
        );

    \I__611\ : InMux
    port map (
            O => \N__5628\,
            I => \N__5618\
        );

    \I__610\ : Span4Mux_v
    port map (
            O => \N__5625\,
            I => \N__5615\
        );

    \I__609\ : InMux
    port map (
            O => \N__5624\,
            I => \N__5610\
        );

    \I__608\ : InMux
    port map (
            O => \N__5623\,
            I => \N__5610\
        );

    \I__607\ : InMux
    port map (
            O => \N__5622\,
            I => \N__5605\
        );

    \I__606\ : InMux
    port map (
            O => \N__5621\,
            I => \N__5605\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__5618\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\
        );

    \I__604\ : Odrv4
    port map (
            O => \N__5615\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__5610\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__5605\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\
        );

    \I__601\ : CascadeMux
    port map (
            O => \N__5596\,
            I => \N__5592\
        );

    \I__600\ : InMux
    port map (
            O => \N__5595\,
            I => \N__5586\
        );

    \I__599\ : InMux
    port map (
            O => \N__5592\,
            I => \N__5583\
        );

    \I__598\ : InMux
    port map (
            O => \N__5591\,
            I => \N__5580\
        );

    \I__597\ : InMux
    port map (
            O => \N__5590\,
            I => \N__5575\
        );

    \I__596\ : InMux
    port map (
            O => \N__5589\,
            I => \N__5575\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__5586\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_1\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__5583\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_1\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__5580\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_1\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__5575\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_1\
        );

    \I__591\ : InMux
    port map (
            O => \N__5566\,
            I => \N__5556\
        );

    \I__590\ : InMux
    port map (
            O => \N__5565\,
            I => \N__5556\
        );

    \I__589\ : InMux
    port map (
            O => \N__5564\,
            I => \N__5556\
        );

    \I__588\ : CascadeMux
    port map (
            O => \N__5563\,
            I => \N__5552\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__5556\,
            I => \N__5549\
        );

    \I__586\ : CascadeMux
    port map (
            O => \N__5555\,
            I => \N__5546\
        );

    \I__585\ : InMux
    port map (
            O => \N__5552\,
            I => \N__5543\
        );

    \I__584\ : Span4Mux_v
    port map (
            O => \N__5549\,
            I => \N__5540\
        );

    \I__583\ : InMux
    port map (
            O => \N__5546\,
            I => \N__5537\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__5543\,
            I => \DUT.fifo_rx_inst.N_148\
        );

    \I__581\ : Odrv4
    port map (
            O => \N__5540\,
            I => \DUT.fifo_rx_inst.N_148\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__5537\,
            I => \DUT.fifo_rx_inst.N_148\
        );

    \I__579\ : InMux
    port map (
            O => \N__5530\,
            I => \N__5527\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__5527\,
            I => \N__5524\
        );

    \I__577\ : Span4Mux_v
    port map (
            O => \N__5524\,
            I => \N__5521\
        );

    \I__576\ : Sp12to4
    port map (
            O => \N__5521\,
            I => \N__5518\
        );

    \I__575\ : Span12Mux_h
    port map (
            O => \N__5518\,
            I => \N__5515\
        );

    \I__574\ : Span12Mux_v
    port map (
            O => \N__5515\,
            I => \N__5512\
        );

    \I__573\ : Odrv12
    port map (
            O => \N__5512\,
            I => \ioFifoData_in_7\
        );

    \I__572\ : InMux
    port map (
            O => \N__5509\,
            I => \N__5506\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__5506\,
            I => \N__5503\
        );

    \I__570\ : Span4Mux_h
    port map (
            O => \N__5503\,
            I => \N__5500\
        );

    \I__569\ : Span4Mux_v
    port map (
            O => \N__5500\,
            I => \N__5497\
        );

    \I__568\ : Odrv4
    port map (
            O => \N__5497\,
            I => \ioFifoData_in_1\
        );

    \I__567\ : InMux
    port map (
            O => \N__5494\,
            I => \N__5491\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__5491\,
            I => \N__5488\
        );

    \I__565\ : Span4Mux_h
    port map (
            O => \N__5488\,
            I => \N__5485\
        );

    \I__564\ : Span4Mux_h
    port map (
            O => \N__5485\,
            I => \N__5482\
        );

    \I__563\ : Span4Mux_v
    port map (
            O => \N__5482\,
            I => \N__5479\
        );

    \I__562\ : Odrv4
    port map (
            O => \N__5479\,
            I => \ioFifoData_in_3\
        );

    \I__561\ : InMux
    port map (
            O => \N__5476\,
            I => \N__5473\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__5473\,
            I => \N__5470\
        );

    \I__559\ : Span4Mux_v
    port map (
            O => \N__5470\,
            I => \N__5467\
        );

    \I__558\ : Span4Mux_h
    port map (
            O => \N__5467\,
            I => \N__5464\
        );

    \I__557\ : Odrv4
    port map (
            O => \N__5464\,
            I => \ioFifoData_in_5\
        );

    \I__556\ : InMux
    port map (
            O => \N__5461\,
            I => \N__5458\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__5458\,
            I => \N__5455\
        );

    \I__554\ : Span4Mux_v
    port map (
            O => \N__5455\,
            I => \N__5452\
        );

    \I__553\ : Span4Mux_h
    port map (
            O => \N__5452\,
            I => \N__5449\
        );

    \I__552\ : Span4Mux_h
    port map (
            O => \N__5449\,
            I => \N__5446\
        );

    \I__551\ : Odrv4
    port map (
            O => \N__5446\,
            I => \ioFifoData_in_2\
        );

    \I__550\ : CascadeMux
    port map (
            O => \N__5443\,
            I => \N__5440\
        );

    \I__549\ : InMux
    port map (
            O => \N__5440\,
            I => \N__5437\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__5437\,
            I => \wRxFifoData_1\
        );

    \I__547\ : CascadeMux
    port map (
            O => \N__5434\,
            I => \N__5431\
        );

    \I__546\ : InMux
    port map (
            O => \N__5431\,
            I => \N__5428\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__5428\,
            I => \N__5425\
        );

    \I__544\ : Odrv4
    port map (
            O => \N__5425\,
            I => \wRxFifoData_2\
        );

    \I__543\ : CascadeMux
    port map (
            O => \N__5422\,
            I => \DUT.uart_inst0.g0_0_5_cascade_\
        );

    \I__542\ : CascadeMux
    port map (
            O => \N__5419\,
            I => \DUT.uart_inst0.g0_6_cascade_\
        );

    \I__541\ : InMux
    port map (
            O => \N__5416\,
            I => \N__5413\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__5413\,
            I => \N__5410\
        );

    \I__539\ : Odrv4
    port map (
            O => \N__5410\,
            I => \DUT.uart_inst0.g0_1_0\
        );

    \I__538\ : CascadeMux
    port map (
            O => \N__5407\,
            I => \DUT.uart_inst0.g3_0_cascade_\
        );

    \I__537\ : InMux
    port map (
            O => \N__5404\,
            I => \N__5401\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__5401\,
            I => \DUT.uart_inst0.g0_0_4\
        );

    \I__535\ : InMux
    port map (
            O => \N__5398\,
            I => \N__5395\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__5395\,
            I => \N__5392\
        );

    \I__533\ : Odrv4
    port map (
            O => \N__5392\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_4\
        );

    \I__532\ : IoInMux
    port map (
            O => \N__5389\,
            I => \N__5386\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__5386\,
            I => \wPllLocked_i\
        );

    \I__530\ : CascadeMux
    port map (
            O => \N__5383\,
            I => \DUT.uart_inst0.N_275_cascade_\
        );

    \I__529\ : CascadeMux
    port map (
            O => \N__5380\,
            I => \DUT.fifo_rx_inst.rReadPtr_RNIDU4H2Z0Z_0_cascade_\
        );

    \I__528\ : InMux
    port map (
            O => \N__5377\,
            I => \N__5374\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__5374\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_6\
        );

    \I__526\ : InMux
    port map (
            O => \N__5371\,
            I => \N__5368\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__5368\,
            I => \N__5365\
        );

    \I__524\ : Odrv4
    port map (
            O => \N__5365\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6\
        );

    \I__523\ : InMux
    port map (
            O => \N__5362\,
            I => \N__5359\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__5359\,
            I => \DUT.fifo_rx_inst.rReadPtr_RNIDU4H2Z0Z_0\
        );

    \I__521\ : CascadeMux
    port map (
            O => \N__5356\,
            I => \N__5353\
        );

    \I__520\ : InMux
    port map (
            O => \N__5353\,
            I => \N__5350\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__5350\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_4\
        );

    \I__518\ : InMux
    port map (
            O => \N__5347\,
            I => \N__5344\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__5344\,
            I => \N__5341\
        );

    \I__516\ : Odrv4
    port map (
            O => \N__5341\,
            I => \DUT.rFifoDatarx_0_4\
        );

    \I__515\ : InMux
    port map (
            O => \N__5338\,
            I => \N__5335\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__5335\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_5\
        );

    \I__513\ : CascadeMux
    port map (
            O => \N__5332\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_\
        );

    \I__512\ : InMux
    port map (
            O => \N__5329\,
            I => \N__5326\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__5326\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_5\
        );

    \I__510\ : InMux
    port map (
            O => \N__5323\,
            I => \N__5320\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__5320\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_6\
        );

    \I__508\ : InMux
    port map (
            O => \N__5317\,
            I => \N__5313\
        );

    \I__507\ : InMux
    port map (
            O => \N__5316\,
            I => \N__5310\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__5313\,
            I => \N__5305\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__5310\,
            I => \N__5305\
        );

    \I__504\ : Odrv4
    port map (
            O => \N__5305\,
            I => \DUT.fifo_rx_inst.rFifoDataro_0\
        );

    \I__503\ : InMux
    port map (
            O => \N__5302\,
            I => \N__5298\
        );

    \I__502\ : InMux
    port map (
            O => \N__5301\,
            I => \N__5295\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__5298\,
            I => \DUT.fifo_rx_inst.rFifoDataro_1\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__5295\,
            I => \DUT.fifo_rx_inst.rFifoDataro_1\
        );

    \I__499\ : InMux
    port map (
            O => \N__5290\,
            I => \N__5287\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__5287\,
            I => \N__5284\
        );

    \I__497\ : Odrv4
    port map (
            O => \N__5284\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_0\
        );

    \I__496\ : InMux
    port map (
            O => \N__5281\,
            I => \N__5278\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__5278\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_6\
        );

    \I__494\ : InMux
    port map (
            O => \N__5275\,
            I => \N__5272\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__5272\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_7\
        );

    \I__492\ : InMux
    port map (
            O => \N__5269\,
            I => \N__5266\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__5266\,
            I => \N__5263\
        );

    \I__490\ : Sp12to4
    port map (
            O => \N__5263\,
            I => \N__5260\
        );

    \I__489\ : Odrv12
    port map (
            O => \N__5260\,
            I => \ioFifoData_in_0\
        );

    \I__488\ : InMux
    port map (
            O => \N__5257\,
            I => \N__5254\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__5254\,
            I => \N__5251\
        );

    \I__486\ : Span4Mux_h
    port map (
            O => \N__5251\,
            I => \N__5248\
        );

    \I__485\ : Span4Mux_h
    port map (
            O => \N__5248\,
            I => \N__5245\
        );

    \I__484\ : Span4Mux_v
    port map (
            O => \N__5245\,
            I => \N__5242\
        );

    \I__483\ : Odrv4
    port map (
            O => \N__5242\,
            I => \ioFifoData_in_4\
        );

    \I__482\ : CascadeMux
    port map (
            O => \N__5239\,
            I => \N__5236\
        );

    \I__481\ : InMux
    port map (
            O => \N__5236\,
            I => \N__5233\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__5233\,
            I => \wRxFifoData_0\
        );

    \I__479\ : InMux
    port map (
            O => \N__5230\,
            I => \N__5227\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__5227\,
            I => \DUT.rFifoDatarx_0\
        );

    \I__477\ : CascadeMux
    port map (
            O => \N__5224\,
            I => \N__5221\
        );

    \I__476\ : InMux
    port map (
            O => \N__5221\,
            I => \N__5218\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__5218\,
            I => \wRxFifoData_4\
        );

    \I__474\ : CascadeMux
    port map (
            O => \N__5215\,
            I => \N__5212\
        );

    \I__473\ : InMux
    port map (
            O => \N__5212\,
            I => \N__5209\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__5209\,
            I => \wRxFifoData_6\
        );

    \I__471\ : InMux
    port map (
            O => \N__5206\,
            I => \N__5203\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__5203\,
            I => \DUT.rFifoDatarx_6\
        );

    \I__469\ : InMux
    port map (
            O => \N__5200\,
            I => \N__5197\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__5197\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_7\
        );

    \I__467\ : CascadeMux
    port map (
            O => \N__5194\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7_cascade_\
        );

    \I__466\ : InMux
    port map (
            O => \N__5191\,
            I => \N__5188\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__5188\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_7\
        );

    \I__464\ : InMux
    port map (
            O => \N__5185\,
            I => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0\
        );

    \I__463\ : InMux
    port map (
            O => \N__5182\,
            I => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1\
        );

    \I__462\ : CascadeMux
    port map (
            O => \N__5179\,
            I => \un1_oRxFlag_0_i_cascade_\
        );

    \I__461\ : InMux
    port map (
            O => \N__5176\,
            I => \N__5173\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__5173\,
            I => \DUT.fifo_rx_inst.rFifoCount_RNITA8H2Z0Z_1\
        );

    \I__459\ : CascadeMux
    port map (
            O => \N__5170\,
            I => \rFifoCount_RNIHH0D1_0_cascade_\
        );

    \I__458\ : InMux
    port map (
            O => \N__5167\,
            I => \N__5164\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__5164\,
            I => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0\
        );

    \I__456\ : InMux
    port map (
            O => \N__5161\,
            I => \N__5158\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__5158\,
            I => \N__5155\
        );

    \I__454\ : Span4Mux_v
    port map (
            O => \N__5155\,
            I => \N__5152\
        );

    \I__453\ : Sp12to4
    port map (
            O => \N__5152\,
            I => \N__5149\
        );

    \I__452\ : Span12Mux_h
    port map (
            O => \N__5149\,
            I => \N__5146\
        );

    \I__451\ : Span12Mux_v
    port map (
            O => \N__5146\,
            I => \N__5143\
        );

    \I__450\ : Odrv12
    port map (
            O => \N__5143\,
            I => \ioFifoData_in_6\
        );

    \I__449\ : CascadeMux
    port map (
            O => \N__5140\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_\
        );

    \I__448\ : CascadeMux
    port map (
            O => \N__5137\,
            I => \N__5134\
        );

    \I__447\ : InMux
    port map (
            O => \N__5134\,
            I => \N__5131\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__5131\,
            I => \N__5128\
        );

    \I__445\ : Odrv4
    port map (
            O => \N__5128\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_0\
        );

    \I__444\ : InMux
    port map (
            O => \N__5125\,
            I => \N__5122\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__5122\,
            I => \N__5119\
        );

    \I__442\ : Odrv4
    port map (
            O => \N__5119\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_1\
        );

    \I__441\ : InMux
    port map (
            O => \N__5116\,
            I => \N__5113\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__5113\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_1\
        );

    \I__439\ : InMux
    port map (
            O => \N__5110\,
            I => \N__5107\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__5107\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_0\
        );

    \I__437\ : InMux
    port map (
            O => \N__5104\,
            I => \N__5101\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__5101\,
            I => \N__5098\
        );

    \I__435\ : Odrv4
    port map (
            O => \N__5098\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_0\
        );

    \I__434\ : InMux
    port map (
            O => \N__5095\,
            I => \N__5092\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__5092\,
            I => \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO\
        );

    \I__432\ : IoInMux
    port map (
            O => \N__5089\,
            I => \N__5086\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__5086\,
            I => \N__5083\
        );

    \I__430\ : Span12Mux_s9_v
    port map (
            O => \N__5083\,
            I => \N__5080\
        );

    \I__429\ : Span12Mux_v
    port map (
            O => \N__5080\,
            I => \N__5077\
        );

    \I__428\ : Odrv12
    port map (
            O => \N__5077\,
            I => \BTN_N_c\
        );

    \IN_MUX_bfv_21_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_9_0_\
        );

    \IN_MUX_bfv_21_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DUT.uart_inst0.tx_clk_divider_cry_7\,
            carryinitout => \bfn_21_10_0_\
        );

    \IN_MUX_bfv_14_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_3_0_\
        );

    \IN_MUX_bfv_15_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_1_0_\
        );

    \IN_MUX_bfv_15_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DUT.uart_inst0.rx_clk_divider_1_cry_7\,
            carryinitout => \bfn_15_2_0_\
        );

    \IN_MUX_bfv_15_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DUT.uart_inst0.rx_clk_divider_1_cry_15\,
            carryinitout => \bfn_15_3_0_\
        );

    \IN_MUX_bfv_16_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_11_0_\
        );

    \IN_MUX_bfv_12_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_4_0_\
        );

    \wPllLocked_i_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5389\,
            GLOBALBUFFEROUTPUT => \wPllLocked_i_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \top_pll_inst.top_pll_inst_RNISDA2\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__10639\,
            GLOBALBUFFEROUTPUT => \wPllLocked_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5095\,
            lcout => \wPllLocked\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7330\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12807\,
            ce => \N__10080\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7372\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12801\,
            ce => \N__7414\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7582\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12793\,
            ce => \N__10071\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_0_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6102\,
            in2 => \_gnd_net_\,
            in3 => \N__5317\,
            lcout => \DUT.fifo_rx_inst.rFifoDataro_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12788\,
            ce => 'H',
            sr => \N__11116\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7591\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12782\,
            ce => \N__7412\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7241\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12794\,
            ce => \N__6697\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_1_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5302\,
            in2 => \_gnd_net_\,
            in3 => \N__6689\,
            lcout => \DUT.fifo_rx_inst.rFifoDataro_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12789\,
            ce => 'H',
            sr => \N__11117\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101000111"
        )
    port map (
            in0 => \N__5110\,
            in1 => \N__5954\,
            in2 => \N__5137\,
            in3 => \N__5874\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI5EJ22_0_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__5875\,
            in1 => \N__5290\,
            in2 => \N__5140\,
            in3 => \N__5104\,
            lcout => \DUT.rFifoDatarx_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7192\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12783\,
            ce => \N__6113\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__5953\,
            in1 => \N__5125\,
            in2 => \N__5886\,
            in3 => \N__5116\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7246\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12783\,
            ce => \N__6113\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8461\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12778\,
            ce => \N__6690\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7024\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12778\,
            ce => \N__6690\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7194\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12778\,
            ce => \N__6690\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7068\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12778\,
            ce => \N__6690\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7198\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12775\,
            ce => \N__6618\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5167\,
            in2 => \N__10417\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_4_0_\,
            carryout => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_1_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5176\,
            in2 => \N__5596\,
            in3 => \N__5185\,
            lcout => \DUT.fifo_rx_inst.rFifoCountZ0Z_1\,
            ltout => OPEN,
            carryin => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0\,
            carryout => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1\,
            clk => \N__12800\,
            ce => 'H',
            sr => \N__11124\
        );

    \DUT.fifo_rx_inst.rFifoCount_2_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011011011001001"
        )
    port map (
            in0 => \N__5662\,
            in1 => \N__5628\,
            in2 => \N__5563\,
            in3 => \N__5182\,
            lcout => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12800\,
            ce => 'H',
            sr => \N__11124\
        );

    \DUT.uart_inst0.un1_oRxFlag_0_i_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10322\,
            in2 => \_gnd_net_\,
            in3 => \N__10233\,
            lcout => OPEN,
            ltout => \un1_oRxFlag_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rTxByte_esr_ctle_7_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__11146\,
            in1 => \_gnd_net_\,
            in2 => \N__5179\,
            in3 => \_gnd_net_\,
            lcout => \un1_oRxFlag_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNITA8H2_1_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__5664\,
            in1 => \_gnd_net_\,
            in2 => \N__5555\,
            in3 => \N__5595\,
            lcout => \DUT.fifo_rx_inst.rFifoCount_RNITA8H2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__10404\,
            in1 => \N__5591\,
            in2 => \_gnd_net_\,
            in3 => \N__5622\,
            lcout => \rFifoCount_RNIHH0D1_0\,
            ltout => \rFifoCount_RNIHH0D1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110011"
        )
    port map (
            in0 => \N__10412\,
            in1 => \N__10451\,
            in2 => \N__5170\,
            in3 => \N__10428\,
            lcout => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNIDQ741_2_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110011001"
        )
    port map (
            in0 => \N__10450\,
            in1 => \N__5663\,
            in2 => \_gnd_net_\,
            in3 => \N__5621\,
            lcout => \DUT.fifo_rx_inst.N_206\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rRxData_esr_6_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5161\,
            lcout => \wRxFifoData_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12787\,
            ce => \N__6454\,
            sr => \N__11115\
        );

    \fifo_inst.ftdi_output_inst.rRxData_esr_0_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5269\,
            lcout => \wRxFifoData_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12787\,
            ce => \N__6454\,
            sr => \N__11115\
        );

    \fifo_inst.ftdi_output_inst.rRxData_esr_4_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5257\,
            lcout => \wRxFifoData_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12787\,
            ce => \N__6454\,
            sr => \N__11115\
        );

    \rTxByte_esr_0_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__6014\,
            in1 => \N__10342\,
            in2 => \N__5239\,
            in3 => \N__5230\,
            lcout => \rTxByteZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12781\,
            ce => \N__5718\,
            sr => \N__11112\
        );

    \rTxByte_esr_4_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__10341\,
            in1 => \N__6015\,
            in2 => \N__5224\,
            in3 => \N__5347\,
            lcout => \rTxByteZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12781\,
            ce => \N__5718\,
            sr => \N__11112\
        );

    \rTxByte_esr_6_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__6016\,
            in1 => \N__5206\,
            in2 => \N__5215\,
            in3 => \N__10343\,
            lcout => \rTxByteZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12781\,
            ce => \N__5718\,
            sr => \N__11112\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIT6K22_6_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__5869\,
            in1 => \N__5281\,
            in2 => \N__6523\,
            in3 => \N__5371\,
            lcout => \DUT.rFifoDatarx_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__5955\,
            in1 => \N__5200\,
            in2 => \N__5885\,
            in3 => \N__5191\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI1BK22_7_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__5275\,
            in1 => \N__6511\,
            in2 => \N__5194\,
            in3 => \N__5870\,
            lcout => \DUT.rFifoDatarx_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7022\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12777\,
            ce => \N__6103\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_0_RNI0AQO1_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110101"
        )
    port map (
            in0 => \N__5316\,
            in1 => \N__5301\,
            in2 => \N__5956\,
            in3 => \N__5865\,
            lcout => \DUT.rFifoDataror_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7193\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12774\,
            ce => \N__6502\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7245\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12774\,
            ce => \N__6502\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8449\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12774\,
            ce => \N__6502\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8510\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12774\,
            ce => \N__6502\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7151\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12774\,
            ce => \N__6502\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7106\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12774\,
            ce => \N__6502\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7061\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12774\,
            ce => \N__6502\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7023\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12774\,
            ce => \N__6502\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rReadPtr_RNIDU4H2_0_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110001111"
        )
    port map (
            in0 => \N__5853\,
            in1 => \N__5943\,
            in2 => \N__12440\,
            in3 => \N__5564\,
            lcout => \DUT.fifo_rx_inst.rReadPtr_RNIDU4H2Z0Z_0\,
            ltout => \DUT.fifo_rx_inst.rReadPtr_RNIDU4H2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rReadPtr_1_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100100001100"
        )
    port map (
            in0 => \N__5566\,
            in1 => \N__5854\,
            in2 => \N__5380\,
            in3 => \N__5949\,
            lcout => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12772\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__5941\,
            in1 => \N__5377\,
            in2 => \N__5876\,
            in3 => \N__5323\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rReadPtr_0_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__5948\,
            in1 => \N__5362\,
            in2 => \_gnd_net_\,
            in3 => \N__5565\,
            lcout => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12772\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNILUJ22_4_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__5398\,
            in1 => \N__5852\,
            in2 => \N__5356\,
            in3 => \N__5767\,
            lcout => \DUT.rFifoDatarx_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111110101"
        )
    port map (
            in0 => \N__5329\,
            in1 => \N__6721\,
            in2 => \N__5879\,
            in3 => \N__5942\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIP2K22_5_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__5338\,
            in1 => \N__6064\,
            in2 => \N__5332\,
            in3 => \N__5851\,
            lcout => \DUT.rFifoDatarx_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7113\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12770\,
            ce => \N__6118\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7069\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12770\,
            ce => \N__6118\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8514\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12769\,
            ce => \N__6622\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7159\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12769\,
            ce => \N__6622\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.wPllLocked_i_LC_12_30_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12439\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \wPllLocked_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIHF7P_0_3_LC_13_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6640\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_2_0_LC_13_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6328\,
            in3 => \N__6361\,
            lcout => \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_0_0_LC_13_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6358\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6316\,
            lcout => \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_0_LC_13_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6327\,
            in3 => \N__6360\,
            lcout => \DUT.uart_inst0.rx_clk_divider_RNIP8N2BZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNI8PF9A_0_LC_13_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8220\,
            in1 => \N__6163\,
            in2 => \N__8260\,
            in3 => \N__6150\,
            lcout => \DUT.uart_inst0.N_275\,
            ltout => \DUT.uart_inst0.N_275_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_0_0_c_RNO_LC_13_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5383\,
            in3 => \N__6357\,
            lcout => \DUT.uart_inst0.rx_countdown_3_cry_0_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_1_0_LC_13_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6359\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6317\,
            lcout => \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_0_LC_13_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111011101"
        )
    port map (
            in0 => \N__12421\,
            in1 => \N__5661\,
            in2 => \N__9856\,
            in3 => \N__8279\,
            lcout => \DUT.uart_inst0.g0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_1_2_LC_13_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9640\,
            in1 => \N__9429\,
            in2 => \N__9504\,
            in3 => \N__9716\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g0_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_2_LC_13_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110011001100"
        )
    port map (
            in0 => \N__8728\,
            in1 => \N__8702\,
            in2 => \N__5422\,
            in3 => \N__5404\,
            lcout => \DUT.uart_inst0.rx_bits_remainingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_1_6_LC_13_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9639\,
            in1 => \N__9428\,
            in2 => \N__9503\,
            in3 => \N__9715\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_6_LC_13_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__9560\,
            in1 => \N__9784\,
            in2 => \N__5419\,
            in3 => \N__8050\,
            lcout => \DUT.wRcvd\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_1_0_LC_13_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6472\,
            in2 => \_gnd_net_\,
            in3 => \N__8032\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_0_LC_13_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__9561\,
            in1 => \N__5416\,
            in2 => \N__5407\,
            in3 => \N__6169\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12814\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_0_2_LC_13_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__8308\,
            in1 => \N__9559\,
            in2 => \N__10626\,
            in3 => \N__8031\,
            lcout => \DUT.uart_inst0.g0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_13_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7290\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12808\,
            ce => \N__10079\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNISS2R41_2_LC_13_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__8524\,
            in1 => \N__8027\,
            in2 => \N__9499\,
            in3 => \N__9416\,
            lcout => \DUT.uart_inst0.g0_8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rRxRead_esr_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__5624\,
            in1 => \N__10408\,
            in2 => \_gnd_net_\,
            in3 => \N__5590\,
            lcout => \rRxReadZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12802\,
            ce => \N__6253\,
            sr => \N__11125\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNIIL8L1_0_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110111"
        )
    port map (
            in0 => \N__5589\,
            in1 => \N__10452\,
            in2 => \N__10413\,
            in3 => \N__5623\,
            lcout => \DUT.fifo_rx_inst.N_148\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rRxData_esr_7_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5530\,
            lcout => \wRxFifoData_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12795\,
            ce => \N__6450\,
            sr => \N__11123\
        );

    \fifo_inst.ftdi_output_inst.rRxData_esr_1_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5509\,
            lcout => \wRxFifoData_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12795\,
            ce => \N__6450\,
            sr => \N__11123\
        );

    \fifo_inst.ftdi_output_inst.rRxData_esr_3_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5494\,
            lcout => \wRxFifoData_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12795\,
            ce => \N__6450\,
            sr => \N__11123\
        );

    \fifo_inst.ftdi_output_inst.rRxData_esr_5_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5476\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \wRxFifoData_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12795\,
            ce => \N__6450\,
            sr => \N__11123\
        );

    \fifo_inst.ftdi_output_inst.rRxData_esr_2_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5461\,
            lcout => \wRxFifoData_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12795\,
            ce => \N__6450\,
            sr => \N__11123\
        );

    \rTxByte_esr_1_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__10334\,
            in1 => \N__6009\,
            in2 => \N__5443\,
            in3 => \N__5683\,
            lcout => \rTxByteZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12790\,
            ce => \N__5719\,
            sr => \N__11118\
        );

    \rTxByte_esr_2_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__6010\,
            in1 => \N__10336\,
            in2 => \N__5434\,
            in3 => \N__6034\,
            lcout => \rTxByteZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12790\,
            ce => \N__5719\,
            sr => \N__11118\
        );

    \rTxByte_esr_3_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__6011\,
            in1 => \N__5761\,
            in2 => \N__10347\,
            in3 => \N__5965\,
            lcout => \rTxByteZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12790\,
            ce => \N__5719\,
            sr => \N__11118\
        );

    \rTxByte_esr_5_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__10335\,
            in1 => \N__5755\,
            in2 => \N__5743\,
            in3 => \N__6012\,
            lcout => \rTxByteZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12790\,
            ce => \N__5719\,
            sr => \N__11118\
        );

    \rTxByte_esr_7_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__5734\,
            in1 => \N__10340\,
            in2 => \N__5728\,
            in3 => \N__6013\,
            lcout => \rTxByteZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12790\,
            ce => \N__5719\,
            sr => \N__11118\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1_1_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__12424\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6500\,
            lcout => \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1\,
            ltout => \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_0_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000101"
        )
    port map (
            in0 => \N__6777\,
            in1 => \_gnd_net_\,
            in2 => \N__5701\,
            in3 => \N__6806\,
            lcout => \DUT.fifo_rx_inst.rWritePtrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12784\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI9IJ22_1_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011001111"
        )
    port map (
            in0 => \N__6529\,
            in1 => \N__5698\,
            in2 => \N__5887\,
            in3 => \N__5692\,
            lcout => \DUT.rFifoDatarx_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI96D91_2_1_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6741\,
            in1 => \N__5670\,
            in2 => \N__6783\,
            in3 => \N__5635\,
            lcout => \DUT.fifo_rx_inst.rFifoData_awe3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_1_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011000110"
        )
    port map (
            in0 => \N__6782\,
            in1 => \N__6743\,
            in2 => \N__6811\,
            in3 => \N__5677\,
            lcout => \DUT.fifo_rx_inst.rWritePtrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12784\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5671\,
            in2 => \_gnd_net_\,
            in3 => \N__5634\,
            lcout => \DUT.fifo_rx_inst.N_194\,
            ltout => \DUT.fifo_rx_inst.N_194_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6776\,
            in2 => \N__6055\,
            in3 => \N__6742\,
            lcout => \DUT.fifo_rx_inst.rFifoData_awe0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111110011"
        )
    port map (
            in0 => \N__6052\,
            in1 => \N__6139\,
            in2 => \N__5881\,
            in3 => \N__5947\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIDMJ22_2_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__6043\,
            in1 => \N__6073\,
            in2 => \N__6037\,
            in3 => \N__5861\,
            lcout => \DUT.rFifoDatarx_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__6802\,
            in1 => \N__6778\,
            in2 => \_gnd_net_\,
            in3 => \N__6744\,
            lcout => \DUT.fifo_rx_inst.rFifoData_awe2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111110111111"
        )
    port map (
            in0 => \N__5946\,
            in1 => \N__6570\,
            in2 => \N__5880\,
            in3 => \N__6483\,
            lcout => OPEN,
            ltout => \DUT.rFifoDataror_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rTxByte_6_0_a2_0_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010101"
        )
    port map (
            in0 => \N__10333\,
            in1 => \_gnd_net_\,
            in2 => \N__6025\,
            in3 => \N__6022\,
            lcout => \DUT.uart_inst0.N_257\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101011011"
        )
    port map (
            in0 => \N__5945\,
            in1 => \N__6130\,
            in2 => \N__5878\,
            in3 => \N__6709\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIHQJ22_3_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__5983\,
            in1 => \N__5977\,
            in2 => \N__5968\,
            in3 => \N__5847\,
            lcout => \DUT.rFifoDatarx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__5944\,
            in1 => \N__6703\,
            in2 => \N__5877\,
            in3 => \N__6124\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8459\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12773\,
            ce => \N__6114\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8515\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12773\,
            ce => \N__6114\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7158\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12773\,
            ce => \N__6114\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8460\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12771\,
            ce => \N__6613\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7114\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12771\,
            ce => \N__6613\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_3_LC_14_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__6639\,
            in1 => \N__9349\,
            in2 => \_gnd_net_\,
            in3 => \N__6326\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12826\,
            ce => \N__12340\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_15_LC_14_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9352\,
            in2 => \_gnd_net_\,
            in3 => \N__6937\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12826\,
            ce => \N__12340\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_0_LC_14_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__9351\,
            in1 => \N__9771\,
            in2 => \_gnd_net_\,
            in3 => \N__9575\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12826\,
            ce => \N__12340\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_LC_14_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__9772\,
            in1 => \N__9354\,
            in2 => \_gnd_net_\,
            in3 => \N__9435\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12826\,
            ce => \N__12340\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_4_LC_14_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9348\,
            in2 => \_gnd_net_\,
            in3 => \N__6901\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12826\,
            ce => \N__12340\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_7_LC_14_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8095\,
            in2 => \_gnd_net_\,
            in3 => \N__9353\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12826\,
            ce => \N__12340\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_6_LC_14_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__9350\,
            in1 => \N__6244\,
            in2 => \_gnd_net_\,
            in3 => \N__6854\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12826\,
            ce => \N__12340\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_LC_14_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__11441\,
            in1 => \N__10867\,
            in2 => \N__9046\,
            in3 => \N__8764\,
            lcout => \P1A7_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12826\,
            ce => \N__12340\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIQ3QE2_14_LC_14_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6875\,
            in1 => \N__8195\,
            in2 => \N__6855\,
            in3 => \N__8234\,
            lcout => \DUT.uart_inst0.rx_clk_divider_5_i_a2_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_14_LC_14_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8196\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9363\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12822\,
            ce => \N__12344\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNO_0_5_LC_14_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6368\,
            in1 => \N__8182\,
            in2 => \N__6856\,
            in3 => \N__6151\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_222_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_5_LC_14_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9362\,
            in2 => \N__6157\,
            in3 => \N__6877\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12822\,
            ce => \N__12344\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNI2VEI1_2_LC_14_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7968\,
            in2 => \_gnd_net_\,
            in3 => \N__6900\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.rx_clk_divider_5_i_a2_11_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIQEH13_10_LC_14_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__8343\,
            in1 => \N__6936\,
            in2 => \N__6154\,
            in3 => \N__8361\,
            lcout => \DUT.uart_inst0.rx_clk_divider_5_i_a2_11_5\,
            ltout => \DUT.uart_inst0.rx_clk_divider_5_i_a2_11_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNO_0_6_LC_14_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6876\,
            in1 => \N__8181\,
            in2 => \N__6247\,
            in3 => \N__6367\,
            lcout => \DUT.uart_inst0.N_221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_16_LC_14_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8235\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9364\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12822\,
            ce => \N__12344\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_0_0_c_LC_14_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6387\,
            in2 => \N__6238\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_3_0_\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_0_0_c_RNIPQVSB_LC_14_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7984\,
            in2 => \N__6229\,
            in3 => \N__6220\,
            lcout => \DUT.uart_inst0.rx_countdown_3_1\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_countdown_3_cry_0\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_1_0_c_RNIRV51C_LC_14_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8374\,
            in2 => \N__6217\,
            in3 => \N__6208\,
            lcout => \DUT.uart_inst0.rx_countdown_3_2\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_countdown_3_cry_1\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_2_0_c_RNIT4CLB_LC_14_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6205\,
            in2 => \N__6196\,
            in3 => \N__6187\,
            lcout => \DUT.uart_inst0.rx_countdown_3_3\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_countdown_3_cry_2\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_3_0_c_RNIV9IPB_LC_14_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6184\,
            in2 => \N__9664\,
            in3 => \N__6178\,
            lcout => \DUT.uart_inst0.rx_countdown_3_4\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_countdown_3_cry_3\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_4_0_c_RNI1FOTB_LC_14_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001010101101010"
        )
    port map (
            in0 => \N__8062\,
            in1 => \N__6324\,
            in2 => \N__6375\,
            in3 => \N__6175\,
            lcout => \DUT.uart_inst0.rx_countdown_3_5\,
            ltout => \DUT.uart_inst0.rx_countdown_3_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_2_0_LC_14_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9486\,
            in1 => \N__9421\,
            in2 => \N__6172\,
            in3 => \N__9714\,
            lcout => \DUT.uart_inst0.g3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNITI4IB_0_LC_14_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__6388\,
            in1 => \_gnd_net_\,
            in2 => \N__6376\,
            in3 => \N__6325\,
            lcout => \DUT.uart_inst0.rx_countdown_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_0_3_LC_14_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__8662\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8605\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_196_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_3_LC_14_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011101011"
        )
    port map (
            in0 => \N__9237\,
            in1 => \N__8631\,
            in2 => \N__6292\,
            in3 => \N__8701\,
            lcout => \DUT.uart_inst0.rx_bits_remainingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12815\,
            ce => \N__6286\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_1_1_LC_14_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101100110"
        )
    port map (
            in0 => \N__8660\,
            in1 => \N__8604\,
            in2 => \_gnd_net_\,
            in3 => \N__9235\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_33_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_0_1_LC_14_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000001"
        )
    port map (
            in0 => \N__9712\,
            in1 => \N__8661\,
            in2 => \N__6289\,
            in3 => \N__9627\,
            lcout => \DUT.uart_inst0.rx_bits_remaining_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_3_0_c_RNIP8I482_LC_14_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__9626\,
            in1 => \N__9552\,
            in2 => \N__6268\,
            in3 => \N__9713\,
            lcout => \DUT.uart_inst0.rx_countdown_3_cry_3_0_c_RNIP8IZ0Z482\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_0_LC_14_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__9236\,
            in1 => \_gnd_net_\,
            in2 => \N__8613\,
            in3 => \_gnd_net_\,
            lcout => \DUT.uart_inst0.rx_bits_remainingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12815\,
            ce => \N__6286\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_1_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011010011110000"
        )
    port map (
            in0 => \N__9576\,
            in1 => \N__6274\,
            in2 => \N__8672\,
            in3 => \N__6267\,
            lcout => \DUT.uart_inst0.rx_bits_remainingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rRxRead_esr_RNO_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__10321\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11148\,
            lcout => \P1A2_c_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_4_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100000"
        )
    port map (
            in0 => \N__6468\,
            in1 => \N__9759\,
            in2 => \N__10640\,
            in3 => \N__7252\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_RNIDTQ4_1_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11147\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10369\,
            lcout => \fifo_inst.ftdi_output_inst.rFifoState_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__6400\,
            in1 => \N__11674\,
            in2 => \N__6421\,
            in3 => \N__11536\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__11675\,
            in1 => \N__6433\,
            in2 => \N__6424\,
            in3 => \N__7336\,
            lcout => \DUT.rFifoDatarx_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7371\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12803\,
            ce => \N__10078\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__11535\,
            in1 => \N__6394\,
            in2 => \N__11680\,
            in3 => \N__6412\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7360\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12796\,
            ce => \N__6559\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7312\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12796\,
            ce => \N__6559\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10141\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12796\,
            ce => \N__6559\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7279\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12796\,
            ce => \N__6559\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7516\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12796\,
            ce => \N__6559\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7438\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12796\,
            ce => \N__6559\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7583\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12796\,
            ce => \N__6559\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10102\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12796\,
            ce => \N__6559\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7237\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12791\,
            ce => \N__6617\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7051\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12791\,
            ce => \N__6617\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7012\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12791\,
            ce => \N__6617\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_3_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6484\,
            in2 => \_gnd_net_\,
            in3 => \N__6501\,
            lcout => \DUT.fifo_rx_inst.rFifoDataro_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12785\,
            ce => 'H',
            sr => \N__11113\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_0_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7717\,
            in2 => \_gnd_net_\,
            in3 => \N__10027\,
            lcout => \DUT.fifo_tx_inst.rFifoDataro_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12785\,
            ce => 'H',
            sr => \N__11113\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_1_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7704\,
            in2 => \_gnd_net_\,
            in3 => \N__6552\,
            lcout => \DUT.fifo_tx_inst.rFifoDataro_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12785\,
            ce => 'H',
            sr => \N__11113\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_3_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7393\,
            in2 => \_gnd_net_\,
            in3 => \N__7729\,
            lcout => \DUT.fifo_tx_inst.rFifoDataro_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12785\,
            ce => 'H',
            sr => \N__11113\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_2_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6571\,
            in2 => \_gnd_net_\,
            in3 => \N__6594\,
            lcout => \DUT.fifo_rx_inst.rFifoDataro_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12785\,
            ce => 'H',
            sr => \N__11113\
        );

    \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_0_1_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__7646\,
            in1 => \N__7612\,
            in2 => \_gnd_net_\,
            in3 => \N__8982\,
            lcout => \DUT.fifo_tx_inst.rFifoData_awe1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_1_1_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__8983\,
            in1 => \_gnd_net_\,
            in2 => \N__7618\,
            in3 => \N__7647\,
            lcout => \DUT.fifo_tx_inst.rFifoData_awe0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_1_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000010010"
        )
    port map (
            in0 => \N__7617\,
            in1 => \N__6538\,
            in2 => \N__7654\,
            in3 => \N__8985\,
            lcout => \DUT.fifo_tx_inst.rWritePtrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12779\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNI8BKM_2_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__7611\,
            in1 => \N__10222\,
            in2 => \N__7653\,
            in3 => \N__9919\,
            lcout => \DUT.fifo_tx_inst.rFifoData_awe3\,
            ltout => \DUT.fifo_tx_inst.rFifoData_awe3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNI4PUO_2_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6541\,
            in3 => \N__12428\,
            lcout => \DUT.fifo_tx_inst.un1_i11_i\,
            ltout => \DUT.fifo_tx_inst.un1_i11_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_0_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000101"
        )
    port map (
            in0 => \N__8984\,
            in1 => \_gnd_net_\,
            in2 => \N__6532\,
            in3 => \N__7648\,
            lcout => \DUT.fifo_tx_inst.rWritePtrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12779\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6810\,
            in1 => \N__6784\,
            in2 => \_gnd_net_\,
            in3 => \N__6748\,
            lcout => \DUT.fifo_rx_inst.rFifoData_awe1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7105\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12776\,
            ce => \N__6682\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8506\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12776\,
            ce => \N__6682\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7150\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12776\,
            ce => \N__6682\,
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_15_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8115\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_1_0_\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNID95P_1_LC_15_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12944\,
            in2 => \N__8071\,
            in3 => \N__6655\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_1\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_0\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIFC6P_2_LC_15_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12953\,
            in2 => \N__7957\,
            in3 => \N__6652\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_2\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_1\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIHF7P_3_LC_15_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12945\,
            in2 => \N__6649\,
            in3 => \N__6625\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_3\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_2\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIJI8P_4_LC_15_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6907\,
            in2 => \N__12996\,
            in3 => \N__6889\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_4\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_3\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNILL9P_5_LC_15_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12949\,
            in2 => \N__6886\,
            in3 => \N__6865\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_5\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_4\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNINOAP_6_LC_15_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6862\,
            in2 => \N__12997\,
            in3 => \N__6835\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_6\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_5\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIPRBP_7_LC_15_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6832\,
            in2 => \N__12998\,
            in3 => \N__6826\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_7\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_6\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIRUCP_8_LC_15_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7759\,
            in2 => \N__13078\,
            in3 => \N__6823\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_8\,
            ltout => OPEN,
            carryin => \bfn_15_2_0_\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIT1EP_9_LC_15_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8152\,
            in2 => \N__13075\,
            in3 => \N__6820\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_9\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_8\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNI6KQI_10_LC_15_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8332\,
            in2 => \N__13076\,
            in3 => \N__6817\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_10\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_9\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIFEUD_11_LC_15_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8137\,
            in2 => \N__13072\,
            in3 => \N__6814\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_11\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_10\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIHHVD_12_LC_15_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8122\,
            in2 => \N__13077\,
            in3 => \N__6961\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_12\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_11\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIJK0E_13_LC_15_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8314\,
            in2 => \N__13073\,
            in3 => \N__6958\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_13\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_12\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNILN1E_14_LC_15_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13055\,
            in2 => \N__6955\,
            in3 => \N__6946\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_14\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_13\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNINQ2E_15_LC_15_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6943\,
            in2 => \N__13074\,
            in3 => \N__6925\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_15\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_14\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIPT3E_16_LC_15_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6922\,
            in2 => \N__13071\,
            in3 => \N__6916\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_16\,
            ltout => OPEN,
            carryin => \bfn_15_3_0_\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIR05E_17_LC_15_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8350\,
            in2 => \_gnd_net_\,
            in3 => \N__6913\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_15_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000100"
        )
    port map (
            in0 => \N__8026\,
            in1 => \N__8556\,
            in2 => \N__9869\,
            in3 => \N__9241\,
            lcout => \DUT.uart_inst0.g0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_2_4_LC_15_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9746\,
            in1 => \N__8022\,
            in2 => \N__9430\,
            in3 => \N__9705\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.recv_state_RNO_2Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_1_4_LC_15_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6910\,
            in3 => \N__9625\,
            lcout => \DUT.uart_inst0.G_11_i_a4_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_2_2_LC_15_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010100000000"
        )
    port map (
            in0 => \N__9747\,
            in1 => \N__9860\,
            in2 => \N__8284\,
            in3 => \N__9487\,
            lcout => \DUT.uart_inst0.g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNI1K9CC_2_LC_15_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10638\,
            in2 => \N__8039\,
            in3 => \N__8555\,
            lcout => \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa_0_a2_0_a2_0_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_15_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__9551\,
            in1 => \_gnd_net_\,
            in2 => \N__9431\,
            in3 => \N__9706\,
            lcout => \DUT.uart_inst0.g0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNIM4BC72_2_LC_15_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__9628\,
            in1 => \N__6982\,
            in2 => \N__9571\,
            in3 => \N__6972\,
            lcout => \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_5_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__8030\,
            in1 => \N__9556\,
            in2 => \_gnd_net_\,
            in3 => \N__9630\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.rx_countdown_8_i_0_o2_1_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_5_LC_15_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__8719\,
            in1 => \N__10633\,
            in2 => \N__6976\,
            in3 => \N__6973\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12818\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_1_0_c_RNINE4G31_LC_15_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9417\,
            in2 => \N__9497\,
            in3 => \N__9707\,
            lcout => \DUT.uart_inst0.recv_state_ns_0_i_0_0_o2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_1_0_c_RNIHVHJ31_LC_15_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__9419\,
            in1 => \N__9479\,
            in2 => \_gnd_net_\,
            in3 => \N__8029\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.G_9_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_3_0_c_RNIEB1T62_LC_15_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__9558\,
            in1 => \N__9629\,
            in2 => \N__6964\,
            in3 => \N__9711\,
            lcout => \DUT.uart_inst0.N_193\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_2_1_LC_15_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__9418\,
            in1 => \N__9316\,
            in2 => \N__9720\,
            in3 => \N__8028\,
            lcout => \DUT.uart_inst0.recv_state_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_4_LC_15_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010100000000"
        )
    port map (
            in0 => \N__9557\,
            in1 => \N__9420\,
            in2 => \N__9498\,
            in3 => \N__7258\,
            lcout => \DUT.uart_inst0.N_4_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_1_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8430\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.wRxByte_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12816\,
            ce => \N__8418\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_0_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7214\,
            lcout => \DUT.wRxByte_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12816\,
            ce => \N__8418\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_3_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7130\,
            lcout => \DUT.wRxByte_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12816\,
            ce => \N__8418\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_4_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7085\,
            lcout => \DUT.wRxByte_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12816\,
            ce => \N__8418\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_5_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7040\,
            lcout => \DUT.wRxByte_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12816\,
            ce => \N__8418\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_6_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7000\,
            lcout => \DUT.wRxByte_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12816\,
            ce => \N__8418\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_7_LC_15_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9855\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.wRxByte_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12816\,
            ce => \N__8418\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7329\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12810\,
            ce => \N__7413\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10158\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12810\,
            ce => \N__7413\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7294\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12810\,
            ce => \N__7413\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7528\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12810\,
            ce => \N__7413\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7456\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12810\,
            ce => \N__7413\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10120\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12810\,
            ce => \N__7413\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7370\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12804\,
            ce => \N__7948\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7322\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12804\,
            ce => \N__7948\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10151\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12804\,
            ce => \N__7948\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7289\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12804\,
            ce => \N__7948\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7526\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12804\,
            ce => \N__7948\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7448\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12804\,
            ce => \N__7948\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7590\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12804\,
            ce => \N__7948\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10112\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12804\,
            ce => \N__7948\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__11540\,
            in1 => \N__7555\,
            in2 => \N__7492\,
            in3 => \N__11661\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__11666\,
            in1 => \N__7549\,
            in2 => \N__7540\,
            in3 => \N__7537\,
            lcout => \DUT.rFifoDatarx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7527\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12797\,
            ce => \N__10061\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111110011"
        )
    port map (
            in0 => \N__7483\,
            in1 => \N__7420\,
            in2 => \N__11678\,
            in3 => \N__11541\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__7477\,
            in1 => \N__7468\,
            in2 => \N__7459\,
            in3 => \N__11665\,
            lcout => \DUT.rFifoDatarx_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7455\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12797\,
            ce => \N__10061\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100100111"
        )
    port map (
            in0 => \N__11539\,
            in1 => \N__7753\,
            in2 => \N__7747\,
            in3 => \N__11660\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111101111111"
        )
    port map (
            in0 => \N__7728\,
            in1 => \N__11522\,
            in2 => \N__11676\,
            in3 => \N__7930\,
            lcout => \DUT.rFifoDataror_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_0_RNI86BE_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100011011"
        )
    port map (
            in0 => \N__11523\,
            in1 => \N__7716\,
            in2 => \N__7705\,
            in3 => \N__11651\,
            lcout => OPEN,
            ltout => \DUT.rFifoDataror_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNIQOK61_0_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7690\,
            in2 => \N__7684\,
            in3 => \N__11434\,
            lcout => \DUT.uart_inst0.N_145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_15_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__11652\,
            in1 => \N__7681\,
            in2 => \N__7672\,
            in3 => \N__7660\,
            lcout => \DUT.rFifoDatarx_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNI7FOF_2_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10217\,
            in2 => \_gnd_net_\,
            in3 => \N__9910\,
            lcout => \DUT.fifo_tx_inst.N_79\,
            ltout => \DUT.fifo_tx_inst.N_79_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_1_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7652\,
            in2 => \N__7621\,
            in3 => \N__7616\,
            lcout => \DUT.fifo_tx_inst.rFifoData_awe2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_RNIFFVH_4_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7895\,
            in2 => \_gnd_net_\,
            in3 => \N__7913\,
            lcout => \fifo_inst.ftdi_output_inst.N_68_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_0_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100110100101"
        )
    port map (
            in0 => \N__10001\,
            in1 => \N__9940\,
            in2 => \N__8989\,
            in3 => \N__11754\,
            lcout => \DUT.fifo_tx_inst.rFifoCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12780\,
            ce => 'H',
            sr => \N__11111\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_2_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7941\,
            in2 => \_gnd_net_\,
            in3 => \N__7929\,
            lcout => \DUT.fifo_tx_inst.rFifoDataro_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12780\,
            ce => 'H',
            sr => \N__11111\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_3_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__11044\,
            in1 => \N__11241\,
            in2 => \_gnd_net_\,
            in3 => \N__10975\,
            lcout => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12780\,
            ce => 'H',
            sr => \N__11111\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_4_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100001010"
        )
    port map (
            in0 => \N__7915\,
            in1 => \_gnd_net_\,
            in2 => \N__7900\,
            in3 => \N__7881\,
            lcout => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12780\,
            ce => 'H',
            sr => \N__11111\
        );

    \fifo_inst.ftdi_output_inst.rWrDelay_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7896\,
            in2 => \_gnd_net_\,
            in3 => \N__7914\,
            lcout => \fifo_inst.ftdi_output_inst.rWrDelayZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12780\,
            ce => 'H',
            sr => \N__11111\
        );

    \fifo_inst.ftdi_output_inst.oTx_n_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__11171\,
            in1 => \N__7847\,
            in2 => \_gnd_net_\,
            in3 => \N__7882\,
            lcout => \P1A4_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12780\,
            ce => 'H',
            sr => \N__11111\
        );

    \fifo_inst.ftdi_output_inst.rTxBusReady_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__7784\,
            in1 => \N__8995\,
            in2 => \_gnd_net_\,
            in3 => \N__11170\,
            lcout => \rTxBusReady\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12780\,
            ce => 'H',
            sr => \N__11111\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIO0PE2_11_LC_16_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7767\,
            in1 => \N__8130\,
            in2 => \N__8166\,
            in3 => \N__8145\,
            lcout => \DUT.uart_inst0.rx_clk_divider_5_i_a2_12_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_8_LC_16_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__9319\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7768\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12832\,
            ce => \N__12345\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_9_LC_16_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8167\,
            in3 => \N__9318\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12832\,
            ce => \N__12345\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_11_LC_16_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__8146\,
            in1 => \_gnd_net_\,
            in2 => \N__9346\,
            in3 => \_gnd_net_\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12832\,
            ce => \N__12345\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_12_LC_16_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9317\,
            in2 => \_gnd_net_\,
            in3 => \N__8131\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12832\,
            ce => \N__12345\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_0_LC_16_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__9320\,
            in1 => \N__8114\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12832\,
            ce => \N__12345\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIS5BA2_0_LC_16_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__8325\,
            in1 => \N__8079\,
            in2 => \N__8116\,
            in3 => \N__8091\,
            lcout => \DUT.uart_inst0.rx_clk_divider_5_i_a2_12_4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_LC_16_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__8080\,
            in1 => \_gnd_net_\,
            in2 => \N__9347\,
            in3 => \_gnd_net_\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12832\,
            ce => \N__12345\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_5_LC_16_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__9311\,
            in1 => \N__9761\,
            in2 => \_gnd_net_\,
            in3 => \N__9651\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12829\,
            ce => \N__12346\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_1_LC_16_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100110011"
        )
    port map (
            in0 => \N__9760\,
            in1 => \N__9313\,
            in2 => \_gnd_net_\,
            in3 => \N__8046\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12829\,
            ce => \N__12346\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_2_LC_16_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9310\,
            in2 => \_gnd_net_\,
            in3 => \N__7972\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12829\,
            ce => \N__12346\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_2_LC_16_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__8395\,
            in1 => \N__8389\,
            in2 => \N__8383\,
            in3 => \N__9652\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12829\,
            ce => \N__12346\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_17_LC_16_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9309\,
            in2 => \_gnd_net_\,
            in3 => \N__8362\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12829\,
            ce => \N__12346\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_10_LC_16_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9312\,
            in2 => \_gnd_net_\,
            in3 => \N__8344\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12829\,
            ce => \N__12346\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_13_LC_16_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9308\,
            in2 => \_gnd_net_\,
            in3 => \N__8326\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12829\,
            ce => \N__12346\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_3_2_LC_16_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__9862\,
            in1 => \N__8554\,
            in2 => \_gnd_net_\,
            in3 => \N__9222\,
            lcout => \DUT.uart_inst0.N_199_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ioFifoData_iobuf_RNO_0_LC_16_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__11266\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_1239_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNI237O_0_LC_16_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9861\,
            in2 => \_gnd_net_\,
            in3 => \N__8280\,
            lcout => \DUT.uart_inst0.N_149\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_3_LC_16_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011000000"
        )
    port map (
            in0 => \N__9802\,
            in1 => \N__8713\,
            in2 => \N__10642\,
            in3 => \N__8569\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12827\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNI2S9L5_0_LC_16_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__8256\,
            in1 => \N__8236\,
            in2 => \N__8221\,
            in3 => \N__8197\,
            lcout => \DUT.uart_inst0.rx_clk_divider_5_i_a2_12_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNO_2_2_LC_16_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111110"
        )
    port map (
            in0 => \N__9223\,
            in1 => \N__8706\,
            in2 => \N__8617\,
            in3 => \N__8674\,
            lcout => \DUT.uart_inst0.N_31_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_1_5_LC_16_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__9882\,
            in1 => \N__9801\,
            in2 => \_gnd_net_\,
            in3 => \N__9220\,
            lcout => \DUT.uart_inst0.N_203\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_3_LC_16_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8552\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8581\,
            lcout => \DUT.uart_inst0.recv_state_ns_0_i_0_0_a3_0_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNIUJI11_3_LC_16_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__8707\,
            in1 => \N__8673\,
            in2 => \N__8635\,
            in3 => \N__8609\,
            lcout => \DUT.uart_inst0.N_215_4\,
            ltout => \DUT.uart_inst0.N_215_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_2_LC_16_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101110"
        )
    port map (
            in0 => \N__9221\,
            in1 => \N__8557\,
            in2 => \N__8575\,
            in3 => \N__9881\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.recv_state_srsts_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_2_LC_16_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__10634\,
            in1 => \N__8553\,
            in2 => \N__8572\,
            in3 => \N__8568\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12823\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNIBTG71_2_LC_16_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010001000"
        )
    port map (
            in0 => \N__12423\,
            in1 => \N__8551\,
            in2 => \N__9883\,
            in3 => \N__9219\,
            lcout => \DUT.uart_inst0.g0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_2_LC_16_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8482\,
            lcout => \DUT.wRxByte_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12819\,
            ce => \N__8419\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__8875\,
            in1 => \N__11659\,
            in2 => \N__8869\,
            in3 => \N__8824\,
            lcout => \DUT.rFifoDatarx_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__11658\,
            in1 => \N__8860\,
            in2 => \N__8854\,
            in3 => \N__8845\,
            lcout => \DUT.rFifoDatarx_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__11537\,
            in1 => \N__8836\,
            in2 => \N__11677\,
            in3 => \N__10126\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111001111"
        )
    port map (
            in0 => \N__8818\,
            in1 => \N__11656\,
            in2 => \N__8806\,
            in3 => \N__11538\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__11657\,
            in1 => \N__8791\,
            in2 => \N__8785\,
            in3 => \N__8782\,
            lcout => \DUT.rFifoDatarx_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_0_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__8776\,
            in1 => \N__9148\,
            in2 => \N__8743\,
            in3 => \N__11436\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12811\,
            ce => \N__9102\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_RNO_0_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111110"
        )
    port map (
            in0 => \N__8902\,
            in1 => \N__8908\,
            in2 => \N__9007\,
            in3 => \N__10859\,
            lcout => \DUT.uart_inst0.tx_out_6_iv_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_1_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__8959\,
            in1 => \N__8749\,
            in2 => \N__11443\,
            in3 => \N__9149\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12811\,
            ce => \N__9102\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_2_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__11435\,
            in1 => \N__8734\,
            in2 => \N__9154\,
            in3 => \N__8947\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12811\,
            ce => \N__9102\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_3_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__8953\,
            in1 => \N__9153\,
            in2 => \N__9172\,
            in3 => \N__11437\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12811\,
            ce => \N__9102\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__11542\,
            in1 => \N__8938\,
            in2 => \N__11679\,
            in3 => \N__10087\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101100001011"
        )
    port map (
            in0 => \N__8926\,
            in1 => \N__11670\,
            in2 => \N__8917\,
            in3 => \N__8914\,
            lcout => \DUT.rFifoDatarx_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNINQKO8_0_0_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000110000"
        )
    port map (
            in0 => \N__11433\,
            in1 => \N__11461\,
            in2 => \N__12441\,
            in3 => \N__10852\,
            lcout => \DUT.uart_inst0.N_22_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_RNO_1_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__11821\,
            in1 => \N__11432\,
            in2 => \N__9081\,
            in3 => \N__10769\,
            lcout => \DUT.uart_inst0.tx_out_6_iv_0_a3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_RNO_3_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010001100"
        )
    port map (
            in0 => \N__10770\,
            in1 => \N__9053\,
            in2 => \N__11442\,
            in3 => \N__11746\,
            lcout => \DUT.uart_inst0.N_101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_5_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__11406\,
            in1 => \N__8896\,
            in2 => \N__8884\,
            in3 => \N__9137\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12798\,
            ce => \N__9109\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_6_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__9138\,
            in1 => \N__8890\,
            in2 => \N__9118\,
            in3 => \N__11408\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12798\,
            ce => \N__9109\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_4_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__9136\,
            in1 => \N__9187\,
            in2 => \N__9181\,
            in3 => \N__11407\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12798\,
            ce => \N__9109\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_7_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9160\,
            in2 => \_gnd_net_\,
            in3 => \N__9135\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12798\,
            ce => \N__9109\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNI0AJL_0_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10218\,
            in2 => \_gnd_net_\,
            in3 => \N__11832\,
            lcout => \DUT.fifo_tx_inst.N_83\,
            ltout => \DUT.fifo_tx_inst.N_83_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNISSQ21_1_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__11749\,
            in1 => \_gnd_net_\,
            in2 => \N__9085\,
            in3 => \N__9963\,
            lcout => \DUT.fifo_tx_inst.rFifoCount_RNISSQ21Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_RNO_2_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011000000"
        )
    port map (
            in0 => \N__9082\,
            in1 => \N__11801\,
            in2 => \N__9064\,
            in3 => \N__11370\,
            lcout => \DUT.uart_inst0.N_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_RNI7AJQ_0_0_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__11054\,
            in1 => \N__11250\,
            in2 => \_gnd_net_\,
            in3 => \N__10939\,
            lcout => \fifo_inst.ftdi_output_inst.rFifoStatec_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNIN9O8_0_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__9906\,
            in1 => \N__9961\,
            in2 => \_gnd_net_\,
            in3 => \N__9993\,
            lcout => \DUT.N_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNIME2J_0_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__9962\,
            in1 => \N__9994\,
            in2 => \N__9915\,
            in3 => \N__11747\,
            lcout => \DUT.fifo_tx_inst.rReadPtr11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__11748\,
            in1 => \N__8981\,
            in2 => \N__10002\,
            in3 => \N__9938\,
            lcout => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10009\,
            in2 => \N__10003\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_11_0_\,
            carryout => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_1_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9964\,
            in2 => \N__9973\,
            in3 => \N__9943\,
            lcout => \DUT.fifo_tx_inst.rFifoCountZ0Z_1\,
            ltout => OPEN,
            carryin => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0\,
            carryout => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1\,
            clk => \N__12786\,
            ce => 'H',
            sr => \N__11114\
        );

    \DUT.fifo_tx_inst.rFifoCount_2_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110010110011010"
        )
    port map (
            in0 => \N__9914\,
            in1 => \N__9939\,
            in2 => \N__11755\,
            in3 => \N__9922\,
            lcout => \DUT.fifo_tx_inst.rFifoCountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12786\,
            ce => 'H',
            sr => \N__11114\
        );

    \DUT.uart_inst0.recv_state_RNO_0_6_LC_17_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9870\,
            in1 => \N__12422\,
            in2 => \_gnd_net_\,
            in3 => \N__9800\,
            lcout => \DUT.uart_inst0.g0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_4_LC_17_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__9770\,
            in1 => \N__9314\,
            in2 => \_gnd_net_\,
            in3 => \N__9721\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12830\,
            ce => \N__12353\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_1_1_LC_17_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9650\,
            in2 => \_gnd_net_\,
            in3 => \N__9586\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.G_10_i_a4_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_1_LC_17_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000010000"
        )
    port map (
            in0 => \N__9577\,
            in1 => \N__9505\,
            in2 => \N__9439\,
            in3 => \N__9436\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_4_i_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_1_LC_17_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001010"
        )
    port map (
            in0 => \N__10641\,
            in1 => \N__9234\,
            in2 => \N__9367\,
            in3 => \N__9315\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12828\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_0_LC_17_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001011001"
        )
    port map (
            in0 => \N__10403\,
            in1 => \N__10456\,
            in2 => \N__10252\,
            in3 => \N__10432\,
            lcout => \DUT.fifo_rx_inst.rFifoCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12824\,
            ce => 'H',
            sr => \N__11130\
        );

    \fifo_inst.ftdi_output_inst.oRxFlag_LC_17_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111001100"
        )
    port map (
            in0 => \N__10790\,
            in1 => \N__10367\,
            in2 => \_gnd_net_\,
            in3 => \N__10302\,
            lcout => \P1A2_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12824\,
            ce => 'H',
            sr => \N__11130\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_2_LC_17_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10368\,
            lcout => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12824\,
            ce => 'H',
            sr => \N__11130\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_1_LC_17_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11059\,
            in2 => \_gnd_net_\,
            in3 => \N__10970\,
            lcout => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12824\,
            ce => 'H',
            sr => \N__11130\
        );

    \rTxWrite_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10301\,
            in2 => \_gnd_net_\,
            in3 => \N__10251\,
            lcout => \rTxWriteZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12820\,
            ce => 'H',
            sr => \N__11129\
        );

    \fifo_inst.ftdi_output_inst.oRx_n_LC_17_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__10791\,
            in1 => \N__10175\,
            in2 => \_gnd_net_\,
            in3 => \N__10906\,
            lcout => \P1A3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12820\,
            ce => 'H',
            sr => \N__11129\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10159\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12817\,
            ce => \N__10081\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10116\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12817\,
            ce => \N__10081\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__10660\,
            in1 => \N__10695\,
            in2 => \N__10683\,
            in3 => \N__10495\,
            lcout => \DUT.uart_inst0.un1_tx_bits_remaining_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_2_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101001"
        )
    port map (
            in0 => \N__10696\,
            in1 => \N__10682\,
            in2 => \N__10501\,
            in3 => \N__10663\,
            lcout => \DUT.uart_inst0.tx_bits_remainingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12812\,
            ce => 'H',
            sr => \N__11845\
        );

    \DUT.uart_inst0.tx_bits_remaining_1_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010100101"
        )
    port map (
            in0 => \N__10662\,
            in1 => \_gnd_net_\,
            in2 => \N__10684\,
            in3 => \N__10497\,
            lcout => \DUT.uart_inst0.tx_bits_remainingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12812\,
            ce => 'H',
            sr => \N__11845\
        );

    \DUT.uart_inst0.tx_bits_remaining_0_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__10496\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10661\,
            lcout => \DUT.uart_inst0.tx_bits_remainingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12812\,
            ce => 'H',
            sr => \N__11845\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_3_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10694\,
            in1 => \N__10675\,
            in2 => \N__10471\,
            in3 => \N__10659\,
            lcout => \DUT.uart_inst0.N_142\,
            ltout => \DUT.uart_inst0.N_142_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNIJ5C81_1_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11804\,
            in2 => \N__10645\,
            in3 => \N__11391\,
            lcout => \DUT.uart_inst0.N_144\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNI6Q5N3_1_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__11392\,
            in1 => \N__10726\,
            in2 => \N__11818\,
            in3 => \N__10771\,
            lcout => \DUT.uart_inst0.N_146\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNI3MLP6_3_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100001010"
        )
    port map (
            in0 => \N__12244\,
            in1 => \_gnd_net_\,
            in2 => \N__10888\,
            in3 => \N__10721\,
            lcout => \DUT.uart_inst0.N_84\,
            ltout => \DUT.uart_inst0.N_84_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNINQKO8_0_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111011101"
        )
    port map (
            in0 => \N__10625\,
            in1 => \N__11459\,
            in2 => \N__10504\,
            in3 => \N__11395\,
            lcout => \DUT.uart_inst0.N_22\,
            ltout => \DUT.uart_inst0.N_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_3_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111110111010111"
        )
    port map (
            in0 => \N__10897\,
            in1 => \N__10470\,
            in2 => \N__10480\,
            in3 => \N__10477\,
            lcout => \DUT.uart_inst0.tx_bits_remainingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNICODU_0_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10768\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11394\,
            lcout => \DUT.uart_inst0.N_143\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_RNO_0_0_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11254\,
            in1 => \N__11055\,
            in2 => \_gnd_net_\,
            in3 => \N__10946\,
            lcout => OPEN,
            ltout => \fifo_inst.ftdi_output_inst.N_78_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_0_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__10795\,
            in1 => \N__12433\,
            in2 => \N__10774\,
            in3 => \N__11182\,
            lcout => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12805\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNIIAMI1_1_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111110001"
        )
    port map (
            in0 => \N__11393\,
            in1 => \N__11712\,
            in2 => \N__11819\,
            in3 => \N__10767\,
            lcout => \DUT.uart_inst0.N_74\,
            ltout => \DUT.uart_inst0.N_74_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNILHU57_1_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__10747\,
            in1 => \N__10883\,
            in2 => \N__10741\,
            in3 => \N__12243\,
            lcout => \DUT.uart_inst0.tx_countdown_7s2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNIFE3O7_0_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000000010000"
        )
    port map (
            in0 => \N__12224\,
            in1 => \N__10725\,
            in2 => \N__10738\,
            in3 => \N__10887\,
            lcout => \DUT.uart_inst0.N_30_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNI45HK1_2_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12133\,
            in1 => \N__12006\,
            in2 => \N__12049\,
            in3 => \N__11976\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNIJKPE2_3_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__11874\,
            in1 => \_gnd_net_\,
            in2 => \N__10729\,
            in3 => \N__12079\,
            lcout => \DUT.uart_inst0.N_75\,
            ltout => \DUT.uart_inst0.N_75_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNIBVOQB_0_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100000"
        )
    port map (
            in0 => \N__11371\,
            in1 => \N__12223\,
            in2 => \N__10705\,
            in3 => \N__10702\,
            lcout => \DUT.uart_inst0.tx_countdown_7_sm0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNI34HK1_2_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__11975\,
            in1 => \N__12132\,
            in2 => \N__12010\,
            in3 => \N__12078\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_state_ns_i_i_o2_a0_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNIJKPE2_0_3_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__12042\,
            in1 => \_gnd_net_\,
            in2 => \N__10891\,
            in3 => \N__11873\,
            lcout => \DUT.uart_inst0.N_69_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_0_2_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111000001111"
        )
    port map (
            in0 => \N__12084\,
            in1 => \N__12046\,
            in2 => \N__12139\,
            in3 => \N__12245\,
            lcout => \DUT.uart_inst0.tx_countdown_7_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100001"
        )
    port map (
            in0 => \N__12045\,
            in1 => \N__12135\,
            in2 => \N__11884\,
            in3 => \N__12083\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_countdown_30_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100001111"
        )
    port map (
            in0 => \N__11882\,
            in1 => \N__12246\,
            in2 => \N__10870\,
            in3 => \N__11917\,
            lcout => \DUT.uart_inst0.tx_countdown_7_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_1_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__10827\,
            in1 => \N__10860\,
            in2 => \_gnd_net_\,
            in3 => \N__11802\,
            lcout => \DUT.tx_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12792\,
            ce => 'H',
            sr => \N__11119\
        );

    \DUT.uart_inst0.tx_state_0_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__10828\,
            in1 => \N__11753\,
            in2 => \N__11427\,
            in3 => \N__11803\,
            lcout => \DUT.tx_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12792\,
            ce => 'H',
            sr => \N__11119\
        );

    \ioFifoData_iobuf_RNO_3_LC_18_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__11275\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_1242_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ioFifoData_iobuf_RNO_1_LC_18_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__11281\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_1240_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rTxBusReady_rep1_i_ess_LC_18_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111010111111111"
        )
    port map (
            in0 => \N__10972\,
            in1 => \_gnd_net_\,
            in2 => \N__11249\,
            in3 => \N__11041\,
            lcout => \rTxBusReady_rep1_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12831\,
            ce => \N__11065\,
            sr => \N__11134\
        );

    \fifo_inst.ftdi_output_inst.rTxBusReady_rep3_i_ess_LC_18_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__11043\,
            in1 => \N__11240\,
            in2 => \_gnd_net_\,
            in3 => \N__10974\,
            lcout => \rTxBusReady_rep3_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12831\,
            ce => \N__11065\,
            sr => \N__11134\
        );

    \fifo_inst.ftdi_output_inst.rTxBusReady_rep0_i_ess_LC_18_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__11040\,
            in1 => \N__11235\,
            in2 => \_gnd_net_\,
            in3 => \N__10971\,
            lcout => \rTxBusReady_rep0_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12831\,
            ce => \N__11065\,
            sr => \N__11134\
        );

    \fifo_inst.ftdi_output_inst.rTxBusReady_rep2_i_ess_LC_18_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__11042\,
            in1 => \N__11239\,
            in2 => \_gnd_net_\,
            in3 => \N__10973\,
            lcout => \rTxBusReady_rep2_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12831\,
            ce => \N__11065\,
            sr => \N__11134\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_RNIMPIC1_0_LC_18_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__11039\,
            in1 => \N__10969\,
            in2 => \N__11248\,
            in3 => \N__11181\,
            lcout => OPEN,
            ltout => \fifo_inst.ftdi_output_inst.un1_oTx_n_1_sqmuxa_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_RNII7TE1_0_LC_18_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__11149\,
            in1 => \_gnd_net_\,
            in2 => \N__11068\,
            in3 => \_gnd_net_\,
            lcout => \fifo_inst.ftdi_output_inst.un1_oTx_n_1_sqmuxa_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_RNIR68B_0_LC_18_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11038\,
            in2 => \_gnd_net_\,
            in3 => \N__10956\,
            lcout => \fifo_inst.ftdi_output_inst.N_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNICU6U_1_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__11808\,
            in1 => \N__11711\,
            in2 => \_gnd_net_\,
            in3 => \N__11428\,
            lcout => \DUT.uart_inst0.N_77\,
            ltout => \DUT.uart_inst0.N_77_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNI8CH01_1_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10900\,
            in3 => \N__12432\,
            lcout => \DUT.uart_inst0.tx_state_RNI8CH01Z0Z_1\,
            ltout => \DUT.uart_inst0.tx_state_RNI8CH01Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNI8CH01_0_1_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11848\,
            in3 => \_gnd_net_\,
            lcout => \DUT.uart_inst0.N_59_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.rTransmit_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__11423\,
            in1 => \N__11839\,
            in2 => \N__11820\,
            in3 => \N__12437\,
            lcout => \DUT.rTransmitZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rReadPtr_1_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__11563\,
            in1 => \N__11603\,
            in2 => \N__11534\,
            in3 => \N__11569\,
            lcout => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rReadPtr_RNILV421_0_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__11602\,
            in1 => \N__11507\,
            in2 => \N__12442\,
            in3 => \N__11561\,
            lcout => \DUT.fifo_tx_inst.un1_i11_2_i\,
            ltout => \DUT.fifo_tx_inst.un1_i11_2_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rReadPtr_0_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__11562\,
            in1 => \_gnd_net_\,
            in2 => \N__11545\,
            in3 => \N__11511\,
            lcout => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12813\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_1_2_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__11953\,
            in1 => \N__11460\,
            in2 => \_gnd_net_\,
            in3 => \N__11422\,
            lcout => \DUT.uart_inst0.N_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_0_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101001000000"
        )
    port map (
            in0 => \N__12085\,
            in1 => \N__12281\,
            in2 => \N__12250\,
            in3 => \N__11920\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12806\,
            ce => \N__12375\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_4_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001101101000100"
        )
    port map (
            in0 => \N__11918\,
            in1 => \N__12109\,
            in2 => \N__12247\,
            in3 => \N__11980\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12806\,
            ce => \N__12375\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_2_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101111111"
        )
    port map (
            in0 => \N__11296\,
            in1 => \N__12230\,
            in2 => \N__11290\,
            in3 => \N__11921\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12806\,
            ce => \N__12375\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_5_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001101101000100"
        )
    port map (
            in0 => \N__11919\,
            in1 => \N__12091\,
            in2 => \N__12248\,
            in3 => \N__12009\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12806\,
            ce => \N__12375\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNIUUGK1_2_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12044\,
            in1 => \N__12134\,
            in2 => \N__11883\,
            in3 => \N__12081\,
            lcout => \DUT.uart_inst0.tx_countdown_0_c4\,
            ltout => \DUT.uart_inst0.tx_countdown_0_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_0_4_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100101110"
        )
    port map (
            in0 => \N__11978\,
            in1 => \N__12157\,
            in2 => \N__12112\,
            in3 => \N__11942\,
            lcout => \DUT.uart_inst0.tx_countdown_7_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_0_1_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011111110"
        )
    port map (
            in0 => \N__11943\,
            in1 => \N__12047\,
            in2 => \N__12163\,
            in3 => \N__12082\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_countdown_7_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_1_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001001011010"
        )
    port map (
            in0 => \N__12048\,
            in1 => \N__12249\,
            in2 => \N__12103\,
            in3 => \N__11925\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12799\,
            ce => \N__12376\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_0_5_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001001110"
        )
    port map (
            in0 => \N__12158\,
            in1 => \N__12008\,
            in2 => \N__12100\,
            in3 => \N__11979\,
            lcout => \DUT.uart_inst0.tx_countdown_7_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_3_2_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__12080\,
            in1 => \N__11875\,
            in2 => \_gnd_net_\,
            in3 => \N__12043\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_countdown_7_m1_0_o2_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_2_2_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12007\,
            in2 => \N__11983\,
            in3 => \N__11977\,
            lcout => \DUT.uart_inst0.N_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_3_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011111110"
        )
    port map (
            in0 => \N__12162\,
            in1 => \N__11944\,
            in2 => \N__11926\,
            in3 => \N__11890\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12799\,
            ce => \N__12376\,
            sr => \_gnd_net_\
        );

    \ioFifoData_iobuf_RNO_2_LC_20_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12478\,
            lcout => \N_1241_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_RNIA7A5_4_LC_20_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12525\,
            in1 => \N__12543\,
            in2 => \N__12511\,
            in3 => \N__12558\,
            lcout => \DUT.uart_inst0.un1_tx_clk_divider_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_RNIHKCN_13_LC_20_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13089\,
            in2 => \_gnd_net_\,
            in3 => \N__13107\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.un1_tx_clk_divider_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_RNITC2S1_0_LC_20_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12454\,
            in1 => \N__12295\,
            in2 => \N__12448\,
            in3 => \N__12289\,
            lcout => \DUT.uart_inst0.un1_tx_clk_divider_0\,
            ltout => \DUT.uart_inst0.un1_tx_clk_divider_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNI5PJS2_1_LC_20_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111111111"
        )
    port map (
            in0 => \N__12283\,
            in1 => \_gnd_net_\,
            in2 => \N__12445\,
            in3 => \N__12438\,
            lcout => \DUT.uart_inst0.N_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_RNIQM95_0_LC_20_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12848\,
            in1 => \N__12612\,
            in2 => \N__12580\,
            in3 => \N__12594\,
            lcout => \DUT.uart_inst0.un1_tx_clk_divider_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_8_LC_20_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13143\,
            in1 => \N__13158\,
            in2 => \N__13128\,
            in3 => \N__12492\,
            lcout => \DUT.uart_inst0.un1_tx_clk_divider_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNI9B9Q2_1_LC_20_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12282\,
            in2 => \_gnd_net_\,
            in3 => \N__12196\,
            lcout => \DUT.uart_inst0.N_147\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_21_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12849\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_21_9_0_\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_1_LC_21_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12613\,
            in2 => \N__13042\,
            in3 => \N__12601\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_1\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_0\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_1\,
            clk => \N__12825\,
            ce => 'H',
            sr => \N__12637\
        );

    \DUT.uart_inst0.tx_clk_divider_2_LC_21_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13008\,
            in2 => \N__12598\,
            in3 => \N__12583\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_2\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_1\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_2\,
            clk => \N__12825\,
            ce => 'H',
            sr => \N__12637\
        );

    \DUT.uart_inst0.tx_clk_divider_3_LC_21_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12579\,
            in2 => \N__13043\,
            in3 => \N__12565\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_3\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_2\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_3\,
            clk => \N__12825\,
            ce => 'H',
            sr => \N__12637\
        );

    \DUT.uart_inst0.tx_clk_divider_4_LC_21_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13012\,
            in2 => \N__12562\,
            in3 => \N__12547\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_4\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_3\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_4\,
            clk => \N__12825\,
            ce => 'H',
            sr => \N__12637\
        );

    \DUT.uart_inst0.tx_clk_divider_5_LC_21_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12544\,
            in2 => \N__13044\,
            in3 => \N__12532\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_5\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_4\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_5\,
            clk => \N__12825\,
            ce => 'H',
            sr => \N__12637\
        );

    \DUT.uart_inst0.tx_clk_divider_6_LC_21_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13016\,
            in2 => \N__12529\,
            in3 => \N__12514\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_6\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_5\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_6\,
            clk => \N__12825\,
            ce => 'H',
            sr => \N__12637\
        );

    \DUT.uart_inst0.tx_clk_divider_7_LC_21_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12510\,
            in2 => \N__13045\,
            in3 => \N__12496\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_7\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_6\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_7\,
            clk => \N__12825\,
            ce => 'H',
            sr => \N__12637\
        );

    \DUT.uart_inst0.tx_clk_divider_8_LC_21_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12493\,
            in2 => \N__13004\,
            in3 => \N__12481\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_21_10_0_\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_8\,
            clk => \N__12821\,
            ce => 'H',
            sr => \N__12636\
        );

    \DUT.uart_inst0.tx_clk_divider_9_LC_21_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12972\,
            in2 => \N__13162\,
            in3 => \N__13147\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_9\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_8\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_9\,
            clk => \N__12821\,
            ce => 'H',
            sr => \N__12636\
        );

    \DUT.uart_inst0.tx_clk_divider_10_LC_21_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13144\,
            in2 => \N__13002\,
            in3 => \N__13132\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_10\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_9\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_10\,
            clk => \N__12821\,
            ce => 'H',
            sr => \N__12636\
        );

    \DUT.uart_inst0.tx_clk_divider_11_LC_21_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12965\,
            in2 => \N__13129\,
            in3 => \N__13111\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_11\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_10\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_11\,
            clk => \N__12821\,
            ce => 'H',
            sr => \N__12636\
        );

    \DUT.uart_inst0.tx_clk_divider_12_LC_21_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13108\,
            in2 => \N__13003\,
            in3 => \N__13096\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_12\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_11\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_12\,
            clk => \N__12821\,
            ce => 'H',
            sr => \N__12636\
        );

    \DUT.uart_inst0.tx_clk_divider_13_LC_21_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13090\,
            in2 => \_gnd_net_\,
            in3 => \N__13093\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12821\,
            ce => 'H',
            sr => \N__12636\
        );

    \DUT.uart_inst0.tx_clk_divider_0_LC_21_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12961\,
            in2 => \_gnd_net_\,
            in3 => \N__12850\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12821\,
            ce => 'H',
            sr => \N__12636\
        );
end \INTERFACE\;
