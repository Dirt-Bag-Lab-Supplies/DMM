-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Mar 28 2020 19:39:19

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    ioFifoData : out std_logic_vector(7 downto 0);
    P1A9 : out std_logic;
    P1A1 : in std_logic;
    P1A8 : out std_logic;
    oRx_n : out std_logic;
    P1A7 : out std_logic;
    P1A3 : out std_logic;
    iTxE_n : in std_logic;
    iRxF_n : in std_logic;
    iClk : in std_logic;
    P1A2 : out std_logic;
    BTN_N : in std_logic;
    BTN1 : in std_logic;
    oTx_n : out std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__13213\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13108\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13012\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12996\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12994\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12985\ : std_logic;
signal \N__12984\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12977\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12947\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12941\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12905\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12898\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12895\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12892\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12884\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12868\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12847\ : std_logic;
signal \N__12842\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12820\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12814\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12785\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12748\ : std_logic;
signal \N__12745\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12730\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12703\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12631\ : std_logic;
signal \N__12628\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12616\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12577\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12557\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12530\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12518\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12494\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12451\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12442\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12388\ : std_logic;
signal \N__12387\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12379\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12338\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12317\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12289\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12230\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12139\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12136\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12100\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11833\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11277\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10771\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10658\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10511\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10177\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9753\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9225\ : std_logic;
signal \N__9222\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8930\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8415\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8406\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8079\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8007\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7972\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7893\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7766\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7712\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7683\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7657\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7648\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7380\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7362\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7101\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6993\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6759\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6378\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6369\ : std_logic;
signal \N__6366\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5017\ : std_logic;
signal \wRamRdData_6\ : std_logic;
signal \wRamRdData_2\ : std_logic;
signal \wRamRdData_3\ : std_logic;
signal \wRamRdData_5\ : std_logic;
signal \BTN_N_c\ : std_logic;
signal \wRamRdData_7\ : std_logic;
signal \wRamRdData_0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \wRamRdData_4\ : std_logic;
signal \wRamRdData_1\ : std_logic;
signal \GNDG0\ : std_logic;
signal \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO\ : std_logic;
signal \DUT.fifo_rx_inst.N_86_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1\ : std_logic;
signal \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1_cascade_\ : std_logic;
signal \oTx_n_c_i\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_5\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_5\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_5\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_6\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_6\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_6\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_awe2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_awe2_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDataro_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDataro_2\ : std_logic;
signal \DUT.fifo_rx_inst.N_42\ : std_logic;
signal \DUT.fifo_rx_inst.rWritePtrZ0Z_0\ : std_logic;
signal \DUT.fifo_rx_inst.N_42_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rWritePtrZ0Z_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_awe1_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.un1_i11_i\ : std_logic;
signal \DUT.fifo_tx_inst.un1_i11_i_cascade_\ : std_logic;
signal \wRxBufferEmpty_i_0_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.un1_rFifoCount16_0_i_0\ : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoCount_RNIK3G92Z0Z_1\ : std_logic;
signal \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0\ : std_logic;
signal \DUT.fifo_rx_inst.un1_rFifoCount_1_axb_2\ : std_logic;
signal \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoCountZ0Z_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoCountZ0Z_1\ : std_logic;
signal \DUT.fifo_tx_inst.N_35_cascade_\ : std_logic;
signal \G_143_cascade_\ : std_logic;
signal \fifo_inst.ftdi_input_inst.SUMZ0Z_2_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.N_86\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram0_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram3_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram2_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_\ : std_logic;
signal \wRxBufferEmpty_i_0_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDataro_1\ : std_logic;
signal \DUT.fifo_rx_inst.rTxByte_42_0\ : std_logic;
signal \DUT.fifo_rx_inst.rTxByte_42_1_cascade_\ : std_logic;
signal \wRxBufferEmpty_i_0\ : std_logic;
signal \rFifoDatarff_0_RNIHJV05\ : std_logic;
signal \DUT.fifo_rx_inst.rReadPtrZ0Z_1\ : std_logic;
signal \DUT.fifo_rx_inst.rReadPtr_RNI4NC92Z0Z_0\ : std_logic;
signal \DUT.fifo_rx_inst.N_73\ : std_logic;
signal \DUT.fifo_rx_inst.rReadPtr_RNI4NC92Z0Z_0_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.rReadPtrZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.recv_state_srsts_1_0_6_cascade_\ : std_logic;
signal \DUT.fifo_rx_inst.un1_rFifoCount16_0_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoCountZ0Z_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_awe0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoDataro_0\ : std_logic;
signal \oTx_n_c\ : std_logic;
signal \P1A2_c\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoCountZ0Z_0\ : std_logic;
signal \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0\ : std_logic;
signal \bfn_14_19_0_\ : std_logic;
signal \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0\ : std_logic;
signal \DUT.fifo_tx_inst.N_35\ : std_logic;
signal \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoDataro_3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoDataro_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoDataro_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoDataro_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoDataror_1_0_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.un1_i11_2_i_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_3\ : std_logic;
signal \DUT.fifo_tx_inst.CO0\ : std_logic;
signal \DUT.fifo_tx_inst.CO0_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.un1_i11_2_i\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_7\ : std_logic;
signal \DUT.fifo_tx_inst.N_33\ : std_logic;
signal \DUT.fifo_tx_inst.N_41\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_2\ : std_logic;
signal \DUT.rFifoDatarx_2_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.N_40\ : std_logic;
signal \G_145_cascade_\ : std_logic;
signal \G_145\ : std_logic;
signal \G_142_cascade_\ : std_logic;
signal \G_144\ : std_logic;
signal \fifo_inst.ftdi_input_inst.SUMZ0Z_3\ : std_logic;
signal \G_147\ : std_logic;
signal \G_142\ : std_logic;
signal \G_141\ : std_logic;
signal \G_141_cascade_\ : std_logic;
signal \G_140\ : std_logic;
signal \fifo_inst_ftdi_input_inst_oTxFull_0\ : std_logic;
signal \G_140_cascade_\ : std_logic;
signal \G_143\ : std_logic;
signal \G_146\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_0\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_1\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_2\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_3\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_4\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_5\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_6\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_ram1_7\ : std_logic;
signal \DUT.fifo_rx_inst.rFifoData_awe1\ : std_logic;
signal \DUT.wRxByte_0\ : std_logic;
signal \DUT.wRxByte_1\ : std_logic;
signal \DUT.wRxByte_2\ : std_logic;
signal \DUT.wRxByte_3\ : std_logic;
signal \DUT.wRxByte_4\ : std_logic;
signal \DUT.wRxByte_5\ : std_logic;
signal \DUT.wRxByte_6\ : std_logic;
signal \DUT.wRxByte_7\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_2_cascade_\ : std_logic;
signal \DUT.wRcvd\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_8_i_o2_2_1_2_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_8_i_o2_2_2_cascade_\ : std_logic;
signal \DUT.uart_inst0.recv_state_RNO_0Z0Z_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.un1_m2_e_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_69\ : std_logic;
signal \DUT.uart_inst0.recv_state_RNITN8GJZ0Z_2_cascade_\ : std_logic;
signal \DUT.uart_inst0.recv_state_RNITN8GJZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remainingZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remainingZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remainingZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.rx_bits_remainingZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.N_98_4_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_m2_e_0\ : std_logic;
signal \DUT.uart_inst0.r_N_5_mux_cascade_\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.N_98_4\ : std_logic;
signal \DUT.uart_inst0.r_N_3_mux_cascade_\ : std_logic;
signal \DUT.uart_inst0.recv_N_5_mux\ : std_logic;
signal \DUT.uart_inst0.g3_cascade_\ : std_logic;
signal \DUT.uart_inst0.g3_1\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_0_c3\ : std_logic;
signal \DUT.uart_inst0.un1_m7_3\ : std_logic;
signal \DUT.uart_inst0.un1_tx_state_0_a4_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_s1_sn_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_7_1_0_3\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_RNO_0Z0Z_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.g0_i_o4_0_4_cascade_\ : std_logic;
signal \DUT.fifo_tx_inst.rWritePtrZ0Z_1\ : std_logic;
signal \DUT.fifo_tx_inst.rWritePtrZ0Z_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoCountZ0Z_2\ : std_logic;
signal \DUT.rFifoDatarxZ0Z_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4\ : std_logic;
signal \DUT.rFifoDatarx_4_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_data_RNO_0Z0Z_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram1_6\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram0_6\ : std_logic;
signal \DUT.fifo_tx_inst.rReadPtrZ0Z_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_data_RNO_0Z0Z_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_0\ : std_logic;
signal \rTxByteZ0Z_2\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_2\ : std_logic;
signal \rTxByteZ0Z_4\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_4\ : std_logic;
signal \rTxByteZ0Z_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_5\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_6\ : std_logic;
signal \rTxByteZ0Z_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_7\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_awe3\ : std_logic;
signal \DUT.rFifoDatarx_7\ : std_logic;
signal \G_152_cascade_\ : std_logic;
signal \G_151\ : std_logic;
signal \G_150\ : std_logic;
signal \fifo_inst.ftdi_input_inst.un1_rWrStateZ0Z_1\ : std_logic;
signal \G_149\ : std_logic;
signal \fifo_inst.ftdi_input_inst.un2_oPacketAvail_iZ0\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_10_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_RNIKU472Z0Z_10\ : std_logic;
signal \DUT.uart_inst0.recv_state_RNO_0Z0Z_0\ : std_logic;
signal \DUT.uart_inst0.recv_state_RNO_1Z0Z_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_10\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_2\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_8_i_o2_1_2_cascade_\ : std_logic;
signal \DUT.uart_inst0.recv_state_RNO_0Z0Z_4_cascade_\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_3\ : std_logic;
signal \P1A1_c\ : std_logic;
signal \DUT.uart_inst0.recv_stateZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.recv_state_srsts_1_5\ : std_logic;
signal \bfn_16_16_0_\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_s1_1\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_0_s1\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_1_s1_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_1_s1\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_s1_3\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_2_s1\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_3_s1\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_cry_4_s1\ : std_logic;
signal \DUT.uart_inst0.N_105\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.N_102\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ1Z_3\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_8_i_o2_1_1_2\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_s1_4\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_RNO_0Z0Z_2\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_8_i_o2_1_2\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_RNO_1Z0Z_2\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_8_i_o2_2_2\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_6_cascade_\ : std_logic;
signal \DUT.uart_inst0.un1_tx_bits_remaining_axbxc2_N_4L5_1_1\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.un1_tx_bits_remaining_axbxc2_N_4L5_1\ : std_logic;
signal \rRxReadZ0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoCountZ0Z_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoCount_RNIBPFMZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.g0_0_0_a3_3_cascade_\ : std_logic;
signal \DUT.uart_inst0.g0_0_0_a3_5_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_159_0_0\ : std_logic;
signal \DUT.N_37\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_0_1_5_cascade_\ : std_logic;
signal \DUT.uart_inst0.g0_i_o4_0_5\ : std_logic;
signal \DUT.uart_inst0.N_14_cascade_\ : std_logic;
signal \P1A7_c\ : std_logic;
signal \DUT.uart_inst0.N_6\ : std_logic;
signal \DUT.uart_inst0.un1_tx_bits_remaining_axbxc2_N_4L5_1_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_1\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_2\ : std_logic;
signal \DUT.rFifoDatarx_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_data_RNO_0Z0Z_1_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.tx_data_RNO_0Z0Z_0\ : std_logic;
signal \DUT.rFifoDatarx_5\ : std_logic;
signal \DUT.uart_inst0.tx_data_RNO_0Z0Z_5_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_5\ : std_logic;
signal \rTxByteZ0Z_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_1\ : std_logic;
signal \rTxByteZ0Z_0\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_0\ : std_logic;
signal \rTxByteZ0Z_6\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_6\ : std_logic;
signal \DUT.uart_inst0.tx_data_8_321_a2_0\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_11\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_12\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_9_cascade_\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_a_13\ : std_logic;
signal \DUT.uart_inst0.rx_countdown_3_s1_5\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.un2_rx_clk_divider_0\ : std_logic;
signal \DUT.uart_inst0.N_70\ : std_logic;
signal \DUT.uart_inst0.rx_countdownZ0Z_3\ : std_logic;
signal \G_148\ : std_logic;
signal \fifo_inst.ftdi_output_inst.N_95_cascade_\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_3\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2\ : std_logic;
signal \fifo_inst.ftdi_output_inst.N_95\ : std_logic;
signal \fifo_inst.ftdi_output_inst.m14_1_cascade_\ : std_logic;
signal \fifo_inst.ftdi_output_inst.N_86_0\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remaining_RNO_1Z0Z_2\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_9\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_8\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_7\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.tx_data_i_m_4_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.tx_countdown_0_c4_i\ : std_logic;
signal \DUT.uart_inst0.tx_state_ns_0_o3_1_0_1\ : std_logic;
signal \DUT.rFifoDatarx_6\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_7\ : std_logic;
signal \DUT.uart_inst0.tx_data_RNO_0Z0Z_6_cascade_\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_6\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_4\ : std_logic;
signal \DUT.rFifoDataror_0\ : std_logic;
signal \DUT.uart_inst0.tx_data_RNO_0Z0Z_3_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_152_0\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.N_159\ : std_logic;
signal \DUT.uart_inst0.tx_dataZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.g0_i_a4_0_4\ : std_logic;
signal \DUT.uart_inst0.tx_countdownZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.g0_i_a4_0_5_cascade_\ : std_logic;
signal \DUT.uart_inst0.N_15\ : std_logic;
signal \DUT.uart_inst0.N_7\ : std_logic;
signal \DUT.fifo_tx_inst.rReadPtrZ0Z_1\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram3_3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3\ : std_logic;
signal \DUT.rFifoDatarx_3\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remainingZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.tx_state_ns_i_i_a2_0_0_0_cascade_\ : std_logic;
signal \DUT.uart_inst0.g0_i_a4_1_0\ : std_logic;
signal \DUT.uart_inst0.d_N_5_mux\ : std_logic;
signal \rTxByteZ0Z_3\ : std_logic;
signal \DUT.fifo_tx_inst.rFifoData_ram2_3\ : std_logic;
signal \DUT.fifo_tx_inst.N_39\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rTxE_nZ0Z_1\ : std_logic;
signal \iTxE_n_c\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rTxE_nZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_1\ : std_logic;
signal \bfn_18_13_0_\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ1Z_1\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_0\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_1\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_2_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_2\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_3\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_4_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_4\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_6\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_5_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_5\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_7\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_6\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_7\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_8\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO\ : std_logic;
signal \bfn_18_14_0_\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_9\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_8\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_10\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_9\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_11\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_10\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_12\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_11\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_13\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_12\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_14\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_13\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_15\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_14\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_15\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_16\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO\ : std_logic;
signal \bfn_18_15_0_\ : std_logic;
signal \DUT.uart_inst0.N_72\ : std_logic;
signal \DUT.uart_inst0.rx_clk_divider_1_cry_16\ : std_logic;
signal \DUT.uart_inst0.rx_clk_dividerZ0Z_17\ : std_logic;
signal \fifo_inst.wRamRdAddr_2\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rWrDelayZ0\ : std_logic;
signal \fifo_inst.ftdi_output_inst.N_3_0\ : std_logic;
signal \fifo_inst.wRamRdAddr_0\ : std_logic;
signal \fifo_inst.ftdi_output_inst.N_3_0_cascade_\ : std_logic;
signal \fifo_inst.wRamRdAddr_1\ : std_logic;
signal \DUT.uart_inst0.tx_state_ns_i_i_a2_0_0_0\ : std_logic;
signal \DUT.uart_inst0.tx_state_0_sqmuxa_i_0\ : std_logic;
signal \wPllLocked_iso_i\ : std_logic;
signal \DUT.uart_inst0.N_345_0_0\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remaining_0_sqmuxa\ : std_logic;
signal \DUT.rTransmitZ0\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_0_sqmuxa\ : std_logic;
signal \wPllLocked\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_0_sqmuxa_cascade_\ : std_logic;
signal \DUT.uart_inst0.un1_tx_clk_divider_0\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rRxF_nZ0Z_1\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_0\ : std_logic;
signal \bfn_18_19_0_\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_0\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_1\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_3\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_2\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_4\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_3\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_5\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_4\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_6\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_5\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_7\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_6\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_7\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_8\ : std_logic;
signal \bfn_18_20_0_\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_9\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_8\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_10\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_9\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_11\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_10\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_12\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_11\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_cry_12\ : std_logic;
signal \DUT.uart_inst0.tx_clk_dividerZ0Z_13\ : std_logic;
signal \DUT.uart_inst0.tx_clk_divider_1_sqmuxa_1_i\ : std_logic;
signal \DUT.uart_inst0.tx_state_ns_i_i_0_0\ : std_logic;
signal \DUT.uart_inst0.N_345_0\ : std_logic;
signal \DUT.uart_inst0.tx_state_ns_i_i_a2_0_1_0\ : std_logic;
signal \DUT.tx_state_0\ : std_logic;
signal \wPllLocked_iso_i_g\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remainingZ0Z_2\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remainingZ0Z_0\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remaining_RNO_0Z0Z_3\ : std_logic;
signal \DUT.tx_state_1\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remainingZ0Z_1\ : std_logic;
signal \DUT.uart_inst0.tx_bits_remaining_RNO_0Z0Z_2\ : std_logic;
signal \iRxF_n_c\ : std_logic;
signal \fifo_inst.ftdi_output_inst.rRxF_nZ0Z_0\ : std_logic;
signal clk_48mhz : std_logic;
signal \wPllLocked_g\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \iClk_wire\ : std_logic;
signal \P1A8_wire\ : std_logic;
signal \ioFifoData_wire\ : std_logic_vector(7 downto 0);
signal \P1A9_wire\ : std_logic;
signal \oRx_n_wire\ : std_logic;
signal \P1A2_wire\ : std_logic;
signal \iRxF_n_wire\ : std_logic;
signal \P1A3_wire\ : std_logic;
signal \P1A7_wire\ : std_logic;
signal \BTN_N_wire\ : std_logic;
signal \oTx_n_wire\ : std_logic;
signal \iTxE_n_wire\ : std_logic;
signal \P1A1_wire\ : std_logic;
signal \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \top_pll_inst.top_pll_inst_pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \iClk_wire\ <= iClk;
    P1A8 <= \P1A8_wire\;
    ioFifoData <= \ioFifoData_wire\;
    P1A9 <= \P1A9_wire\;
    oRx_n <= \oRx_n_wire\;
    P1A2 <= \P1A2_wire\;
    \iRxF_n_wire\ <= iRxF_n;
    P1A3 <= \P1A3_wire\;
    P1A7 <= \P1A7_wire\;
    \BTN_N_wire\ <= BTN_N;
    oTx_n <= \oTx_n_wire\;
    \iTxE_n_wire\ <= iTxE_n;
    \P1A1_wire\ <= P1A1;
    \wRamRdData_7\ <= \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RDATA_wire\(14);
    \wRamRdData_6\ <= \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RDATA_wire\(12);
    \wRamRdData_5\ <= \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RDATA_wire\(10);
    \wRamRdData_4\ <= \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RDATA_wire\(8);
    \wRamRdData_3\ <= \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RDATA_wire\(6);
    \wRamRdData_2\ <= \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RDATA_wire\(4);
    \wRamRdData_1\ <= \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RDATA_wire\(2);
    \wRamRdData_0\ <= \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RDATA_wire\(0);
    \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__11068\&\N__10945\&\N__10975\;
    \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__7876\&\N__7855\&\N__7819\;
    \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \top_pll_inst.top_pll_inst_pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \fifo_inst.ftdi_input_inst.ram512x8_inst_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 1,
            READ_MODE => 1,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RDATA_wire\,
            RADDR => \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_RADDR_wire\,
            WADDR => \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_WADDR_wire\,
            MASK => \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_MASK_wire\,
            WDATA => \fifo_inst.ftdi_input_inst.ram512x8_inst_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \GNDG0\,
            RE => \N__13008\,
            WCLKE => 'H',
            WCLK => \N__12139\,
            WE => \N__6523\
        );

    \top_pll_inst.top_pll_inst_pll\ : PLL40
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "0111111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            PLLOUTGLOBAL => clk_48mhz,
            SDI => \GNDG0\,
            BYPASS => \GNDG0\,
            RESETB => \N__5137\,
            PLLOUTCORE => OPEN,
            LOCK => \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO\,
            SDO => OPEN,
            SCLK => \GNDG0\,
            LATCHINPUTVALUE => \GNDG0\,
            EXTFEEDBACK => \GNDG0\,
            DYNAMICDELAY => \top_pll_inst.top_pll_inst_pll_DYNAMICDELAY_wire\,
            PLLIN => \N__13213\
        );

    \top_pll_inst.top_pll_inst_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \VCCG0\,
            DIN => '0',
            DOUT => \N__13213\,
            PACKAGEPIN => \iClk_wire\
        );

    \P1A8_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13199\,
            DIN => \N__13198\,
            DOUT => \N__13197\,
            PACKAGEPIN => \P1A8_wire\
        );

    \P1A8_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13199\,
            PADOUT => \N__13198\,
            PADIN => \N__13197\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13190\,
            DIN => \N__13189\,
            DOUT => \N__13188\,
            PACKAGEPIN => \ioFifoData_wire\(1)
        );

    \ioFifoData_obuft_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13190\,
            PADOUT => \N__13189\,
            PADIN => \N__13188\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5229\,
            DIN0 => OPEN,
            DOUT0 => \N__5161\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A9_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13181\,
            DIN => \N__13180\,
            DOUT => \N__13179\,
            PACKAGEPIN => \P1A9_wire\
        );

    \P1A9_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13181\,
            PADOUT => \N__13180\,
            PADIN => \N__13179\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13172\,
            DIN => \N__13171\,
            DOUT => \N__13170\,
            PACKAGEPIN => \ioFifoData_wire\(4)
        );

    \ioFifoData_obuft_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13172\,
            PADOUT => \N__13171\,
            PADIN => \N__13170\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5243\,
            DIN0 => OPEN,
            DOUT0 => \N__5086\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13163\,
            DIN => \N__13162\,
            DOUT => \N__13161\,
            PACKAGEPIN => \ioFifoData_wire\(0)
        );

    \ioFifoData_obuft_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13163\,
            PADOUT => \N__13162\,
            PADIN => \N__13161\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5216\,
            DIN0 => OPEN,
            DOUT0 => \N__5107\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \oRx_n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13154\,
            DIN => \N__13153\,
            DOUT => \N__13152\,
            PACKAGEPIN => \oRx_n_wire\
        );

    \oRx_n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13154\,
            PADOUT => \N__13153\,
            PADIN => \N__13152\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__13018\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13145\,
            DIN => \N__13144\,
            DOUT => \N__13143\,
            PACKAGEPIN => \P1A2_wire\
        );

    \P1A2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13145\,
            PADOUT => \N__13144\,
            PADIN => \N__13143\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6181\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13136\,
            DIN => \N__13135\,
            DOUT => \N__13134\,
            PACKAGEPIN => \ioFifoData_wire\(7)
        );

    \ioFifoData_obuft_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13136\,
            PADOUT => \N__13135\,
            PADIN => \N__13134\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5215\,
            DIN0 => OPEN,
            DOUT0 => \N__5122\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \iRxF_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13127\,
            DIN => \N__13126\,
            DOUT => \N__13125\,
            PACKAGEPIN => \iRxF_n_wire\
        );

    \iRxF_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13127\,
            PADOUT => \N__13126\,
            PADIN => \N__13125\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \iRxF_n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13118\,
            DIN => \N__13117\,
            DOUT => \N__13116\,
            PACKAGEPIN => \P1A3_wire\
        );

    \P1A3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13118\,
            PADOUT => \N__13117\,
            PADIN => \N__13116\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A7_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13109\,
            DIN => \N__13108\,
            DOUT => \N__13107\,
            PACKAGEPIN => \P1A7_wire\
        );

    \P1A7_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13109\,
            PADOUT => \N__13108\,
            PADIN => \N__13107\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8809\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BTN_N_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13100\,
            DIN => \N__13099\,
            DOUT => \N__13098\,
            PACKAGEPIN => \BTN_N_wire\
        );

    \BTN_N_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13100\,
            PADOUT => \N__13099\,
            PADIN => \N__13098\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \BTN_N_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13091\,
            DIN => \N__13090\,
            DOUT => \N__13089\,
            PACKAGEPIN => \ioFifoData_wire\(3)
        );

    \ioFifoData_obuft_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13091\,
            PADOUT => \N__13090\,
            PADIN => \N__13089\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5250\,
            DIN0 => OPEN,
            DOUT0 => \N__5044\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13082\,
            DIN => \N__13081\,
            DOUT => \N__13080\,
            PACKAGEPIN => \ioFifoData_wire\(6)
        );

    \ioFifoData_obuft_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13082\,
            PADOUT => \N__13081\,
            PADIN => \N__13080\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5214\,
            DIN0 => OPEN,
            DOUT0 => \N__5074\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13073\,
            DIN => \N__13072\,
            DOUT => \N__13071\,
            PACKAGEPIN => \ioFifoData_wire\(5)
        );

    \ioFifoData_obuft_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13073\,
            PADOUT => \N__13072\,
            PADIN => \N__13071\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5242\,
            DIN0 => OPEN,
            DOUT0 => \N__5026\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \oTx_n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13064\,
            DIN => \N__13063\,
            DOUT => \N__13062\,
            PACKAGEPIN => \oTx_n_wire\
        );

    \oTx_n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13064\,
            PADOUT => \N__13063\,
            PADIN => \N__13062\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6214\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \iTxE_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13055\,
            DIN => \N__13054\,
            DOUT => \N__13053\,
            PACKAGEPIN => \iTxE_n_wire\
        );

    \iTxE_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13055\,
            PADOUT => \N__13054\,
            PADIN => \N__13053\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \iTxE_n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ioFifoData_obuft_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13046\,
            DIN => \N__13045\,
            DOUT => \N__13044\,
            PACKAGEPIN => \ioFifoData_wire\(2)
        );

    \ioFifoData_obuft_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13046\,
            PADOUT => \N__13045\,
            PADIN => \N__13044\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5251\,
            DIN0 => OPEN,
            DOUT0 => \N__5062\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \P1A1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13037\,
            DIN => \N__13036\,
            DOUT => \N__13035\,
            PACKAGEPIN => \P1A1_wire\
        );

    \P1A1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13037\,
            PADOUT => \N__13036\,
            PADIN => \N__13035\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \P1A1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__3084\ : IoInMux
    port map (
            O => \N__13018\,
            I => \N__13015\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__13015\,
            I => \N__13012\
        );

    \I__3082\ : IoSpan4Mux
    port map (
            O => \N__13012\,
            I => \N__13009\
        );

    \I__3081\ : Span4Mux_s3_v
    port map (
            O => \N__13009\,
            I => \N__13005\
        );

    \I__3080\ : SRMux
    port map (
            O => \N__13008\,
            I => \N__13002\
        );

    \I__3079\ : Span4Mux_v
    port map (
            O => \N__13005\,
            I => \N__12972\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__13002\,
            I => \N__12972\
        );

    \I__3077\ : InMux
    port map (
            O => \N__13001\,
            I => \N__12967\
        );

    \I__3076\ : InMux
    port map (
            O => \N__13000\,
            I => \N__12967\
        );

    \I__3075\ : InMux
    port map (
            O => \N__12999\,
            I => \N__12960\
        );

    \I__3074\ : InMux
    port map (
            O => \N__12998\,
            I => \N__12960\
        );

    \I__3073\ : InMux
    port map (
            O => \N__12997\,
            I => \N__12960\
        );

    \I__3072\ : CascadeMux
    port map (
            O => \N__12996\,
            I => \N__12957\
        );

    \I__3071\ : CascadeMux
    port map (
            O => \N__12995\,
            I => \N__12954\
        );

    \I__3070\ : CascadeMux
    port map (
            O => \N__12994\,
            I => \N__12951\
        );

    \I__3069\ : CascadeMux
    port map (
            O => \N__12993\,
            I => \N__12948\
        );

    \I__3068\ : CascadeMux
    port map (
            O => \N__12992\,
            I => \N__12944\
        );

    \I__3067\ : CascadeMux
    port map (
            O => \N__12991\,
            I => \N__12941\
        );

    \I__3066\ : CascadeMux
    port map (
            O => \N__12990\,
            I => \N__12938\
        );

    \I__3065\ : CascadeMux
    port map (
            O => \N__12989\,
            I => \N__12935\
        );

    \I__3064\ : CascadeMux
    port map (
            O => \N__12988\,
            I => \N__12932\
        );

    \I__3063\ : CascadeMux
    port map (
            O => \N__12987\,
            I => \N__12929\
        );

    \I__3062\ : CascadeMux
    port map (
            O => \N__12986\,
            I => \N__12926\
        );

    \I__3061\ : CascadeMux
    port map (
            O => \N__12985\,
            I => \N__12923\
        );

    \I__3060\ : CascadeMux
    port map (
            O => \N__12984\,
            I => \N__12920\
        );

    \I__3059\ : CascadeMux
    port map (
            O => \N__12983\,
            I => \N__12917\
        );

    \I__3058\ : CascadeMux
    port map (
            O => \N__12982\,
            I => \N__12914\
        );

    \I__3057\ : CascadeMux
    port map (
            O => \N__12981\,
            I => \N__12911\
        );

    \I__3056\ : CascadeMux
    port map (
            O => \N__12980\,
            I => \N__12908\
        );

    \I__3055\ : CascadeMux
    port map (
            O => \N__12979\,
            I => \N__12905\
        );

    \I__3054\ : CascadeMux
    port map (
            O => \N__12978\,
            I => \N__12902\
        );

    \I__3053\ : CascadeMux
    port map (
            O => \N__12977\,
            I => \N__12899\
        );

    \I__3052\ : Span4Mux_v
    port map (
            O => \N__12972\,
            I => \N__12889\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__12967\,
            I => \N__12884\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__12960\,
            I => \N__12884\
        );

    \I__3049\ : InMux
    port map (
            O => \N__12957\,
            I => \N__12879\
        );

    \I__3048\ : InMux
    port map (
            O => \N__12954\,
            I => \N__12879\
        );

    \I__3047\ : InMux
    port map (
            O => \N__12951\,
            I => \N__12868\
        );

    \I__3046\ : InMux
    port map (
            O => \N__12948\,
            I => \N__12868\
        );

    \I__3045\ : InMux
    port map (
            O => \N__12947\,
            I => \N__12868\
        );

    \I__3044\ : InMux
    port map (
            O => \N__12944\,
            I => \N__12868\
        );

    \I__3043\ : InMux
    port map (
            O => \N__12941\,
            I => \N__12868\
        );

    \I__3042\ : InMux
    port map (
            O => \N__12938\,
            I => \N__12859\
        );

    \I__3041\ : InMux
    port map (
            O => \N__12935\,
            I => \N__12859\
        );

    \I__3040\ : InMux
    port map (
            O => \N__12932\,
            I => \N__12859\
        );

    \I__3039\ : InMux
    port map (
            O => \N__12929\,
            I => \N__12859\
        );

    \I__3038\ : InMux
    port map (
            O => \N__12926\,
            I => \N__12850\
        );

    \I__3037\ : InMux
    port map (
            O => \N__12923\,
            I => \N__12850\
        );

    \I__3036\ : InMux
    port map (
            O => \N__12920\,
            I => \N__12850\
        );

    \I__3035\ : InMux
    port map (
            O => \N__12917\,
            I => \N__12850\
        );

    \I__3034\ : InMux
    port map (
            O => \N__12914\,
            I => \N__12847\
        );

    \I__3033\ : InMux
    port map (
            O => \N__12911\,
            I => \N__12842\
        );

    \I__3032\ : InMux
    port map (
            O => \N__12908\,
            I => \N__12842\
        );

    \I__3031\ : InMux
    port map (
            O => \N__12905\,
            I => \N__12835\
        );

    \I__3030\ : InMux
    port map (
            O => \N__12902\,
            I => \N__12835\
        );

    \I__3029\ : InMux
    port map (
            O => \N__12899\,
            I => \N__12835\
        );

    \I__3028\ : CascadeMux
    port map (
            O => \N__12898\,
            I => \N__12832\
        );

    \I__3027\ : CascadeMux
    port map (
            O => \N__12897\,
            I => \N__12829\
        );

    \I__3026\ : CascadeMux
    port map (
            O => \N__12896\,
            I => \N__12826\
        );

    \I__3025\ : CascadeMux
    port map (
            O => \N__12895\,
            I => \N__12823\
        );

    \I__3024\ : CascadeMux
    port map (
            O => \N__12894\,
            I => \N__12820\
        );

    \I__3023\ : CascadeMux
    port map (
            O => \N__12893\,
            I => \N__12817\
        );

    \I__3022\ : CascadeMux
    port map (
            O => \N__12892\,
            I => \N__12814\
        );

    \I__3021\ : Span4Mux_v
    port map (
            O => \N__12889\,
            I => \N__12811\
        );

    \I__3020\ : Span4Mux_v
    port map (
            O => \N__12884\,
            I => \N__12808\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__12879\,
            I => \N__12799\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__12868\,
            I => \N__12799\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__12859\,
            I => \N__12799\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__12850\,
            I => \N__12799\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__12847\,
            I => \N__12792\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__12842\,
            I => \N__12792\
        );

    \I__3013\ : LocalMux
    port map (
            O => \N__12835\,
            I => \N__12792\
        );

    \I__3012\ : InMux
    port map (
            O => \N__12832\,
            I => \N__12785\
        );

    \I__3011\ : InMux
    port map (
            O => \N__12829\,
            I => \N__12785\
        );

    \I__3010\ : InMux
    port map (
            O => \N__12826\,
            I => \N__12785\
        );

    \I__3009\ : InMux
    port map (
            O => \N__12823\,
            I => \N__12776\
        );

    \I__3008\ : InMux
    port map (
            O => \N__12820\,
            I => \N__12776\
        );

    \I__3007\ : InMux
    port map (
            O => \N__12817\,
            I => \N__12776\
        );

    \I__3006\ : InMux
    port map (
            O => \N__12814\,
            I => \N__12776\
        );

    \I__3005\ : Odrv4
    port map (
            O => \N__12811\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3004\ : Odrv4
    port map (
            O => \N__12808\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3003\ : Odrv12
    port map (
            O => \N__12799\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3002\ : Odrv12
    port map (
            O => \N__12792\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__12785\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__12776\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2999\ : InMux
    port map (
            O => \N__12763\,
            I => \N__12759\
        );

    \I__2998\ : InMux
    port map (
            O => \N__12762\,
            I => \N__12756\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__12759\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_12\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__12756\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_12\
        );

    \I__2995\ : InMux
    port map (
            O => \N__12751\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_11\
        );

    \I__2994\ : InMux
    port map (
            O => \N__12748\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_12\
        );

    \I__2993\ : CascadeMux
    port map (
            O => \N__12745\,
            I => \N__12741\
        );

    \I__2992\ : InMux
    port map (
            O => \N__12744\,
            I => \N__12738\
        );

    \I__2991\ : InMux
    port map (
            O => \N__12741\,
            I => \N__12735\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__12738\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_13\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__12735\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_13\
        );

    \I__2988\ : SRMux
    port map (
            O => \N__12730\,
            I => \N__12726\
        );

    \I__2987\ : SRMux
    port map (
            O => \N__12729\,
            I => \N__12723\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__12726\,
            I => \N__12720\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__12723\,
            I => \N__12717\
        );

    \I__2984\ : Span4Mux_h
    port map (
            O => \N__12720\,
            I => \N__12711\
        );

    \I__2983\ : Span4Mux_h
    port map (
            O => \N__12717\,
            I => \N__12711\
        );

    \I__2982\ : SRMux
    port map (
            O => \N__12716\,
            I => \N__12708\
        );

    \I__2981\ : Odrv4
    port map (
            O => \N__12711\,
            I => \DUT.uart_inst0.tx_clk_divider_1_sqmuxa_1_i\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__12708\,
            I => \DUT.uart_inst0.tx_clk_divider_1_sqmuxa_1_i\
        );

    \I__2979\ : InMux
    port map (
            O => \N__12703\,
            I => \N__12700\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__12700\,
            I => \DUT.uart_inst0.tx_state_ns_i_i_0_0\
        );

    \I__2977\ : InMux
    port map (
            O => \N__12697\,
            I => \N__12694\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__12694\,
            I => \N__12690\
        );

    \I__2975\ : InMux
    port map (
            O => \N__12693\,
            I => \N__12687\
        );

    \I__2974\ : Odrv4
    port map (
            O => \N__12690\,
            I => \DUT.uart_inst0.N_345_0\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__12687\,
            I => \DUT.uart_inst0.N_345_0\
        );

    \I__2972\ : InMux
    port map (
            O => \N__12682\,
            I => \N__12679\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__12679\,
            I => \DUT.uart_inst0.tx_state_ns_i_i_a2_0_1_0\
        );

    \I__2970\ : CascadeMux
    port map (
            O => \N__12676\,
            I => \N__12667\
        );

    \I__2969\ : CascadeMux
    port map (
            O => \N__12675\,
            I => \N__12663\
        );

    \I__2968\ : InMux
    port map (
            O => \N__12674\,
            I => \N__12659\
        );

    \I__2967\ : CascadeMux
    port map (
            O => \N__12673\,
            I => \N__12656\
        );

    \I__2966\ : InMux
    port map (
            O => \N__12672\,
            I => \N__12650\
        );

    \I__2965\ : CascadeMux
    port map (
            O => \N__12671\,
            I => \N__12647\
        );

    \I__2964\ : InMux
    port map (
            O => \N__12670\,
            I => \N__12642\
        );

    \I__2963\ : InMux
    port map (
            O => \N__12667\,
            I => \N__12639\
        );

    \I__2962\ : InMux
    port map (
            O => \N__12666\,
            I => \N__12636\
        );

    \I__2961\ : InMux
    port map (
            O => \N__12663\,
            I => \N__12631\
        );

    \I__2960\ : InMux
    port map (
            O => \N__12662\,
            I => \N__12631\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__12659\,
            I => \N__12628\
        );

    \I__2958\ : InMux
    port map (
            O => \N__12656\,
            I => \N__12625\
        );

    \I__2957\ : InMux
    port map (
            O => \N__12655\,
            I => \N__12620\
        );

    \I__2956\ : InMux
    port map (
            O => \N__12654\,
            I => \N__12620\
        );

    \I__2955\ : InMux
    port map (
            O => \N__12653\,
            I => \N__12611\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__12650\,
            I => \N__12608\
        );

    \I__2953\ : InMux
    port map (
            O => \N__12647\,
            I => \N__12601\
        );

    \I__2952\ : InMux
    port map (
            O => \N__12646\,
            I => \N__12601\
        );

    \I__2951\ : InMux
    port map (
            O => \N__12645\,
            I => \N__12601\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__12642\,
            I => \N__12592\
        );

    \I__2949\ : LocalMux
    port map (
            O => \N__12639\,
            I => \N__12592\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__12636\,
            I => \N__12592\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__12631\,
            I => \N__12592\
        );

    \I__2946\ : Span4Mux_v
    port map (
            O => \N__12628\,
            I => \N__12584\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__12625\,
            I => \N__12584\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__12620\,
            I => \N__12584\
        );

    \I__2943\ : InMux
    port map (
            O => \N__12619\,
            I => \N__12577\
        );

    \I__2942\ : InMux
    port map (
            O => \N__12618\,
            I => \N__12577\
        );

    \I__2941\ : InMux
    port map (
            O => \N__12617\,
            I => \N__12577\
        );

    \I__2940\ : InMux
    port map (
            O => \N__12616\,
            I => \N__12570\
        );

    \I__2939\ : InMux
    port map (
            O => \N__12615\,
            I => \N__12570\
        );

    \I__2938\ : InMux
    port map (
            O => \N__12614\,
            I => \N__12570\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__12611\,
            I => \N__12567\
        );

    \I__2936\ : Span4Mux_v
    port map (
            O => \N__12608\,
            I => \N__12560\
        );

    \I__2935\ : LocalMux
    port map (
            O => \N__12601\,
            I => \N__12560\
        );

    \I__2934\ : Span4Mux_v
    port map (
            O => \N__12592\,
            I => \N__12560\
        );

    \I__2933\ : InMux
    port map (
            O => \N__12591\,
            I => \N__12557\
        );

    \I__2932\ : Span4Mux_h
    port map (
            O => \N__12584\,
            I => \N__12554\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__12577\,
            I => \DUT.tx_state_0\
        );

    \I__2930\ : LocalMux
    port map (
            O => \N__12570\,
            I => \DUT.tx_state_0\
        );

    \I__2929\ : Odrv4
    port map (
            O => \N__12567\,
            I => \DUT.tx_state_0\
        );

    \I__2928\ : Odrv4
    port map (
            O => \N__12560\,
            I => \DUT.tx_state_0\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__12557\,
            I => \DUT.tx_state_0\
        );

    \I__2926\ : Odrv4
    port map (
            O => \N__12554\,
            I => \DUT.tx_state_0\
        );

    \I__2925\ : CascadeMux
    port map (
            O => \N__12541\,
            I => \N__12536\
        );

    \I__2924\ : CascadeMux
    port map (
            O => \N__12540\,
            I => \N__12531\
        );

    \I__2923\ : InMux
    port map (
            O => \N__12539\,
            I => \N__12521\
        );

    \I__2922\ : InMux
    port map (
            O => \N__12536\,
            I => \N__12521\
        );

    \I__2921\ : InMux
    port map (
            O => \N__12535\,
            I => \N__12521\
        );

    \I__2920\ : InMux
    port map (
            O => \N__12534\,
            I => \N__12518\
        );

    \I__2919\ : InMux
    port map (
            O => \N__12531\,
            I => \N__12513\
        );

    \I__2918\ : InMux
    port map (
            O => \N__12530\,
            I => \N__12513\
        );

    \I__2917\ : InMux
    port map (
            O => \N__12529\,
            I => \N__12508\
        );

    \I__2916\ : InMux
    port map (
            O => \N__12528\,
            I => \N__12508\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__12521\,
            I => \N__12505\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__12518\,
            I => \N__12502\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__12513\,
            I => \N__12499\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__12508\,
            I => \N__12496\
        );

    \I__2911\ : Glb2LocalMux
    port map (
            O => \N__12505\,
            I => \N__12451\
        );

    \I__2910\ : Glb2LocalMux
    port map (
            O => \N__12502\,
            I => \N__12451\
        );

    \I__2909\ : Glb2LocalMux
    port map (
            O => \N__12499\,
            I => \N__12451\
        );

    \I__2908\ : Glb2LocalMux
    port map (
            O => \N__12496\,
            I => \N__12451\
        );

    \I__2907\ : SRMux
    port map (
            O => \N__12495\,
            I => \N__12451\
        );

    \I__2906\ : SRMux
    port map (
            O => \N__12494\,
            I => \N__12451\
        );

    \I__2905\ : SRMux
    port map (
            O => \N__12493\,
            I => \N__12451\
        );

    \I__2904\ : SRMux
    port map (
            O => \N__12492\,
            I => \N__12451\
        );

    \I__2903\ : SRMux
    port map (
            O => \N__12491\,
            I => \N__12451\
        );

    \I__2902\ : SRMux
    port map (
            O => \N__12490\,
            I => \N__12451\
        );

    \I__2901\ : SRMux
    port map (
            O => \N__12489\,
            I => \N__12451\
        );

    \I__2900\ : SRMux
    port map (
            O => \N__12488\,
            I => \N__12451\
        );

    \I__2899\ : SRMux
    port map (
            O => \N__12487\,
            I => \N__12451\
        );

    \I__2898\ : SRMux
    port map (
            O => \N__12486\,
            I => \N__12451\
        );

    \I__2897\ : SRMux
    port map (
            O => \N__12485\,
            I => \N__12451\
        );

    \I__2896\ : SRMux
    port map (
            O => \N__12484\,
            I => \N__12451\
        );

    \I__2895\ : GlobalMux
    port map (
            O => \N__12451\,
            I => \N__12448\
        );

    \I__2894\ : gio2CtrlBuf
    port map (
            O => \N__12448\,
            I => \wPllLocked_iso_i_g\
        );

    \I__2893\ : InMux
    port map (
            O => \N__12445\,
            I => \N__12439\
        );

    \I__2892\ : InMux
    port map (
            O => \N__12444\,
            I => \N__12436\
        );

    \I__2891\ : InMux
    port map (
            O => \N__12443\,
            I => \N__12432\
        );

    \I__2890\ : InMux
    port map (
            O => \N__12442\,
            I => \N__12429\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__12439\,
            I => \N__12426\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__12436\,
            I => \N__12423\
        );

    \I__2887\ : InMux
    port map (
            O => \N__12435\,
            I => \N__12420\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__12432\,
            I => \N__12417\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__12429\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_2\
        );

    \I__2884\ : Odrv4
    port map (
            O => \N__12426\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_2\
        );

    \I__2883\ : Odrv4
    port map (
            O => \N__12423\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_2\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__12420\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_2\
        );

    \I__2881\ : Odrv4
    port map (
            O => \N__12417\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_2\
        );

    \I__2880\ : InMux
    port map (
            O => \N__12406\,
            I => \N__12401\
        );

    \I__2879\ : CascadeMux
    port map (
            O => \N__12405\,
            I => \N__12397\
        );

    \I__2878\ : InMux
    port map (
            O => \N__12404\,
            I => \N__12393\
        );

    \I__2877\ : LocalMux
    port map (
            O => \N__12401\,
            I => \N__12390\
        );

    \I__2876\ : InMux
    port map (
            O => \N__12400\,
            I => \N__12384\
        );

    \I__2875\ : InMux
    port map (
            O => \N__12397\,
            I => \N__12379\
        );

    \I__2874\ : InMux
    port map (
            O => \N__12396\,
            I => \N__12379\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__12393\,
            I => \N__12376\
        );

    \I__2872\ : Span4Mux_v
    port map (
            O => \N__12390\,
            I => \N__12373\
        );

    \I__2871\ : InMux
    port map (
            O => \N__12389\,
            I => \N__12370\
        );

    \I__2870\ : InMux
    port map (
            O => \N__12388\,
            I => \N__12365\
        );

    \I__2869\ : InMux
    port map (
            O => \N__12387\,
            I => \N__12365\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__12384\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_0\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__12379\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_0\
        );

    \I__2866\ : Odrv12
    port map (
            O => \N__12376\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_0\
        );

    \I__2865\ : Odrv4
    port map (
            O => \N__12373\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_0\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__12370\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_0\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__12365\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_0\
        );

    \I__2862\ : CascadeMux
    port map (
            O => \N__12352\,
            I => \N__12349\
        );

    \I__2861\ : InMux
    port map (
            O => \N__12349\,
            I => \N__12346\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__12346\,
            I => \N__12343\
        );

    \I__2859\ : Odrv4
    port map (
            O => \N__12343\,
            I => \DUT.uart_inst0.tx_bits_remaining_RNO_0Z0Z_3\
        );

    \I__2858\ : InMux
    port map (
            O => \N__12340\,
            I => \N__12334\
        );

    \I__2857\ : InMux
    port map (
            O => \N__12339\,
            I => \N__12329\
        );

    \I__2856\ : InMux
    port map (
            O => \N__12338\,
            I => \N__12329\
        );

    \I__2855\ : CascadeMux
    port map (
            O => \N__12337\,
            I => \N__12325\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__12334\,
            I => \N__12312\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__12329\,
            I => \N__12312\
        );

    \I__2852\ : InMux
    port map (
            O => \N__12328\,
            I => \N__12307\
        );

    \I__2851\ : InMux
    port map (
            O => \N__12325\,
            I => \N__12307\
        );

    \I__2850\ : InMux
    port map (
            O => \N__12324\,
            I => \N__12304\
        );

    \I__2849\ : InMux
    port map (
            O => \N__12323\,
            I => \N__12299\
        );

    \I__2848\ : InMux
    port map (
            O => \N__12322\,
            I => \N__12299\
        );

    \I__2847\ : InMux
    port map (
            O => \N__12321\,
            I => \N__12296\
        );

    \I__2846\ : InMux
    port map (
            O => \N__12320\,
            I => \N__12289\
        );

    \I__2845\ : InMux
    port map (
            O => \N__12319\,
            I => \N__12289\
        );

    \I__2844\ : InMux
    port map (
            O => \N__12318\,
            I => \N__12289\
        );

    \I__2843\ : InMux
    port map (
            O => \N__12317\,
            I => \N__12286\
        );

    \I__2842\ : Span4Mux_v
    port map (
            O => \N__12312\,
            I => \N__12283\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__12307\,
            I => \N__12278\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__12304\,
            I => \N__12278\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__12299\,
            I => \N__12275\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__12296\,
            I => \N__12270\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__12289\,
            I => \N__12270\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__12286\,
            I => \N__12267\
        );

    \I__2835\ : Span4Mux_h
    port map (
            O => \N__12283\,
            I => \N__12262\
        );

    \I__2834\ : Span4Mux_v
    port map (
            O => \N__12278\,
            I => \N__12259\
        );

    \I__2833\ : Span4Mux_h
    port map (
            O => \N__12275\,
            I => \N__12256\
        );

    \I__2832\ : Span4Mux_v
    port map (
            O => \N__12270\,
            I => \N__12251\
        );

    \I__2831\ : Span4Mux_h
    port map (
            O => \N__12267\,
            I => \N__12251\
        );

    \I__2830\ : InMux
    port map (
            O => \N__12266\,
            I => \N__12246\
        );

    \I__2829\ : InMux
    port map (
            O => \N__12265\,
            I => \N__12246\
        );

    \I__2828\ : Odrv4
    port map (
            O => \N__12262\,
            I => \DUT.tx_state_1\
        );

    \I__2827\ : Odrv4
    port map (
            O => \N__12259\,
            I => \DUT.tx_state_1\
        );

    \I__2826\ : Odrv4
    port map (
            O => \N__12256\,
            I => \DUT.tx_state_1\
        );

    \I__2825\ : Odrv4
    port map (
            O => \N__12251\,
            I => \DUT.tx_state_1\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__12246\,
            I => \DUT.tx_state_1\
        );

    \I__2823\ : InMux
    port map (
            O => \N__12235\,
            I => \N__12230\
        );

    \I__2822\ : InMux
    port map (
            O => \N__12234\,
            I => \N__12225\
        );

    \I__2821\ : InMux
    port map (
            O => \N__12233\,
            I => \N__12225\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__12230\,
            I => \N__12218\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__12225\,
            I => \N__12218\
        );

    \I__2818\ : InMux
    port map (
            O => \N__12224\,
            I => \N__12213\
        );

    \I__2817\ : InMux
    port map (
            O => \N__12223\,
            I => \N__12210\
        );

    \I__2816\ : Span4Mux_v
    port map (
            O => \N__12218\,
            I => \N__12207\
        );

    \I__2815\ : InMux
    port map (
            O => \N__12217\,
            I => \N__12204\
        );

    \I__2814\ : InMux
    port map (
            O => \N__12216\,
            I => \N__12201\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__12213\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_1\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__12210\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_1\
        );

    \I__2811\ : Odrv4
    port map (
            O => \N__12207\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_1\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__12204\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_1\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__12201\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_1\
        );

    \I__2808\ : CascadeMux
    port map (
            O => \N__12190\,
            I => \N__12187\
        );

    \I__2807\ : InMux
    port map (
            O => \N__12187\,
            I => \N__12184\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__12184\,
            I => \N__12181\
        );

    \I__2805\ : Span4Mux_h
    port map (
            O => \N__12181\,
            I => \N__12178\
        );

    \I__2804\ : Odrv4
    port map (
            O => \N__12178\,
            I => \DUT.uart_inst0.tx_bits_remaining_RNO_0Z0Z_2\
        );

    \I__2803\ : InMux
    port map (
            O => \N__12175\,
            I => \N__12172\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__12172\,
            I => \N__12169\
        );

    \I__2801\ : Odrv12
    port map (
            O => \N__12169\,
            I => \iRxF_n_c\
        );

    \I__2800\ : CascadeMux
    port map (
            O => \N__12166\,
            I => \N__12161\
        );

    \I__2799\ : InMux
    port map (
            O => \N__12165\,
            I => \N__12158\
        );

    \I__2798\ : InMux
    port map (
            O => \N__12164\,
            I => \N__12155\
        );

    \I__2797\ : InMux
    port map (
            O => \N__12161\,
            I => \N__12152\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__12158\,
            I => \N__12147\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__12155\,
            I => \N__12147\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__12152\,
            I => \N__12142\
        );

    \I__2793\ : Sp12to4
    port map (
            O => \N__12147\,
            I => \N__12142\
        );

    \I__2792\ : Odrv12
    port map (
            O => \N__12142\,
            I => \fifo_inst.ftdi_output_inst.rRxF_nZ0Z_0\
        );

    \I__2791\ : ClkMux
    port map (
            O => \N__12139\,
            I => \N__11944\
        );

    \I__2790\ : ClkMux
    port map (
            O => \N__12138\,
            I => \N__11944\
        );

    \I__2789\ : ClkMux
    port map (
            O => \N__12137\,
            I => \N__11944\
        );

    \I__2788\ : ClkMux
    port map (
            O => \N__12136\,
            I => \N__11944\
        );

    \I__2787\ : ClkMux
    port map (
            O => \N__12135\,
            I => \N__11944\
        );

    \I__2786\ : ClkMux
    port map (
            O => \N__12134\,
            I => \N__11944\
        );

    \I__2785\ : ClkMux
    port map (
            O => \N__12133\,
            I => \N__11944\
        );

    \I__2784\ : ClkMux
    port map (
            O => \N__12132\,
            I => \N__11944\
        );

    \I__2783\ : ClkMux
    port map (
            O => \N__12131\,
            I => \N__11944\
        );

    \I__2782\ : ClkMux
    port map (
            O => \N__12130\,
            I => \N__11944\
        );

    \I__2781\ : ClkMux
    port map (
            O => \N__12129\,
            I => \N__11944\
        );

    \I__2780\ : ClkMux
    port map (
            O => \N__12128\,
            I => \N__11944\
        );

    \I__2779\ : ClkMux
    port map (
            O => \N__12127\,
            I => \N__11944\
        );

    \I__2778\ : ClkMux
    port map (
            O => \N__12126\,
            I => \N__11944\
        );

    \I__2777\ : ClkMux
    port map (
            O => \N__12125\,
            I => \N__11944\
        );

    \I__2776\ : ClkMux
    port map (
            O => \N__12124\,
            I => \N__11944\
        );

    \I__2775\ : ClkMux
    port map (
            O => \N__12123\,
            I => \N__11944\
        );

    \I__2774\ : ClkMux
    port map (
            O => \N__12122\,
            I => \N__11944\
        );

    \I__2773\ : ClkMux
    port map (
            O => \N__12121\,
            I => \N__11944\
        );

    \I__2772\ : ClkMux
    port map (
            O => \N__12120\,
            I => \N__11944\
        );

    \I__2771\ : ClkMux
    port map (
            O => \N__12119\,
            I => \N__11944\
        );

    \I__2770\ : ClkMux
    port map (
            O => \N__12118\,
            I => \N__11944\
        );

    \I__2769\ : ClkMux
    port map (
            O => \N__12117\,
            I => \N__11944\
        );

    \I__2768\ : ClkMux
    port map (
            O => \N__12116\,
            I => \N__11944\
        );

    \I__2767\ : ClkMux
    port map (
            O => \N__12115\,
            I => \N__11944\
        );

    \I__2766\ : ClkMux
    port map (
            O => \N__12114\,
            I => \N__11944\
        );

    \I__2765\ : ClkMux
    port map (
            O => \N__12113\,
            I => \N__11944\
        );

    \I__2764\ : ClkMux
    port map (
            O => \N__12112\,
            I => \N__11944\
        );

    \I__2763\ : ClkMux
    port map (
            O => \N__12111\,
            I => \N__11944\
        );

    \I__2762\ : ClkMux
    port map (
            O => \N__12110\,
            I => \N__11944\
        );

    \I__2761\ : ClkMux
    port map (
            O => \N__12109\,
            I => \N__11944\
        );

    \I__2760\ : ClkMux
    port map (
            O => \N__12108\,
            I => \N__11944\
        );

    \I__2759\ : ClkMux
    port map (
            O => \N__12107\,
            I => \N__11944\
        );

    \I__2758\ : ClkMux
    port map (
            O => \N__12106\,
            I => \N__11944\
        );

    \I__2757\ : ClkMux
    port map (
            O => \N__12105\,
            I => \N__11944\
        );

    \I__2756\ : ClkMux
    port map (
            O => \N__12104\,
            I => \N__11944\
        );

    \I__2755\ : ClkMux
    port map (
            O => \N__12103\,
            I => \N__11944\
        );

    \I__2754\ : ClkMux
    port map (
            O => \N__12102\,
            I => \N__11944\
        );

    \I__2753\ : ClkMux
    port map (
            O => \N__12101\,
            I => \N__11944\
        );

    \I__2752\ : ClkMux
    port map (
            O => \N__12100\,
            I => \N__11944\
        );

    \I__2751\ : ClkMux
    port map (
            O => \N__12099\,
            I => \N__11944\
        );

    \I__2750\ : ClkMux
    port map (
            O => \N__12098\,
            I => \N__11944\
        );

    \I__2749\ : ClkMux
    port map (
            O => \N__12097\,
            I => \N__11944\
        );

    \I__2748\ : ClkMux
    port map (
            O => \N__12096\,
            I => \N__11944\
        );

    \I__2747\ : ClkMux
    port map (
            O => \N__12095\,
            I => \N__11944\
        );

    \I__2746\ : ClkMux
    port map (
            O => \N__12094\,
            I => \N__11944\
        );

    \I__2745\ : ClkMux
    port map (
            O => \N__12093\,
            I => \N__11944\
        );

    \I__2744\ : ClkMux
    port map (
            O => \N__12092\,
            I => \N__11944\
        );

    \I__2743\ : ClkMux
    port map (
            O => \N__12091\,
            I => \N__11944\
        );

    \I__2742\ : ClkMux
    port map (
            O => \N__12090\,
            I => \N__11944\
        );

    \I__2741\ : ClkMux
    port map (
            O => \N__12089\,
            I => \N__11944\
        );

    \I__2740\ : ClkMux
    port map (
            O => \N__12088\,
            I => \N__11944\
        );

    \I__2739\ : ClkMux
    port map (
            O => \N__12087\,
            I => \N__11944\
        );

    \I__2738\ : ClkMux
    port map (
            O => \N__12086\,
            I => \N__11944\
        );

    \I__2737\ : ClkMux
    port map (
            O => \N__12085\,
            I => \N__11944\
        );

    \I__2736\ : ClkMux
    port map (
            O => \N__12084\,
            I => \N__11944\
        );

    \I__2735\ : ClkMux
    port map (
            O => \N__12083\,
            I => \N__11944\
        );

    \I__2734\ : ClkMux
    port map (
            O => \N__12082\,
            I => \N__11944\
        );

    \I__2733\ : ClkMux
    port map (
            O => \N__12081\,
            I => \N__11944\
        );

    \I__2732\ : ClkMux
    port map (
            O => \N__12080\,
            I => \N__11944\
        );

    \I__2731\ : ClkMux
    port map (
            O => \N__12079\,
            I => \N__11944\
        );

    \I__2730\ : ClkMux
    port map (
            O => \N__12078\,
            I => \N__11944\
        );

    \I__2729\ : ClkMux
    port map (
            O => \N__12077\,
            I => \N__11944\
        );

    \I__2728\ : ClkMux
    port map (
            O => \N__12076\,
            I => \N__11944\
        );

    \I__2727\ : ClkMux
    port map (
            O => \N__12075\,
            I => \N__11944\
        );

    \I__2726\ : GlobalMux
    port map (
            O => \N__11944\,
            I => clk_48mhz
        );

    \I__2725\ : CascadeMux
    port map (
            O => \N__11941\,
            I => \N__11932\
        );

    \I__2724\ : CascadeMux
    port map (
            O => \N__11940\,
            I => \N__11926\
        );

    \I__2723\ : InMux
    port map (
            O => \N__11939\,
            I => \N__11915\
        );

    \I__2722\ : InMux
    port map (
            O => \N__11938\,
            I => \N__11908\
        );

    \I__2721\ : InMux
    port map (
            O => \N__11937\,
            I => \N__11908\
        );

    \I__2720\ : InMux
    port map (
            O => \N__11936\,
            I => \N__11908\
        );

    \I__2719\ : InMux
    port map (
            O => \N__11935\,
            I => \N__11905\
        );

    \I__2718\ : InMux
    port map (
            O => \N__11932\,
            I => \N__11898\
        );

    \I__2717\ : InMux
    port map (
            O => \N__11931\,
            I => \N__11898\
        );

    \I__2716\ : InMux
    port map (
            O => \N__11930\,
            I => \N__11898\
        );

    \I__2715\ : InMux
    port map (
            O => \N__11929\,
            I => \N__11893\
        );

    \I__2714\ : InMux
    port map (
            O => \N__11926\,
            I => \N__11893\
        );

    \I__2713\ : InMux
    port map (
            O => \N__11925\,
            I => \N__11890\
        );

    \I__2712\ : InMux
    port map (
            O => \N__11924\,
            I => \N__11887\
        );

    \I__2711\ : InMux
    port map (
            O => \N__11923\,
            I => \N__11884\
        );

    \I__2710\ : InMux
    port map (
            O => \N__11922\,
            I => \N__11881\
        );

    \I__2709\ : InMux
    port map (
            O => \N__11921\,
            I => \N__11878\
        );

    \I__2708\ : InMux
    port map (
            O => \N__11920\,
            I => \N__11875\
        );

    \I__2707\ : InMux
    port map (
            O => \N__11919\,
            I => \N__11872\
        );

    \I__2706\ : InMux
    port map (
            O => \N__11918\,
            I => \N__11869\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__11915\,
            I => \N__11863\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__11908\,
            I => \N__11859\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__11905\,
            I => \N__11856\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__11898\,
            I => \N__11853\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__11893\,
            I => \N__11850\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__11890\,
            I => \N__11840\
        );

    \I__2699\ : LocalMux
    port map (
            O => \N__11887\,
            I => \N__11837\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__11884\,
            I => \N__11833\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__11881\,
            I => \N__11829\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__11878\,
            I => \N__11826\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__11875\,
            I => \N__11823\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__11872\,
            I => \N__11820\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__11869\,
            I => \N__11817\
        );

    \I__2692\ : CEMux
    port map (
            O => \N__11868\,
            I => \N__11764\
        );

    \I__2691\ : CEMux
    port map (
            O => \N__11867\,
            I => \N__11764\
        );

    \I__2690\ : CEMux
    port map (
            O => \N__11866\,
            I => \N__11764\
        );

    \I__2689\ : Glb2LocalMux
    port map (
            O => \N__11863\,
            I => \N__11764\
        );

    \I__2688\ : CEMux
    port map (
            O => \N__11862\,
            I => \N__11764\
        );

    \I__2687\ : Glb2LocalMux
    port map (
            O => \N__11859\,
            I => \N__11764\
        );

    \I__2686\ : Glb2LocalMux
    port map (
            O => \N__11856\,
            I => \N__11764\
        );

    \I__2685\ : Glb2LocalMux
    port map (
            O => \N__11853\,
            I => \N__11764\
        );

    \I__2684\ : Glb2LocalMux
    port map (
            O => \N__11850\,
            I => \N__11764\
        );

    \I__2683\ : CEMux
    port map (
            O => \N__11849\,
            I => \N__11764\
        );

    \I__2682\ : CEMux
    port map (
            O => \N__11848\,
            I => \N__11764\
        );

    \I__2681\ : CEMux
    port map (
            O => \N__11847\,
            I => \N__11764\
        );

    \I__2680\ : CEMux
    port map (
            O => \N__11846\,
            I => \N__11764\
        );

    \I__2679\ : CEMux
    port map (
            O => \N__11845\,
            I => \N__11764\
        );

    \I__2678\ : CEMux
    port map (
            O => \N__11844\,
            I => \N__11764\
        );

    \I__2677\ : CEMux
    port map (
            O => \N__11843\,
            I => \N__11764\
        );

    \I__2676\ : Glb2LocalMux
    port map (
            O => \N__11840\,
            I => \N__11764\
        );

    \I__2675\ : Glb2LocalMux
    port map (
            O => \N__11837\,
            I => \N__11764\
        );

    \I__2674\ : CEMux
    port map (
            O => \N__11836\,
            I => \N__11764\
        );

    \I__2673\ : Glb2LocalMux
    port map (
            O => \N__11833\,
            I => \N__11764\
        );

    \I__2672\ : CEMux
    port map (
            O => \N__11832\,
            I => \N__11764\
        );

    \I__2671\ : Glb2LocalMux
    port map (
            O => \N__11829\,
            I => \N__11764\
        );

    \I__2670\ : Glb2LocalMux
    port map (
            O => \N__11826\,
            I => \N__11764\
        );

    \I__2669\ : Glb2LocalMux
    port map (
            O => \N__11823\,
            I => \N__11764\
        );

    \I__2668\ : Glb2LocalMux
    port map (
            O => \N__11820\,
            I => \N__11764\
        );

    \I__2667\ : Glb2LocalMux
    port map (
            O => \N__11817\,
            I => \N__11764\
        );

    \I__2666\ : GlobalMux
    port map (
            O => \N__11764\,
            I => \N__11761\
        );

    \I__2665\ : gio2CtrlBuf
    port map (
            O => \N__11761\,
            I => \wPllLocked_g\
        );

    \I__2664\ : InMux
    port map (
            O => \N__11758\,
            I => \N__11754\
        );

    \I__2663\ : InMux
    port map (
            O => \N__11757\,
            I => \N__11751\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__11754\,
            I => \N__11748\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__11751\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_4\
        );

    \I__2660\ : Odrv4
    port map (
            O => \N__11748\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_4\
        );

    \I__2659\ : InMux
    port map (
            O => \N__11743\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_3\
        );

    \I__2658\ : InMux
    port map (
            O => \N__11740\,
            I => \N__11736\
        );

    \I__2657\ : InMux
    port map (
            O => \N__11739\,
            I => \N__11733\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__11736\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_5\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__11733\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_5\
        );

    \I__2654\ : InMux
    port map (
            O => \N__11728\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_4\
        );

    \I__2653\ : InMux
    port map (
            O => \N__11725\,
            I => \N__11721\
        );

    \I__2652\ : InMux
    port map (
            O => \N__11724\,
            I => \N__11718\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__11721\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_6\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__11718\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_6\
        );

    \I__2649\ : InMux
    port map (
            O => \N__11713\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_5\
        );

    \I__2648\ : InMux
    port map (
            O => \N__11710\,
            I => \N__11706\
        );

    \I__2647\ : InMux
    port map (
            O => \N__11709\,
            I => \N__11703\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__11706\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_7\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__11703\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_7\
        );

    \I__2644\ : InMux
    port map (
            O => \N__11698\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_6\
        );

    \I__2643\ : InMux
    port map (
            O => \N__11695\,
            I => \N__11691\
        );

    \I__2642\ : InMux
    port map (
            O => \N__11694\,
            I => \N__11688\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__11691\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_8\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__11688\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_8\
        );

    \I__2639\ : InMux
    port map (
            O => \N__11683\,
            I => \bfn_18_20_0_\
        );

    \I__2638\ : InMux
    port map (
            O => \N__11680\,
            I => \N__11676\
        );

    \I__2637\ : InMux
    port map (
            O => \N__11679\,
            I => \N__11673\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__11676\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_9\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__11673\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_9\
        );

    \I__2634\ : InMux
    port map (
            O => \N__11668\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_8\
        );

    \I__2633\ : InMux
    port map (
            O => \N__11665\,
            I => \N__11661\
        );

    \I__2632\ : InMux
    port map (
            O => \N__11664\,
            I => \N__11658\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__11661\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_10\
        );

    \I__2630\ : LocalMux
    port map (
            O => \N__11658\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_10\
        );

    \I__2629\ : InMux
    port map (
            O => \N__11653\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_9\
        );

    \I__2628\ : CascadeMux
    port map (
            O => \N__11650\,
            I => \N__11646\
        );

    \I__2627\ : InMux
    port map (
            O => \N__11649\,
            I => \N__11643\
        );

    \I__2626\ : InMux
    port map (
            O => \N__11646\,
            I => \N__11640\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__11643\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_11\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__11640\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_11\
        );

    \I__2623\ : InMux
    port map (
            O => \N__11635\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_10\
        );

    \I__2622\ : SRMux
    port map (
            O => \N__11632\,
            I => \N__11629\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__11629\,
            I => \N__11626\
        );

    \I__2620\ : Odrv12
    port map (
            O => \N__11626\,
            I => \DUT.uart_inst0.tx_bits_remaining_0_sqmuxa\
        );

    \I__2619\ : CascadeMux
    port map (
            O => \N__11623\,
            I => \N__11614\
        );

    \I__2618\ : InMux
    port map (
            O => \N__11622\,
            I => \N__11611\
        );

    \I__2617\ : InMux
    port map (
            O => \N__11621\,
            I => \N__11603\
        );

    \I__2616\ : InMux
    port map (
            O => \N__11620\,
            I => \N__11603\
        );

    \I__2615\ : InMux
    port map (
            O => \N__11619\,
            I => \N__11599\
        );

    \I__2614\ : InMux
    port map (
            O => \N__11618\,
            I => \N__11596\
        );

    \I__2613\ : InMux
    port map (
            O => \N__11617\,
            I => \N__11593\
        );

    \I__2612\ : InMux
    port map (
            O => \N__11614\,
            I => \N__11590\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__11611\,
            I => \N__11587\
        );

    \I__2610\ : InMux
    port map (
            O => \N__11610\,
            I => \N__11579\
        );

    \I__2609\ : InMux
    port map (
            O => \N__11609\,
            I => \N__11579\
        );

    \I__2608\ : InMux
    port map (
            O => \N__11608\,
            I => \N__11579\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__11603\,
            I => \N__11576\
        );

    \I__2606\ : InMux
    port map (
            O => \N__11602\,
            I => \N__11573\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__11599\,
            I => \N__11566\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__11596\,
            I => \N__11566\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__11593\,
            I => \N__11566\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__11590\,
            I => \N__11561\
        );

    \I__2601\ : Span4Mux_h
    port map (
            O => \N__11587\,
            I => \N__11561\
        );

    \I__2600\ : InMux
    port map (
            O => \N__11586\,
            I => \N__11558\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__11579\,
            I => \N__11553\
        );

    \I__2598\ : Span4Mux_h
    port map (
            O => \N__11576\,
            I => \N__11553\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__11573\,
            I => \DUT.rTransmitZ0\
        );

    \I__2596\ : Odrv12
    port map (
            O => \N__11566\,
            I => \DUT.rTransmitZ0\
        );

    \I__2595\ : Odrv4
    port map (
            O => \N__11561\,
            I => \DUT.rTransmitZ0\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__11558\,
            I => \DUT.rTransmitZ0\
        );

    \I__2593\ : Odrv4
    port map (
            O => \N__11553\,
            I => \DUT.rTransmitZ0\
        );

    \I__2592\ : InMux
    port map (
            O => \N__11542\,
            I => \N__11539\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__11539\,
            I => \DUT.uart_inst0.tx_clk_divider_0_sqmuxa\
        );

    \I__2590\ : IoInMux
    port map (
            O => \N__11536\,
            I => \N__11532\
        );

    \I__2589\ : CascadeMux
    port map (
            O => \N__11535\,
            I => \N__11528\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__11532\,
            I => \N__11521\
        );

    \I__2587\ : InMux
    port map (
            O => \N__11531\,
            I => \N__11517\
        );

    \I__2586\ : InMux
    port map (
            O => \N__11528\,
            I => \N__11512\
        );

    \I__2585\ : InMux
    port map (
            O => \N__11527\,
            I => \N__11512\
        );

    \I__2584\ : InMux
    port map (
            O => \N__11526\,
            I => \N__11507\
        );

    \I__2583\ : InMux
    port map (
            O => \N__11525\,
            I => \N__11507\
        );

    \I__2582\ : CascadeMux
    port map (
            O => \N__11524\,
            I => \N__11503\
        );

    \I__2581\ : Span4Mux_s1_v
    port map (
            O => \N__11521\,
            I => \N__11498\
        );

    \I__2580\ : CascadeMux
    port map (
            O => \N__11520\,
            I => \N__11495\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__11517\,
            I => \N__11489\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__11512\,
            I => \N__11489\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__11507\,
            I => \N__11486\
        );

    \I__2576\ : InMux
    port map (
            O => \N__11506\,
            I => \N__11483\
        );

    \I__2575\ : InMux
    port map (
            O => \N__11503\,
            I => \N__11478\
        );

    \I__2574\ : InMux
    port map (
            O => \N__11502\,
            I => \N__11478\
        );

    \I__2573\ : InMux
    port map (
            O => \N__11501\,
            I => \N__11475\
        );

    \I__2572\ : Sp12to4
    port map (
            O => \N__11498\,
            I => \N__11472\
        );

    \I__2571\ : InMux
    port map (
            O => \N__11495\,
            I => \N__11469\
        );

    \I__2570\ : InMux
    port map (
            O => \N__11494\,
            I => \N__11466\
        );

    \I__2569\ : Span4Mux_v
    port map (
            O => \N__11489\,
            I => \N__11463\
        );

    \I__2568\ : Span4Mux_v
    port map (
            O => \N__11486\,
            I => \N__11460\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__11483\,
            I => \N__11457\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__11478\,
            I => \N__11454\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__11475\,
            I => \N__11451\
        );

    \I__2564\ : Span12Mux_h
    port map (
            O => \N__11472\,
            I => \N__11448\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__11469\,
            I => \N__11445\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__11466\,
            I => \N__11442\
        );

    \I__2561\ : Span4Mux_h
    port map (
            O => \N__11463\,
            I => \N__11435\
        );

    \I__2560\ : Span4Mux_h
    port map (
            O => \N__11460\,
            I => \N__11435\
        );

    \I__2559\ : Span4Mux_v
    port map (
            O => \N__11457\,
            I => \N__11435\
        );

    \I__2558\ : Span4Mux_v
    port map (
            O => \N__11454\,
            I => \N__11430\
        );

    \I__2557\ : Span4Mux_v
    port map (
            O => \N__11451\,
            I => \N__11430\
        );

    \I__2556\ : Span12Mux_v
    port map (
            O => \N__11448\,
            I => \N__11427\
        );

    \I__2555\ : Span12Mux_v
    port map (
            O => \N__11445\,
            I => \N__11424\
        );

    \I__2554\ : Span12Mux_h
    port map (
            O => \N__11442\,
            I => \N__11417\
        );

    \I__2553\ : Sp12to4
    port map (
            O => \N__11435\,
            I => \N__11417\
        );

    \I__2552\ : Sp12to4
    port map (
            O => \N__11430\,
            I => \N__11417\
        );

    \I__2551\ : Span12Mux_v
    port map (
            O => \N__11427\,
            I => \N__11412\
        );

    \I__2550\ : Span12Mux_h
    port map (
            O => \N__11424\,
            I => \N__11412\
        );

    \I__2549\ : Span12Mux_h
    port map (
            O => \N__11417\,
            I => \N__11409\
        );

    \I__2548\ : Odrv12
    port map (
            O => \N__11412\,
            I => \wPllLocked\
        );

    \I__2547\ : Odrv12
    port map (
            O => \N__11409\,
            I => \wPllLocked\
        );

    \I__2546\ : CascadeMux
    port map (
            O => \N__11404\,
            I => \DUT.uart_inst0.tx_clk_divider_0_sqmuxa_cascade_\
        );

    \I__2545\ : InMux
    port map (
            O => \N__11401\,
            I => \N__11389\
        );

    \I__2544\ : InMux
    port map (
            O => \N__11400\,
            I => \N__11383\
        );

    \I__2543\ : InMux
    port map (
            O => \N__11399\,
            I => \N__11383\
        );

    \I__2542\ : InMux
    port map (
            O => \N__11398\,
            I => \N__11380\
        );

    \I__2541\ : InMux
    port map (
            O => \N__11397\,
            I => \N__11377\
        );

    \I__2540\ : InMux
    port map (
            O => \N__11396\,
            I => \N__11372\
        );

    \I__2539\ : InMux
    port map (
            O => \N__11395\,
            I => \N__11363\
        );

    \I__2538\ : InMux
    port map (
            O => \N__11394\,
            I => \N__11363\
        );

    \I__2537\ : InMux
    port map (
            O => \N__11393\,
            I => \N__11363\
        );

    \I__2536\ : InMux
    port map (
            O => \N__11392\,
            I => \N__11363\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__11389\,
            I => \N__11360\
        );

    \I__2534\ : InMux
    port map (
            O => \N__11388\,
            I => \N__11357\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__11383\,
            I => \N__11352\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__11380\,
            I => \N__11352\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__11377\,
            I => \N__11349\
        );

    \I__2530\ : InMux
    port map (
            O => \N__11376\,
            I => \N__11344\
        );

    \I__2529\ : InMux
    port map (
            O => \N__11375\,
            I => \N__11344\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__11372\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__11363\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0\
        );

    \I__2526\ : Odrv4
    port map (
            O => \N__11360\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__11357\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0\
        );

    \I__2524\ : Odrv4
    port map (
            O => \N__11352\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0\
        );

    \I__2523\ : Odrv4
    port map (
            O => \N__11349\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__11344\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0\
        );

    \I__2521\ : InMux
    port map (
            O => \N__11329\,
            I => \N__11323\
        );

    \I__2520\ : InMux
    port map (
            O => \N__11328\,
            I => \N__11323\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__11323\,
            I => \N__11319\
        );

    \I__2518\ : InMux
    port map (
            O => \N__11322\,
            I => \N__11316\
        );

    \I__2517\ : Odrv4
    port map (
            O => \N__11319\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__11316\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0\
        );

    \I__2515\ : InMux
    port map (
            O => \N__11311\,
            I => \N__11308\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__11308\,
            I => \N__11304\
        );

    \I__2513\ : InMux
    port map (
            O => \N__11307\,
            I => \N__11301\
        );

    \I__2512\ : Odrv4
    port map (
            O => \N__11304\,
            I => \fifo_inst.ftdi_output_inst.rRxF_nZ0Z_1\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__11301\,
            I => \fifo_inst.ftdi_output_inst.rRxF_nZ0Z_1\
        );

    \I__2510\ : InMux
    port map (
            O => \N__11296\,
            I => \N__11293\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__11293\,
            I => \N__11289\
        );

    \I__2508\ : InMux
    port map (
            O => \N__11292\,
            I => \N__11286\
        );

    \I__2507\ : Odrv12
    port map (
            O => \N__11289\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__11286\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1\
        );

    \I__2505\ : InMux
    port map (
            O => \N__11281\,
            I => \N__11278\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__11278\,
            I => \N__11273\
        );

    \I__2503\ : InMux
    port map (
            O => \N__11277\,
            I => \N__11270\
        );

    \I__2502\ : InMux
    port map (
            O => \N__11276\,
            I => \N__11267\
        );

    \I__2501\ : Span4Mux_h
    port map (
            O => \N__11273\,
            I => \N__11262\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__11270\,
            I => \N__11262\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__11267\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_0\
        );

    \I__2498\ : Odrv4
    port map (
            O => \N__11262\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_0\
        );

    \I__2497\ : InMux
    port map (
            O => \N__11257\,
            I => \N__11254\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__11254\,
            I => \N__11250\
        );

    \I__2495\ : InMux
    port map (
            O => \N__11253\,
            I => \N__11247\
        );

    \I__2494\ : Span4Mux_v
    port map (
            O => \N__11250\,
            I => \N__11244\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__11247\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_1\
        );

    \I__2492\ : Odrv4
    port map (
            O => \N__11244\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_1\
        );

    \I__2491\ : InMux
    port map (
            O => \N__11239\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_0\
        );

    \I__2490\ : CascadeMux
    port map (
            O => \N__11236\,
            I => \N__11232\
        );

    \I__2489\ : InMux
    port map (
            O => \N__11235\,
            I => \N__11229\
        );

    \I__2488\ : InMux
    port map (
            O => \N__11232\,
            I => \N__11226\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__11229\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_2\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__11226\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_2\
        );

    \I__2485\ : InMux
    port map (
            O => \N__11221\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_1\
        );

    \I__2484\ : InMux
    port map (
            O => \N__11218\,
            I => \N__11214\
        );

    \I__2483\ : InMux
    port map (
            O => \N__11217\,
            I => \N__11211\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__11214\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_3\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__11211\,
            I => \DUT.uart_inst0.tx_clk_dividerZ0Z_3\
        );

    \I__2480\ : InMux
    port map (
            O => \N__11206\,
            I => \DUT.uart_inst0.tx_clk_divider_cry_2\
        );

    \I__2479\ : CascadeMux
    port map (
            O => \N__11203\,
            I => \N__11197\
        );

    \I__2478\ : InMux
    port map (
            O => \N__11202\,
            I => \N__11191\
        );

    \I__2477\ : InMux
    port map (
            O => \N__11201\,
            I => \N__11182\
        );

    \I__2476\ : InMux
    port map (
            O => \N__11200\,
            I => \N__11182\
        );

    \I__2475\ : InMux
    port map (
            O => \N__11197\,
            I => \N__11182\
        );

    \I__2474\ : InMux
    port map (
            O => \N__11196\,
            I => \N__11182\
        );

    \I__2473\ : InMux
    port map (
            O => \N__11195\,
            I => \N__11169\
        );

    \I__2472\ : InMux
    port map (
            O => \N__11194\,
            I => \N__11169\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__11191\,
            I => \N__11164\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__11182\,
            I => \N__11164\
        );

    \I__2469\ : CascadeMux
    port map (
            O => \N__11181\,
            I => \N__11157\
        );

    \I__2468\ : CascadeMux
    port map (
            O => \N__11180\,
            I => \N__11153\
        );

    \I__2467\ : CascadeMux
    port map (
            O => \N__11179\,
            I => \N__11150\
        );

    \I__2466\ : CascadeMux
    port map (
            O => \N__11178\,
            I => \N__11147\
        );

    \I__2465\ : InMux
    port map (
            O => \N__11177\,
            I => \N__11138\
        );

    \I__2464\ : InMux
    port map (
            O => \N__11176\,
            I => \N__11138\
        );

    \I__2463\ : InMux
    port map (
            O => \N__11175\,
            I => \N__11138\
        );

    \I__2462\ : InMux
    port map (
            O => \N__11174\,
            I => \N__11135\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__11169\,
            I => \N__11132\
        );

    \I__2460\ : Span4Mux_h
    port map (
            O => \N__11164\,
            I => \N__11129\
        );

    \I__2459\ : InMux
    port map (
            O => \N__11163\,
            I => \N__11114\
        );

    \I__2458\ : InMux
    port map (
            O => \N__11162\,
            I => \N__11114\
        );

    \I__2457\ : InMux
    port map (
            O => \N__11161\,
            I => \N__11114\
        );

    \I__2456\ : InMux
    port map (
            O => \N__11160\,
            I => \N__11114\
        );

    \I__2455\ : InMux
    port map (
            O => \N__11157\,
            I => \N__11114\
        );

    \I__2454\ : InMux
    port map (
            O => \N__11156\,
            I => \N__11114\
        );

    \I__2453\ : InMux
    port map (
            O => \N__11153\,
            I => \N__11114\
        );

    \I__2452\ : InMux
    port map (
            O => \N__11150\,
            I => \N__11105\
        );

    \I__2451\ : InMux
    port map (
            O => \N__11147\,
            I => \N__11105\
        );

    \I__2450\ : InMux
    port map (
            O => \N__11146\,
            I => \N__11105\
        );

    \I__2449\ : InMux
    port map (
            O => \N__11145\,
            I => \N__11105\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__11138\,
            I => \N__11102\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__11135\,
            I => \N__11097\
        );

    \I__2446\ : Span4Mux_h
    port map (
            O => \N__11132\,
            I => \N__11097\
        );

    \I__2445\ : Odrv4
    port map (
            O => \N__11129\,
            I => \DUT.uart_inst0.N_72\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__11114\,
            I => \DUT.uart_inst0.N_72\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__11105\,
            I => \DUT.uart_inst0.N_72\
        );

    \I__2442\ : Odrv12
    port map (
            O => \N__11102\,
            I => \DUT.uart_inst0.N_72\
        );

    \I__2441\ : Odrv4
    port map (
            O => \N__11097\,
            I => \DUT.uart_inst0.N_72\
        );

    \I__2440\ : InMux
    port map (
            O => \N__11086\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_16\
        );

    \I__2439\ : CascadeMux
    port map (
            O => \N__11083\,
            I => \N__11079\
        );

    \I__2438\ : InMux
    port map (
            O => \N__11082\,
            I => \N__11076\
        );

    \I__2437\ : InMux
    port map (
            O => \N__11079\,
            I => \N__11073\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__11076\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_17\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__11073\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_17\
        );

    \I__2434\ : CascadeMux
    port map (
            O => \N__11068\,
            I => \N__11065\
        );

    \I__2433\ : InMux
    port map (
            O => \N__11065\,
            I => \N__11062\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__11062\,
            I => \N__11058\
        );

    \I__2431\ : CascadeMux
    port map (
            O => \N__11061\,
            I => \N__11055\
        );

    \I__2430\ : Span4Mux_v
    port map (
            O => \N__11058\,
            I => \N__11052\
        );

    \I__2429\ : InMux
    port map (
            O => \N__11055\,
            I => \N__11049\
        );

    \I__2428\ : Odrv4
    port map (
            O => \N__11052\,
            I => \fifo_inst.wRamRdAddr_2\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__11049\,
            I => \fifo_inst.wRamRdAddr_2\
        );

    \I__2426\ : InMux
    port map (
            O => \N__11044\,
            I => \N__11040\
        );

    \I__2425\ : CascadeMux
    port map (
            O => \N__11043\,
            I => \N__11037\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__11040\,
            I => \N__11031\
        );

    \I__2423\ : InMux
    port map (
            O => \N__11037\,
            I => \N__11026\
        );

    \I__2422\ : InMux
    port map (
            O => \N__11036\,
            I => \N__11026\
        );

    \I__2421\ : InMux
    port map (
            O => \N__11035\,
            I => \N__11021\
        );

    \I__2420\ : InMux
    port map (
            O => \N__11034\,
            I => \N__11021\
        );

    \I__2419\ : Odrv4
    port map (
            O => \N__11031\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__11026\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__11021\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4\
        );

    \I__2416\ : InMux
    port map (
            O => \N__11014\,
            I => \N__11006\
        );

    \I__2415\ : InMux
    port map (
            O => \N__11013\,
            I => \N__11006\
        );

    \I__2414\ : InMux
    port map (
            O => \N__11012\,
            I => \N__11000\
        );

    \I__2413\ : InMux
    port map (
            O => \N__11011\,
            I => \N__11000\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__11006\,
            I => \N__10997\
        );

    \I__2411\ : InMux
    port map (
            O => \N__11005\,
            I => \N__10994\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__11000\,
            I => \N__10991\
        );

    \I__2409\ : Span4Mux_h
    port map (
            O => \N__10997\,
            I => \N__10988\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__10994\,
            I => \fifo_inst.ftdi_output_inst.rWrDelayZ0\
        );

    \I__2407\ : Odrv4
    port map (
            O => \N__10991\,
            I => \fifo_inst.ftdi_output_inst.rWrDelayZ0\
        );

    \I__2406\ : Odrv4
    port map (
            O => \N__10988\,
            I => \fifo_inst.ftdi_output_inst.rWrDelayZ0\
        );

    \I__2405\ : InMux
    port map (
            O => \N__10981\,
            I => \N__10978\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__10978\,
            I => \fifo_inst.ftdi_output_inst.N_3_0\
        );

    \I__2403\ : CascadeMux
    port map (
            O => \N__10975\,
            I => \N__10972\
        );

    \I__2402\ : InMux
    port map (
            O => \N__10972\,
            I => \N__10969\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__10969\,
            I => \N__10966\
        );

    \I__2400\ : Span4Mux_v
    port map (
            O => \N__10966\,
            I => \N__10960\
        );

    \I__2399\ : InMux
    port map (
            O => \N__10965\,
            I => \N__10953\
        );

    \I__2398\ : InMux
    port map (
            O => \N__10964\,
            I => \N__10953\
        );

    \I__2397\ : InMux
    port map (
            O => \N__10963\,
            I => \N__10953\
        );

    \I__2396\ : Odrv4
    port map (
            O => \N__10960\,
            I => \fifo_inst.wRamRdAddr_0\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__10953\,
            I => \fifo_inst.wRamRdAddr_0\
        );

    \I__2394\ : CascadeMux
    port map (
            O => \N__10948\,
            I => \fifo_inst.ftdi_output_inst.N_3_0_cascade_\
        );

    \I__2393\ : CascadeMux
    port map (
            O => \N__10945\,
            I => \N__10942\
        );

    \I__2392\ : InMux
    port map (
            O => \N__10942\,
            I => \N__10939\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__10939\,
            I => \N__10936\
        );

    \I__2390\ : Span4Mux_v
    port map (
            O => \N__10936\,
            I => \N__10933\
        );

    \I__2389\ : Span4Mux_v
    port map (
            O => \N__10933\,
            I => \N__10928\
        );

    \I__2388\ : InMux
    port map (
            O => \N__10932\,
            I => \N__10923\
        );

    \I__2387\ : InMux
    port map (
            O => \N__10931\,
            I => \N__10923\
        );

    \I__2386\ : Odrv4
    port map (
            O => \N__10928\,
            I => \fifo_inst.wRamRdAddr_1\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__10923\,
            I => \fifo_inst.wRamRdAddr_1\
        );

    \I__2384\ : InMux
    port map (
            O => \N__10918\,
            I => \N__10915\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__10915\,
            I => \N__10912\
        );

    \I__2382\ : Span4Mux_h
    port map (
            O => \N__10912\,
            I => \N__10909\
        );

    \I__2381\ : Odrv4
    port map (
            O => \N__10909\,
            I => \DUT.uart_inst0.tx_state_ns_i_i_a2_0_0_0\
        );

    \I__2380\ : CascadeMux
    port map (
            O => \N__10906\,
            I => \N__10901\
        );

    \I__2379\ : InMux
    port map (
            O => \N__10905\,
            I => \N__10893\
        );

    \I__2378\ : InMux
    port map (
            O => \N__10904\,
            I => \N__10890\
        );

    \I__2377\ : InMux
    port map (
            O => \N__10901\,
            I => \N__10883\
        );

    \I__2376\ : InMux
    port map (
            O => \N__10900\,
            I => \N__10883\
        );

    \I__2375\ : InMux
    port map (
            O => \N__10899\,
            I => \N__10883\
        );

    \I__2374\ : InMux
    port map (
            O => \N__10898\,
            I => \N__10878\
        );

    \I__2373\ : InMux
    port map (
            O => \N__10897\,
            I => \N__10878\
        );

    \I__2372\ : InMux
    port map (
            O => \N__10896\,
            I => \N__10875\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__10893\,
            I => \N__10872\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__10890\,
            I => \N__10864\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__10883\,
            I => \N__10864\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__10878\,
            I => \N__10859\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__10875\,
            I => \N__10859\
        );

    \I__2366\ : Span4Mux_h
    port map (
            O => \N__10872\,
            I => \N__10856\
        );

    \I__2365\ : InMux
    port map (
            O => \N__10871\,
            I => \N__10849\
        );

    \I__2364\ : InMux
    port map (
            O => \N__10870\,
            I => \N__10849\
        );

    \I__2363\ : InMux
    port map (
            O => \N__10869\,
            I => \N__10849\
        );

    \I__2362\ : Span4Mux_v
    port map (
            O => \N__10864\,
            I => \N__10846\
        );

    \I__2361\ : Span4Mux_h
    port map (
            O => \N__10859\,
            I => \N__10843\
        );

    \I__2360\ : Span4Mux_v
    port map (
            O => \N__10856\,
            I => \N__10840\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__10849\,
            I => \DUT.uart_inst0.tx_state_0_sqmuxa_i_0\
        );

    \I__2358\ : Odrv4
    port map (
            O => \N__10846\,
            I => \DUT.uart_inst0.tx_state_0_sqmuxa_i_0\
        );

    \I__2357\ : Odrv4
    port map (
            O => \N__10843\,
            I => \DUT.uart_inst0.tx_state_0_sqmuxa_i_0\
        );

    \I__2356\ : Odrv4
    port map (
            O => \N__10840\,
            I => \DUT.uart_inst0.tx_state_0_sqmuxa_i_0\
        );

    \I__2355\ : InMux
    port map (
            O => \N__10831\,
            I => \N__10827\
        );

    \I__2354\ : IoInMux
    port map (
            O => \N__10830\,
            I => \N__10824\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__10827\,
            I => \N__10821\
        );

    \I__2352\ : LocalMux
    port map (
            O => \N__10824\,
            I => \N__10818\
        );

    \I__2351\ : Span4Mux_v
    port map (
            O => \N__10821\,
            I => \N__10815\
        );

    \I__2350\ : Span12Mux_s10_v
    port map (
            O => \N__10818\,
            I => \N__10812\
        );

    \I__2349\ : Span4Mux_h
    port map (
            O => \N__10815\,
            I => \N__10809\
        );

    \I__2348\ : Odrv12
    port map (
            O => \N__10812\,
            I => \wPllLocked_iso_i\
        );

    \I__2347\ : Odrv4
    port map (
            O => \N__10809\,
            I => \wPllLocked_iso_i\
        );

    \I__2346\ : CEMux
    port map (
            O => \N__10804\,
            I => \N__10801\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__10801\,
            I => \DUT.uart_inst0.N_345_0_0\
        );

    \I__2344\ : InMux
    port map (
            O => \N__10798\,
            I => \N__10793\
        );

    \I__2343\ : InMux
    port map (
            O => \N__10797\,
            I => \N__10790\
        );

    \I__2342\ : InMux
    port map (
            O => \N__10796\,
            I => \N__10787\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__10793\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_9\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__10790\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_9\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__10787\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_9\
        );

    \I__2338\ : InMux
    port map (
            O => \N__10780\,
            I => \N__10777\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__10777\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO\
        );

    \I__2336\ : InMux
    port map (
            O => \N__10774\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_8\
        );

    \I__2335\ : InMux
    port map (
            O => \N__10771\,
            I => \N__10766\
        );

    \I__2334\ : InMux
    port map (
            O => \N__10770\,
            I => \N__10761\
        );

    \I__2333\ : InMux
    port map (
            O => \N__10769\,
            I => \N__10761\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__10766\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_10\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__10761\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_10\
        );

    \I__2330\ : InMux
    port map (
            O => \N__10756\,
            I => \N__10753\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__10753\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO\
        );

    \I__2328\ : InMux
    port map (
            O => \N__10750\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_9\
        );

    \I__2327\ : InMux
    port map (
            O => \N__10747\,
            I => \N__10742\
        );

    \I__2326\ : InMux
    port map (
            O => \N__10746\,
            I => \N__10737\
        );

    \I__2325\ : InMux
    port map (
            O => \N__10745\,
            I => \N__10737\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__10742\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_11\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__10737\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_11\
        );

    \I__2322\ : InMux
    port map (
            O => \N__10732\,
            I => \N__10729\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__10729\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO\
        );

    \I__2320\ : InMux
    port map (
            O => \N__10726\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_10\
        );

    \I__2319\ : CascadeMux
    port map (
            O => \N__10723\,
            I => \N__10718\
        );

    \I__2318\ : InMux
    port map (
            O => \N__10722\,
            I => \N__10715\
        );

    \I__2317\ : InMux
    port map (
            O => \N__10721\,
            I => \N__10710\
        );

    \I__2316\ : InMux
    port map (
            O => \N__10718\,
            I => \N__10710\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__10715\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_12\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__10710\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_12\
        );

    \I__2313\ : InMux
    port map (
            O => \N__10705\,
            I => \N__10702\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__10702\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO\
        );

    \I__2311\ : InMux
    port map (
            O => \N__10699\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_11\
        );

    \I__2310\ : InMux
    port map (
            O => \N__10696\,
            I => \N__10691\
        );

    \I__2309\ : InMux
    port map (
            O => \N__10695\,
            I => \N__10686\
        );

    \I__2308\ : InMux
    port map (
            O => \N__10694\,
            I => \N__10686\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__10691\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_13\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__10686\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_13\
        );

    \I__2305\ : CascadeMux
    port map (
            O => \N__10681\,
            I => \N__10678\
        );

    \I__2304\ : InMux
    port map (
            O => \N__10678\,
            I => \N__10675\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__10675\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO\
        );

    \I__2302\ : InMux
    port map (
            O => \N__10672\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_12\
        );

    \I__2301\ : InMux
    port map (
            O => \N__10669\,
            I => \N__10664\
        );

    \I__2300\ : InMux
    port map (
            O => \N__10668\,
            I => \N__10661\
        );

    \I__2299\ : InMux
    port map (
            O => \N__10667\,
            I => \N__10658\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__10664\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_14\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__10661\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_14\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__10658\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_14\
        );

    \I__2295\ : InMux
    port map (
            O => \N__10651\,
            I => \N__10648\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__10648\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO\
        );

    \I__2293\ : InMux
    port map (
            O => \N__10645\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_13\
        );

    \I__2292\ : InMux
    port map (
            O => \N__10642\,
            I => \N__10637\
        );

    \I__2291\ : InMux
    port map (
            O => \N__10641\,
            I => \N__10632\
        );

    \I__2290\ : InMux
    port map (
            O => \N__10640\,
            I => \N__10632\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__10637\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_15\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__10632\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_15\
        );

    \I__2287\ : CascadeMux
    port map (
            O => \N__10627\,
            I => \N__10624\
        );

    \I__2286\ : InMux
    port map (
            O => \N__10624\,
            I => \N__10621\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__10621\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO\
        );

    \I__2284\ : InMux
    port map (
            O => \N__10618\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_14\
        );

    \I__2283\ : InMux
    port map (
            O => \N__10615\,
            I => \N__10610\
        );

    \I__2282\ : InMux
    port map (
            O => \N__10614\,
            I => \N__10607\
        );

    \I__2281\ : InMux
    port map (
            O => \N__10613\,
            I => \N__10604\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__10610\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_16\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__10607\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_16\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__10604\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_16\
        );

    \I__2277\ : InMux
    port map (
            O => \N__10597\,
            I => \N__10594\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__10594\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO\
        );

    \I__2275\ : InMux
    port map (
            O => \N__10591\,
            I => \bfn_18_15_0_\
        );

    \I__2274\ : InMux
    port map (
            O => \N__10588\,
            I => \N__10583\
        );

    \I__2273\ : InMux
    port map (
            O => \N__10587\,
            I => \N__10580\
        );

    \I__2272\ : InMux
    port map (
            O => \N__10586\,
            I => \N__10577\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__10583\,
            I => \DUT.uart_inst0.rx_clk_dividerZ1Z_1\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__10580\,
            I => \DUT.uart_inst0.rx_clk_dividerZ1Z_1\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__10577\,
            I => \DUT.uart_inst0.rx_clk_dividerZ1Z_1\
        );

    \I__2268\ : InMux
    port map (
            O => \N__10570\,
            I => \N__10567\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__10567\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO\
        );

    \I__2266\ : InMux
    port map (
            O => \N__10564\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_0\
        );

    \I__2265\ : InMux
    port map (
            O => \N__10561\,
            I => \N__10558\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__10558\,
            I => \N__10553\
        );

    \I__2263\ : InMux
    port map (
            O => \N__10557\,
            I => \N__10548\
        );

    \I__2262\ : InMux
    port map (
            O => \N__10556\,
            I => \N__10548\
        );

    \I__2261\ : Odrv4
    port map (
            O => \N__10553\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_2\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__10548\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_2\
        );

    \I__2259\ : InMux
    port map (
            O => \N__10543\,
            I => \N__10540\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__10540\,
            I => \N__10537\
        );

    \I__2257\ : Odrv4
    port map (
            O => \N__10537\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO\
        );

    \I__2256\ : InMux
    port map (
            O => \N__10534\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_1\
        );

    \I__2255\ : InMux
    port map (
            O => \N__10531\,
            I => \N__10527\
        );

    \I__2254\ : CascadeMux
    port map (
            O => \N__10530\,
            I => \N__10523\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__10527\,
            I => \N__10520\
        );

    \I__2252\ : InMux
    port map (
            O => \N__10526\,
            I => \N__10517\
        );

    \I__2251\ : InMux
    port map (
            O => \N__10523\,
            I => \N__10514\
        );

    \I__2250\ : Span4Mux_h
    port map (
            O => \N__10520\,
            I => \N__10511\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__10517\,
            I => \N__10508\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__10514\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_3\
        );

    \I__2247\ : Odrv4
    port map (
            O => \N__10511\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_3\
        );

    \I__2246\ : Odrv4
    port map (
            O => \N__10508\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_3\
        );

    \I__2245\ : InMux
    port map (
            O => \N__10501\,
            I => \N__10498\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__10498\,
            I => \N__10495\
        );

    \I__2243\ : Span4Mux_v
    port map (
            O => \N__10495\,
            I => \N__10492\
        );

    \I__2242\ : Odrv4
    port map (
            O => \N__10492\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_2_THRU_CO\
        );

    \I__2241\ : InMux
    port map (
            O => \N__10489\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_2\
        );

    \I__2240\ : CascadeMux
    port map (
            O => \N__10486\,
            I => \N__10481\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__10485\,
            I => \N__10478\
        );

    \I__2238\ : InMux
    port map (
            O => \N__10484\,
            I => \N__10475\
        );

    \I__2237\ : InMux
    port map (
            O => \N__10481\,
            I => \N__10472\
        );

    \I__2236\ : InMux
    port map (
            O => \N__10478\,
            I => \N__10469\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__10475\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_4\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__10472\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_4\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__10469\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_4\
        );

    \I__2232\ : InMux
    port map (
            O => \N__10462\,
            I => \N__10459\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__10459\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO\
        );

    \I__2230\ : InMux
    port map (
            O => \N__10456\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_3\
        );

    \I__2229\ : InMux
    port map (
            O => \N__10453\,
            I => \N__10448\
        );

    \I__2228\ : InMux
    port map (
            O => \N__10452\,
            I => \N__10445\
        );

    \I__2227\ : InMux
    port map (
            O => \N__10451\,
            I => \N__10442\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__10448\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_5\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__10445\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_5\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__10442\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_5\
        );

    \I__2223\ : InMux
    port map (
            O => \N__10435\,
            I => \N__10432\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__10432\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_4_THRU_CO\
        );

    \I__2221\ : InMux
    port map (
            O => \N__10429\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_4\
        );

    \I__2220\ : InMux
    port map (
            O => \N__10426\,
            I => \N__10421\
        );

    \I__2219\ : InMux
    port map (
            O => \N__10425\,
            I => \N__10418\
        );

    \I__2218\ : InMux
    port map (
            O => \N__10424\,
            I => \N__10415\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__10421\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_6\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__10418\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_6\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__10415\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_6\
        );

    \I__2214\ : InMux
    port map (
            O => \N__10408\,
            I => \N__10405\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__10405\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_5_THRU_CO\
        );

    \I__2212\ : InMux
    port map (
            O => \N__10402\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_5\
        );

    \I__2211\ : InMux
    port map (
            O => \N__10399\,
            I => \N__10394\
        );

    \I__2210\ : InMux
    port map (
            O => \N__10398\,
            I => \N__10391\
        );

    \I__2209\ : InMux
    port map (
            O => \N__10397\,
            I => \N__10388\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__10394\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_7\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__10391\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_7\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__10388\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_7\
        );

    \I__2205\ : InMux
    port map (
            O => \N__10381\,
            I => \N__10378\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__10378\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO\
        );

    \I__2203\ : InMux
    port map (
            O => \N__10375\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_6\
        );

    \I__2202\ : CascadeMux
    port map (
            O => \N__10372\,
            I => \N__10368\
        );

    \I__2201\ : InMux
    port map (
            O => \N__10371\,
            I => \N__10364\
        );

    \I__2200\ : InMux
    port map (
            O => \N__10368\,
            I => \N__10361\
        );

    \I__2199\ : InMux
    port map (
            O => \N__10367\,
            I => \N__10358\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__10364\,
            I => \N__10355\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__10361\,
            I => \N__10352\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__10358\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_8\
        );

    \I__2195\ : Odrv4
    port map (
            O => \N__10355\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_8\
        );

    \I__2194\ : Odrv4
    port map (
            O => \N__10352\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_8\
        );

    \I__2193\ : InMux
    port map (
            O => \N__10345\,
            I => \N__10342\
        );

    \I__2192\ : LocalMux
    port map (
            O => \N__10342\,
            I => \N__10339\
        );

    \I__2191\ : Odrv4
    port map (
            O => \N__10339\,
            I => \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO\
        );

    \I__2190\ : InMux
    port map (
            O => \N__10336\,
            I => \bfn_18_14_0_\
        );

    \I__2189\ : CascadeMux
    port map (
            O => \N__10333\,
            I => \N__10328\
        );

    \I__2188\ : InMux
    port map (
            O => \N__10332\,
            I => \N__10324\
        );

    \I__2187\ : CascadeMux
    port map (
            O => \N__10331\,
            I => \N__10321\
        );

    \I__2186\ : InMux
    port map (
            O => \N__10328\,
            I => \N__10318\
        );

    \I__2185\ : InMux
    port map (
            O => \N__10327\,
            I => \N__10315\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__10324\,
            I => \N__10312\
        );

    \I__2183\ : InMux
    port map (
            O => \N__10321\,
            I => \N__10309\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__10318\,
            I => \N__10306\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__10315\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_3\
        );

    \I__2180\ : Odrv4
    port map (
            O => \N__10312\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_3\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__10309\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_3\
        );

    \I__2178\ : Odrv4
    port map (
            O => \N__10306\,
            I => \DUT.uart_inst0.tx_bits_remainingZ0Z_3\
        );

    \I__2177\ : CascadeMux
    port map (
            O => \N__10297\,
            I => \DUT.uart_inst0.tx_state_ns_i_i_a2_0_0_0_cascade_\
        );

    \I__2176\ : InMux
    port map (
            O => \N__10294\,
            I => \N__10291\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__10291\,
            I => \DUT.uart_inst0.g0_i_a4_1_0\
        );

    \I__2174\ : InMux
    port map (
            O => \N__10288\,
            I => \N__10285\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__10285\,
            I => \N__10282\
        );

    \I__2172\ : Span4Mux_h
    port map (
            O => \N__10282\,
            I => \N__10279\
        );

    \I__2171\ : Odrv4
    port map (
            O => \N__10279\,
            I => \DUT.uart_inst0.d_N_5_mux\
        );

    \I__2170\ : InMux
    port map (
            O => \N__10276\,
            I => \N__10272\
        );

    \I__2169\ : InMux
    port map (
            O => \N__10275\,
            I => \N__10269\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__10272\,
            I => \N__10262\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__10269\,
            I => \N__10262\
        );

    \I__2166\ : InMux
    port map (
            O => \N__10268\,
            I => \N__10259\
        );

    \I__2165\ : InMux
    port map (
            O => \N__10267\,
            I => \N__10256\
        );

    \I__2164\ : Span12Mux_h
    port map (
            O => \N__10262\,
            I => \N__10249\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__10259\,
            I => \N__10249\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__10256\,
            I => \N__10249\
        );

    \I__2161\ : Odrv12
    port map (
            O => \N__10249\,
            I => \rTxByteZ0Z_3\
        );

    \I__2160\ : InMux
    port map (
            O => \N__10246\,
            I => \N__10243\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__10243\,
            I => \N__10240\
        );

    \I__2158\ : Odrv4
    port map (
            O => \N__10240\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_3\
        );

    \I__2157\ : CEMux
    port map (
            O => \N__10237\,
            I => \N__10234\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__10234\,
            I => \N__10230\
        );

    \I__2155\ : CEMux
    port map (
            O => \N__10233\,
            I => \N__10226\
        );

    \I__2154\ : Span4Mux_v
    port map (
            O => \N__10230\,
            I => \N__10223\
        );

    \I__2153\ : CEMux
    port map (
            O => \N__10229\,
            I => \N__10220\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__10226\,
            I => \N__10217\
        );

    \I__2151\ : Span4Mux_h
    port map (
            O => \N__10223\,
            I => \N__10212\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__10220\,
            I => \N__10212\
        );

    \I__2149\ : Span12Mux_h
    port map (
            O => \N__10217\,
            I => \N__10208\
        );

    \I__2148\ : Span4Mux_v
    port map (
            O => \N__10212\,
            I => \N__10205\
        );

    \I__2147\ : CEMux
    port map (
            O => \N__10211\,
            I => \N__10202\
        );

    \I__2146\ : Odrv12
    port map (
            O => \N__10208\,
            I => \DUT.fifo_tx_inst.N_39\
        );

    \I__2145\ : Odrv4
    port map (
            O => \N__10205\,
            I => \DUT.fifo_tx_inst.N_39\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__10202\,
            I => \DUT.fifo_tx_inst.N_39\
        );

    \I__2143\ : InMux
    port map (
            O => \N__10195\,
            I => \N__10192\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__10192\,
            I => \N__10189\
        );

    \I__2141\ : Span4Mux_v
    port map (
            O => \N__10189\,
            I => \N__10186\
        );

    \I__2140\ : Odrv4
    port map (
            O => \N__10186\,
            I => \fifo_inst.ftdi_output_inst.rTxE_nZ0Z_1\
        );

    \I__2139\ : InMux
    port map (
            O => \N__10183\,
            I => \N__10180\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__10180\,
            I => \N__10177\
        );

    \I__2137\ : Span4Mux_v
    port map (
            O => \N__10177\,
            I => \N__10174\
        );

    \I__2136\ : Odrv4
    port map (
            O => \N__10174\,
            I => \iTxE_n_c\
        );

    \I__2135\ : InMux
    port map (
            O => \N__10171\,
            I => \N__10168\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__10168\,
            I => \N__10164\
        );

    \I__2133\ : InMux
    port map (
            O => \N__10167\,
            I => \N__10161\
        );

    \I__2132\ : Span4Mux_v
    port map (
            O => \N__10164\,
            I => \N__10158\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__10161\,
            I => \fifo_inst.ftdi_output_inst.rTxE_nZ0Z_0\
        );

    \I__2130\ : Odrv4
    port map (
            O => \N__10158\,
            I => \fifo_inst.ftdi_output_inst.rTxE_nZ0Z_0\
        );

    \I__2129\ : InMux
    port map (
            O => \N__10153\,
            I => \N__10148\
        );

    \I__2128\ : InMux
    port map (
            O => \N__10152\,
            I => \N__10145\
        );

    \I__2127\ : InMux
    port map (
            O => \N__10151\,
            I => \N__10142\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__10148\,
            I => \N__10139\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__10145\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_1\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__10142\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_1\
        );

    \I__2123\ : Odrv4
    port map (
            O => \N__10139\,
            I => \DUT.uart_inst0.rx_clk_dividerZ0Z_1\
        );

    \I__2122\ : InMux
    port map (
            O => \N__10132\,
            I => \N__10129\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__10129\,
            I => \N__10126\
        );

    \I__2120\ : Span4Mux_h
    port map (
            O => \N__10126\,
            I => \N__10123\
        );

    \I__2119\ : Odrv4
    port map (
            O => \N__10123\,
            I => \DUT.rFifoDatarx_6\
        );

    \I__2118\ : CascadeMux
    port map (
            O => \N__10120\,
            I => \N__10117\
        );

    \I__2117\ : InMux
    port map (
            O => \N__10117\,
            I => \N__10113\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__10116\,
            I => \N__10110\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__10113\,
            I => \N__10107\
        );

    \I__2114\ : InMux
    port map (
            O => \N__10110\,
            I => \N__10104\
        );

    \I__2113\ : Span4Mux_h
    port map (
            O => \N__10107\,
            I => \N__10101\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__10104\,
            I => \DUT.uart_inst0.tx_dataZ0Z_7\
        );

    \I__2111\ : Odrv4
    port map (
            O => \N__10101\,
            I => \DUT.uart_inst0.tx_dataZ0Z_7\
        );

    \I__2110\ : CascadeMux
    port map (
            O => \N__10096\,
            I => \DUT.uart_inst0.tx_data_RNO_0Z0Z_6_cascade_\
        );

    \I__2109\ : InMux
    port map (
            O => \N__10093\,
            I => \N__10090\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__10090\,
            I => \N__10086\
        );

    \I__2107\ : InMux
    port map (
            O => \N__10089\,
            I => \N__10083\
        );

    \I__2106\ : Span4Mux_h
    port map (
            O => \N__10086\,
            I => \N__10080\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__10083\,
            I => \DUT.uart_inst0.tx_dataZ0Z_6\
        );

    \I__2104\ : Odrv4
    port map (
            O => \N__10080\,
            I => \DUT.uart_inst0.tx_dataZ0Z_6\
        );

    \I__2103\ : CascadeMux
    port map (
            O => \N__10075\,
            I => \N__10071\
        );

    \I__2102\ : CascadeMux
    port map (
            O => \N__10074\,
            I => \N__10068\
        );

    \I__2101\ : InMux
    port map (
            O => \N__10071\,
            I => \N__10065\
        );

    \I__2100\ : InMux
    port map (
            O => \N__10068\,
            I => \N__10062\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__10065\,
            I => \N__10057\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__10062\,
            I => \N__10057\
        );

    \I__2097\ : Odrv4
    port map (
            O => \N__10057\,
            I => \DUT.uart_inst0.tx_dataZ0Z_4\
        );

    \I__2096\ : InMux
    port map (
            O => \N__10054\,
            I => \N__10049\
        );

    \I__2095\ : InMux
    port map (
            O => \N__10053\,
            I => \N__10044\
        );

    \I__2094\ : InMux
    port map (
            O => \N__10052\,
            I => \N__10044\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__10049\,
            I => \N__10036\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__10044\,
            I => \N__10036\
        );

    \I__2091\ : InMux
    port map (
            O => \N__10043\,
            I => \N__10031\
        );

    \I__2090\ : InMux
    port map (
            O => \N__10042\,
            I => \N__10031\
        );

    \I__2089\ : InMux
    port map (
            O => \N__10041\,
            I => \N__10027\
        );

    \I__2088\ : Span4Mux_v
    port map (
            O => \N__10036\,
            I => \N__10023\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__10031\,
            I => \N__10020\
        );

    \I__2086\ : InMux
    port map (
            O => \N__10030\,
            I => \N__10017\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__10027\,
            I => \N__10014\
        );

    \I__2084\ : InMux
    port map (
            O => \N__10026\,
            I => \N__10011\
        );

    \I__2083\ : Odrv4
    port map (
            O => \N__10023\,
            I => \DUT.rFifoDataror_0\
        );

    \I__2082\ : Odrv4
    port map (
            O => \N__10020\,
            I => \DUT.rFifoDataror_0\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__10017\,
            I => \DUT.rFifoDataror_0\
        );

    \I__2080\ : Odrv4
    port map (
            O => \N__10014\,
            I => \DUT.rFifoDataror_0\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__10011\,
            I => \DUT.rFifoDataror_0\
        );

    \I__2078\ : CascadeMux
    port map (
            O => \N__10000\,
            I => \DUT.uart_inst0.tx_data_RNO_0Z0Z_3_cascade_\
        );

    \I__2077\ : CEMux
    port map (
            O => \N__9997\,
            I => \N__9994\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__9994\,
            I => \N__9979\
        );

    \I__2075\ : InMux
    port map (
            O => \N__9993\,
            I => \N__9976\
        );

    \I__2074\ : InMux
    port map (
            O => \N__9992\,
            I => \N__9969\
        );

    \I__2073\ : InMux
    port map (
            O => \N__9991\,
            I => \N__9969\
        );

    \I__2072\ : InMux
    port map (
            O => \N__9990\,
            I => \N__9969\
        );

    \I__2071\ : InMux
    port map (
            O => \N__9989\,
            I => \N__9961\
        );

    \I__2070\ : InMux
    port map (
            O => \N__9988\,
            I => \N__9956\
        );

    \I__2069\ : InMux
    port map (
            O => \N__9987\,
            I => \N__9956\
        );

    \I__2068\ : InMux
    port map (
            O => \N__9986\,
            I => \N__9953\
        );

    \I__2067\ : InMux
    port map (
            O => \N__9985\,
            I => \N__9944\
        );

    \I__2066\ : InMux
    port map (
            O => \N__9984\,
            I => \N__9944\
        );

    \I__2065\ : InMux
    port map (
            O => \N__9983\,
            I => \N__9944\
        );

    \I__2064\ : InMux
    port map (
            O => \N__9982\,
            I => \N__9944\
        );

    \I__2063\ : Span4Mux_v
    port map (
            O => \N__9979\,
            I => \N__9937\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__9976\,
            I => \N__9937\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__9969\,
            I => \N__9937\
        );

    \I__2060\ : InMux
    port map (
            O => \N__9968\,
            I => \N__9932\
        );

    \I__2059\ : InMux
    port map (
            O => \N__9967\,
            I => \N__9932\
        );

    \I__2058\ : InMux
    port map (
            O => \N__9966\,
            I => \N__9925\
        );

    \I__2057\ : InMux
    port map (
            O => \N__9965\,
            I => \N__9925\
        );

    \I__2056\ : InMux
    port map (
            O => \N__9964\,
            I => \N__9925\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__9961\,
            I => \DUT.uart_inst0.N_152_0\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__9956\,
            I => \DUT.uart_inst0.N_152_0\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__9953\,
            I => \DUT.uart_inst0.N_152_0\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__9944\,
            I => \DUT.uart_inst0.N_152_0\
        );

    \I__2051\ : Odrv4
    port map (
            O => \N__9937\,
            I => \DUT.uart_inst0.N_152_0\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__9932\,
            I => \DUT.uart_inst0.N_152_0\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__9925\,
            I => \DUT.uart_inst0.N_152_0\
        );

    \I__2048\ : InMux
    port map (
            O => \N__9910\,
            I => \N__9907\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__9907\,
            I => \N__9904\
        );

    \I__2046\ : Span4Mux_v
    port map (
            O => \N__9904\,
            I => \N__9900\
        );

    \I__2045\ : InMux
    port map (
            O => \N__9903\,
            I => \N__9897\
        );

    \I__2044\ : Span4Mux_h
    port map (
            O => \N__9900\,
            I => \N__9894\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__9897\,
            I => \DUT.uart_inst0.tx_dataZ0Z_3\
        );

    \I__2042\ : Odrv4
    port map (
            O => \N__9894\,
            I => \DUT.uart_inst0.tx_dataZ0Z_3\
        );

    \I__2041\ : InMux
    port map (
            O => \N__9889\,
            I => \N__9886\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__9886\,
            I => \N__9882\
        );

    \I__2039\ : InMux
    port map (
            O => \N__9885\,
            I => \N__9879\
        );

    \I__2038\ : Odrv4
    port map (
            O => \N__9882\,
            I => \DUT.uart_inst0.N_159\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__9879\,
            I => \DUT.uart_inst0.N_159\
        );

    \I__2036\ : CascadeMux
    port map (
            O => \N__9874\,
            I => \N__9871\
        );

    \I__2035\ : InMux
    port map (
            O => \N__9871\,
            I => \N__9867\
        );

    \I__2034\ : InMux
    port map (
            O => \N__9870\,
            I => \N__9864\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__9867\,
            I => \N__9861\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__9864\,
            I => \DUT.uart_inst0.tx_dataZ0Z_0\
        );

    \I__2031\ : Odrv4
    port map (
            O => \N__9861\,
            I => \DUT.uart_inst0.tx_dataZ0Z_0\
        );

    \I__2030\ : InMux
    port map (
            O => \N__9856\,
            I => \N__9852\
        );

    \I__2029\ : InMux
    port map (
            O => \N__9855\,
            I => \N__9846\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__9852\,
            I => \N__9843\
        );

    \I__2027\ : InMux
    port map (
            O => \N__9851\,
            I => \N__9839\
        );

    \I__2026\ : CascadeMux
    port map (
            O => \N__9850\,
            I => \N__9834\
        );

    \I__2025\ : InMux
    port map (
            O => \N__9849\,
            I => \N__9828\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__9846\,
            I => \N__9825\
        );

    \I__2023\ : Span4Mux_h
    port map (
            O => \N__9843\,
            I => \N__9822\
        );

    \I__2022\ : InMux
    port map (
            O => \N__9842\,
            I => \N__9819\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__9839\,
            I => \N__9816\
        );

    \I__2020\ : InMux
    port map (
            O => \N__9838\,
            I => \N__9813\
        );

    \I__2019\ : InMux
    port map (
            O => \N__9837\,
            I => \N__9804\
        );

    \I__2018\ : InMux
    port map (
            O => \N__9834\,
            I => \N__9804\
        );

    \I__2017\ : InMux
    port map (
            O => \N__9833\,
            I => \N__9804\
        );

    \I__2016\ : InMux
    port map (
            O => \N__9832\,
            I => \N__9804\
        );

    \I__2015\ : InMux
    port map (
            O => \N__9831\,
            I => \N__9801\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__9828\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__2013\ : Odrv4
    port map (
            O => \N__9825\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__2012\ : Odrv4
    port map (
            O => \N__9822\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__9819\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__2010\ : Odrv12
    port map (
            O => \N__9816\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__9813\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__9804\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__9801\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_1\
        );

    \I__2006\ : InMux
    port map (
            O => \N__9784\,
            I => \N__9781\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__9781\,
            I => \N__9778\
        );

    \I__2004\ : Span4Mux_h
    port map (
            O => \N__9778\,
            I => \N__9775\
        );

    \I__2003\ : Odrv4
    port map (
            O => \N__9775\,
            I => \DUT.uart_inst0.g0_i_a4_0_4\
        );

    \I__2002\ : InMux
    port map (
            O => \N__9772\,
            I => \N__9768\
        );

    \I__2001\ : InMux
    port map (
            O => \N__9771\,
            I => \N__9760\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__9768\,
            I => \N__9756\
        );

    \I__1999\ : InMux
    port map (
            O => \N__9767\,
            I => \N__9748\
        );

    \I__1998\ : InMux
    port map (
            O => \N__9766\,
            I => \N__9748\
        );

    \I__1997\ : CascadeMux
    port map (
            O => \N__9765\,
            I => \N__9745\
        );

    \I__1996\ : CascadeMux
    port map (
            O => \N__9764\,
            I => \N__9742\
        );

    \I__1995\ : InMux
    port map (
            O => \N__9763\,
            I => \N__9737\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__9760\,
            I => \N__9734\
        );

    \I__1993\ : InMux
    port map (
            O => \N__9759\,
            I => \N__9731\
        );

    \I__1992\ : Span4Mux_v
    port map (
            O => \N__9756\,
            I => \N__9728\
        );

    \I__1991\ : InMux
    port map (
            O => \N__9755\,
            I => \N__9725\
        );

    \I__1990\ : InMux
    port map (
            O => \N__9754\,
            I => \N__9720\
        );

    \I__1989\ : InMux
    port map (
            O => \N__9753\,
            I => \N__9720\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__9748\,
            I => \N__9717\
        );

    \I__1987\ : InMux
    port map (
            O => \N__9745\,
            I => \N__9708\
        );

    \I__1986\ : InMux
    port map (
            O => \N__9742\,
            I => \N__9708\
        );

    \I__1985\ : InMux
    port map (
            O => \N__9741\,
            I => \N__9708\
        );

    \I__1984\ : InMux
    port map (
            O => \N__9740\,
            I => \N__9708\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__9737\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__1982\ : Odrv4
    port map (
            O => \N__9734\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__9731\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__1980\ : Odrv4
    port map (
            O => \N__9728\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__9725\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__9720\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__1977\ : Odrv12
    port map (
            O => \N__9717\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__9708\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_0\
        );

    \I__1975\ : CascadeMux
    port map (
            O => \N__9691\,
            I => \DUT.uart_inst0.g0_i_a4_0_5_cascade_\
        );

    \I__1974\ : InMux
    port map (
            O => \N__9688\,
            I => \N__9685\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__9685\,
            I => \DUT.uart_inst0.N_15\
        );

    \I__1972\ : InMux
    port map (
            O => \N__9682\,
            I => \N__9679\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__9679\,
            I => \DUT.uart_inst0.N_7\
        );

    \I__1970\ : InMux
    port map (
            O => \N__9676\,
            I => \N__9667\
        );

    \I__1969\ : InMux
    port map (
            O => \N__9675\,
            I => \N__9664\
        );

    \I__1968\ : CascadeMux
    port map (
            O => \N__9674\,
            I => \N__9661\
        );

    \I__1967\ : CascadeMux
    port map (
            O => \N__9673\,
            I => \N__9653\
        );

    \I__1966\ : CascadeMux
    port map (
            O => \N__9672\,
            I => \N__9644\
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__9671\,
            I => \N__9639\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__9670\,
            I => \N__9636\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__9667\,
            I => \N__9631\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__9664\,
            I => \N__9631\
        );

    \I__1961\ : InMux
    port map (
            O => \N__9661\,
            I => \N__9628\
        );

    \I__1960\ : InMux
    port map (
            O => \N__9660\,
            I => \N__9621\
        );

    \I__1959\ : InMux
    port map (
            O => \N__9659\,
            I => \N__9621\
        );

    \I__1958\ : InMux
    port map (
            O => \N__9658\,
            I => \N__9621\
        );

    \I__1957\ : InMux
    port map (
            O => \N__9657\,
            I => \N__9612\
        );

    \I__1956\ : InMux
    port map (
            O => \N__9656\,
            I => \N__9612\
        );

    \I__1955\ : InMux
    port map (
            O => \N__9653\,
            I => \N__9612\
        );

    \I__1954\ : InMux
    port map (
            O => \N__9652\,
            I => \N__9612\
        );

    \I__1953\ : InMux
    port map (
            O => \N__9651\,
            I => \N__9599\
        );

    \I__1952\ : InMux
    port map (
            O => \N__9650\,
            I => \N__9599\
        );

    \I__1951\ : InMux
    port map (
            O => \N__9649\,
            I => \N__9599\
        );

    \I__1950\ : InMux
    port map (
            O => \N__9648\,
            I => \N__9599\
        );

    \I__1949\ : InMux
    port map (
            O => \N__9647\,
            I => \N__9599\
        );

    \I__1948\ : InMux
    port map (
            O => \N__9644\,
            I => \N__9599\
        );

    \I__1947\ : InMux
    port map (
            O => \N__9643\,
            I => \N__9590\
        );

    \I__1946\ : InMux
    port map (
            O => \N__9642\,
            I => \N__9590\
        );

    \I__1945\ : InMux
    port map (
            O => \N__9639\,
            I => \N__9590\
        );

    \I__1944\ : InMux
    port map (
            O => \N__9636\,
            I => \N__9590\
        );

    \I__1943\ : Odrv4
    port map (
            O => \N__9631\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__9628\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__9621\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__9612\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__9599\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__9590\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__9577\,
            I => \N__9574\
        );

    \I__1936\ : InMux
    port map (
            O => \N__9574\,
            I => \N__9571\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__9571\,
            I => \N__9568\
        );

    \I__1934\ : Span4Mux_h
    port map (
            O => \N__9568\,
            I => \N__9565\
        );

    \I__1933\ : Odrv4
    port map (
            O => \N__9565\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_3\
        );

    \I__1932\ : InMux
    port map (
            O => \N__9562\,
            I => \N__9559\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__9559\,
            I => \N__9556\
        );

    \I__1930\ : Odrv4
    port map (
            O => \N__9556\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3\
        );

    \I__1929\ : InMux
    port map (
            O => \N__9553\,
            I => \N__9550\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__9550\,
            I => \DUT.rFifoDatarx_3\
        );

    \I__1927\ : InMux
    port map (
            O => \N__9547\,
            I => \N__9544\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__9544\,
            I => \DUT.uart_inst0.tx_bits_remaining_RNO_1Z0Z_2\
        );

    \I__1925\ : InMux
    port map (
            O => \N__9541\,
            I => \N__9538\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__9538\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_9\
        );

    \I__1923\ : InMux
    port map (
            O => \N__9535\,
            I => \N__9532\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__9532\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_8\
        );

    \I__1921\ : InMux
    port map (
            O => \N__9529\,
            I => \N__9526\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__9526\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_7\
        );

    \I__1919\ : CascadeMux
    port map (
            O => \N__9523\,
            I => \N__9518\
        );

    \I__1918\ : InMux
    port map (
            O => \N__9522\,
            I => \N__9514\
        );

    \I__1917\ : CascadeMux
    port map (
            O => \N__9521\,
            I => \N__9510\
        );

    \I__1916\ : InMux
    port map (
            O => \N__9518\,
            I => \N__9506\
        );

    \I__1915\ : CascadeMux
    port map (
            O => \N__9517\,
            I => \N__9500\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__9514\,
            I => \N__9497\
        );

    \I__1913\ : InMux
    port map (
            O => \N__9513\,
            I => \N__9490\
        );

    \I__1912\ : InMux
    port map (
            O => \N__9510\,
            I => \N__9490\
        );

    \I__1911\ : InMux
    port map (
            O => \N__9509\,
            I => \N__9490\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__9506\,
            I => \N__9487\
        );

    \I__1909\ : InMux
    port map (
            O => \N__9505\,
            I => \N__9484\
        );

    \I__1908\ : InMux
    port map (
            O => \N__9504\,
            I => \N__9481\
        );

    \I__1907\ : InMux
    port map (
            O => \N__9503\,
            I => \N__9476\
        );

    \I__1906\ : InMux
    port map (
            O => \N__9500\,
            I => \N__9476\
        );

    \I__1905\ : Odrv4
    port map (
            O => \N__9497\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__9490\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__1903\ : Odrv12
    port map (
            O => \N__9487\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__9484\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__9481\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__9476\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_3\
        );

    \I__1899\ : CascadeMux
    port map (
            O => \N__9463\,
            I => \N__9458\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__9462\,
            I => \N__9453\
        );

    \I__1897\ : InMux
    port map (
            O => \N__9461\,
            I => \N__9446\
        );

    \I__1896\ : InMux
    port map (
            O => \N__9458\,
            I => \N__9446\
        );

    \I__1895\ : CascadeMux
    port map (
            O => \N__9457\,
            I => \N__9443\
        );

    \I__1894\ : CascadeMux
    port map (
            O => \N__9456\,
            I => \N__9440\
        );

    \I__1893\ : InMux
    port map (
            O => \N__9453\,
            I => \N__9437\
        );

    \I__1892\ : InMux
    port map (
            O => \N__9452\,
            I => \N__9434\
        );

    \I__1891\ : InMux
    port map (
            O => \N__9451\,
            I => \N__9431\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__9446\,
            I => \N__9428\
        );

    \I__1889\ : InMux
    port map (
            O => \N__9443\,
            I => \N__9425\
        );

    \I__1888\ : InMux
    port map (
            O => \N__9440\,
            I => \N__9422\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__9437\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_5\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__9434\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_5\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__9431\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_5\
        );

    \I__1884\ : Odrv4
    port map (
            O => \N__9428\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_5\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__9425\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_5\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__9422\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_5\
        );

    \I__1881\ : InMux
    port map (
            O => \N__9409\,
            I => \N__9406\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__9406\,
            I => \N__9396\
        );

    \I__1879\ : InMux
    port map (
            O => \N__9405\,
            I => \N__9387\
        );

    \I__1878\ : InMux
    port map (
            O => \N__9404\,
            I => \N__9387\
        );

    \I__1877\ : InMux
    port map (
            O => \N__9403\,
            I => \N__9387\
        );

    \I__1876\ : InMux
    port map (
            O => \N__9402\,
            I => \N__9387\
        );

    \I__1875\ : InMux
    port map (
            O => \N__9401\,
            I => \N__9382\
        );

    \I__1874\ : InMux
    port map (
            O => \N__9400\,
            I => \N__9379\
        );

    \I__1873\ : InMux
    port map (
            O => \N__9399\,
            I => \N__9376\
        );

    \I__1872\ : Span4Mux_h
    port map (
            O => \N__9396\,
            I => \N__9373\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__9387\,
            I => \N__9370\
        );

    \I__1870\ : InMux
    port map (
            O => \N__9386\,
            I => \N__9365\
        );

    \I__1869\ : InMux
    port map (
            O => \N__9385\,
            I => \N__9365\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__9382\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_2\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__9379\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_2\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__9376\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_2\
        );

    \I__1865\ : Odrv4
    port map (
            O => \N__9373\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_2\
        );

    \I__1864\ : Odrv4
    port map (
            O => \N__9370\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_2\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__9365\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_2\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__9352\,
            I => \DUT.uart_inst0.tx_data_i_m_4_0_cascade_\
        );

    \I__1861\ : InMux
    port map (
            O => \N__9349\,
            I => \N__9344\
        );

    \I__1860\ : InMux
    port map (
            O => \N__9348\,
            I => \N__9340\
        );

    \I__1859\ : InMux
    port map (
            O => \N__9347\,
            I => \N__9336\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__9344\,
            I => \N__9330\
        );

    \I__1857\ : InMux
    port map (
            O => \N__9343\,
            I => \N__9327\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__9340\,
            I => \N__9324\
        );

    \I__1855\ : InMux
    port map (
            O => \N__9339\,
            I => \N__9321\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__9336\,
            I => \N__9318\
        );

    \I__1853\ : InMux
    port map (
            O => \N__9335\,
            I => \N__9311\
        );

    \I__1852\ : InMux
    port map (
            O => \N__9334\,
            I => \N__9311\
        );

    \I__1851\ : InMux
    port map (
            O => \N__9333\,
            I => \N__9311\
        );

    \I__1850\ : Span4Mux_h
    port map (
            O => \N__9330\,
            I => \N__9308\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__9327\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_4\
        );

    \I__1848\ : Odrv4
    port map (
            O => \N__9324\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_4\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__9321\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_4\
        );

    \I__1846\ : Odrv4
    port map (
            O => \N__9318\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_4\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__9311\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_4\
        );

    \I__1844\ : Odrv4
    port map (
            O => \N__9308\,
            I => \DUT.uart_inst0.tx_countdownZ0Z_4\
        );

    \I__1843\ : CascadeMux
    port map (
            O => \N__9295\,
            I => \N__9292\
        );

    \I__1842\ : InMux
    port map (
            O => \N__9292\,
            I => \N__9288\
        );

    \I__1841\ : InMux
    port map (
            O => \N__9291\,
            I => \N__9285\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__9288\,
            I => \N__9282\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__9285\,
            I => \DUT.uart_inst0.tx_countdown_0_c4_i\
        );

    \I__1838\ : Odrv4
    port map (
            O => \N__9282\,
            I => \DUT.uart_inst0.tx_countdown_0_c4_i\
        );

    \I__1837\ : InMux
    port map (
            O => \N__9277\,
            I => \N__9274\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__9274\,
            I => \DUT.uart_inst0.tx_state_ns_0_o3_1_0_1\
        );

    \I__1835\ : InMux
    port map (
            O => \N__9271\,
            I => \N__9268\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__9268\,
            I => \N__9265\
        );

    \I__1833\ : Span4Mux_v
    port map (
            O => \N__9265\,
            I => \N__9261\
        );

    \I__1832\ : InMux
    port map (
            O => \N__9264\,
            I => \N__9258\
        );

    \I__1831\ : Odrv4
    port map (
            O => \N__9261\,
            I => \G_148\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__9258\,
            I => \G_148\
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__9253\,
            I => \fifo_inst.ftdi_output_inst.N_95_cascade_\
        );

    \I__1828\ : InMux
    port map (
            O => \N__9250\,
            I => \N__9246\
        );

    \I__1827\ : InMux
    port map (
            O => \N__9249\,
            I => \N__9243\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__9246\,
            I => \N__9240\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__9243\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_3\
        );

    \I__1824\ : Odrv4
    port map (
            O => \N__9240\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_3\
        );

    \I__1823\ : InMux
    port map (
            O => \N__9235\,
            I => \N__9232\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__9232\,
            I => \N__9229\
        );

    \I__1821\ : Span4Mux_h
    port map (
            O => \N__9229\,
            I => \N__9225\
        );

    \I__1820\ : InMux
    port map (
            O => \N__9228\,
            I => \N__9222\
        );

    \I__1819\ : Odrv4
    port map (
            O => \N__9225\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__9222\,
            I => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2\
        );

    \I__1817\ : InMux
    port map (
            O => \N__9217\,
            I => \N__9214\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__9214\,
            I => \fifo_inst.ftdi_output_inst.N_95\
        );

    \I__1815\ : CascadeMux
    port map (
            O => \N__9211\,
            I => \fifo_inst.ftdi_output_inst.m14_1_cascade_\
        );

    \I__1814\ : InMux
    port map (
            O => \N__9208\,
            I => \N__9202\
        );

    \I__1813\ : InMux
    port map (
            O => \N__9207\,
            I => \N__9202\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__9202\,
            I => \fifo_inst.ftdi_output_inst.N_86_0\
        );

    \I__1811\ : CascadeMux
    port map (
            O => \N__9199\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_9_cascade_\
        );

    \I__1810\ : InMux
    port map (
            O => \N__9196\,
            I => \N__9193\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__9193\,
            I => \N__9189\
        );

    \I__1808\ : InMux
    port map (
            O => \N__9192\,
            I => \N__9186\
        );

    \I__1807\ : Odrv4
    port map (
            O => \N__9189\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_13\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__9186\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_13\
        );

    \I__1805\ : InMux
    port map (
            O => \N__9181\,
            I => \N__9177\
        );

    \I__1804\ : InMux
    port map (
            O => \N__9180\,
            I => \N__9174\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__9177\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_5\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__9174\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_5\
        );

    \I__1801\ : CascadeMux
    port map (
            O => \N__9169\,
            I => \N__9166\
        );

    \I__1800\ : InMux
    port map (
            O => \N__9166\,
            I => \N__9162\
        );

    \I__1799\ : InMux
    port map (
            O => \N__9165\,
            I => \N__9158\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__9162\,
            I => \N__9155\
        );

    \I__1797\ : InMux
    port map (
            O => \N__9161\,
            I => \N__9152\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__9158\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_5\
        );

    \I__1795\ : Odrv4
    port map (
            O => \N__9155\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_5\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__9152\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_5\
        );

    \I__1793\ : InMux
    port map (
            O => \N__9145\,
            I => \N__9137\
        );

    \I__1792\ : InMux
    port map (
            O => \N__9144\,
            I => \N__9137\
        );

    \I__1791\ : InMux
    port map (
            O => \N__9143\,
            I => \N__9132\
        );

    \I__1790\ : InMux
    port map (
            O => \N__9142\,
            I => \N__9132\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__9137\,
            I => \N__9124\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__9132\,
            I => \N__9121\
        );

    \I__1787\ : InMux
    port map (
            O => \N__9131\,
            I => \N__9116\
        );

    \I__1786\ : InMux
    port map (
            O => \N__9130\,
            I => \N__9116\
        );

    \I__1785\ : InMux
    port map (
            O => \N__9129\,
            I => \N__9111\
        );

    \I__1784\ : InMux
    port map (
            O => \N__9128\,
            I => \N__9111\
        );

    \I__1783\ : InMux
    port map (
            O => \N__9127\,
            I => \N__9108\
        );

    \I__1782\ : Odrv4
    port map (
            O => \N__9124\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__1781\ : Odrv4
    port map (
            O => \N__9121\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__9116\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__9111\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__9108\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0\
        );

    \I__1777\ : CascadeMux
    port map (
            O => \N__9097\,
            I => \N__9094\
        );

    \I__1776\ : InMux
    port map (
            O => \N__9094\,
            I => \N__9087\
        );

    \I__1775\ : InMux
    port map (
            O => \N__9093\,
            I => \N__9087\
        );

    \I__1774\ : InMux
    port map (
            O => \N__9092\,
            I => \N__9084\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__9087\,
            I => \N__9081\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__9084\,
            I => \N__9078\
        );

    \I__1771\ : Span4Mux_h
    port map (
            O => \N__9081\,
            I => \N__9075\
        );

    \I__1770\ : Odrv4
    port map (
            O => \N__9078\,
            I => \DUT.uart_inst0.N_70\
        );

    \I__1769\ : Odrv4
    port map (
            O => \N__9075\,
            I => \DUT.uart_inst0.N_70\
        );

    \I__1768\ : InMux
    port map (
            O => \N__9070\,
            I => \N__9063\
        );

    \I__1767\ : InMux
    port map (
            O => \N__9069\,
            I => \N__9063\
        );

    \I__1766\ : InMux
    port map (
            O => \N__9068\,
            I => \N__9059\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__9063\,
            I => \N__9056\
        );

    \I__1764\ : InMux
    port map (
            O => \N__9062\,
            I => \N__9053\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__9059\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__1762\ : Odrv12
    port map (
            O => \N__9056\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__9053\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_3\
        );

    \I__1760\ : InMux
    port map (
            O => \N__9046\,
            I => \N__9042\
        );

    \I__1759\ : InMux
    port map (
            O => \N__9045\,
            I => \N__9039\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__9042\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_11\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__9039\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_11\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__9034\,
            I => \N__9031\
        );

    \I__1755\ : InMux
    port map (
            O => \N__9031\,
            I => \N__9027\
        );

    \I__1754\ : InMux
    port map (
            O => \N__9030\,
            I => \N__9024\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__9027\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_12\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__9024\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_12\
        );

    \I__1751\ : InMux
    port map (
            O => \N__9019\,
            I => \N__9016\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__9016\,
            I => \N__9013\
        );

    \I__1749\ : Odrv4
    port map (
            O => \N__9013\,
            I => \DUT.rFifoDatarx_5\
        );

    \I__1748\ : CascadeMux
    port map (
            O => \N__9010\,
            I => \DUT.uart_inst0.tx_data_RNO_0Z0Z_5_cascade_\
        );

    \I__1747\ : InMux
    port map (
            O => \N__9007\,
            I => \N__9003\
        );

    \I__1746\ : InMux
    port map (
            O => \N__9006\,
            I => \N__9000\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__9003\,
            I => \N__8997\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__9000\,
            I => \DUT.uart_inst0.tx_dataZ0Z_5\
        );

    \I__1743\ : Odrv4
    port map (
            O => \N__8997\,
            I => \DUT.uart_inst0.tx_dataZ0Z_5\
        );

    \I__1742\ : InMux
    port map (
            O => \N__8992\,
            I => \N__8988\
        );

    \I__1741\ : InMux
    port map (
            O => \N__8991\,
            I => \N__8985\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__8988\,
            I => \N__8978\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__8985\,
            I => \N__8978\
        );

    \I__1738\ : InMux
    port map (
            O => \N__8984\,
            I => \N__8975\
        );

    \I__1737\ : InMux
    port map (
            O => \N__8983\,
            I => \N__8972\
        );

    \I__1736\ : Span4Mux_h
    port map (
            O => \N__8978\,
            I => \N__8967\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__8975\,
            I => \N__8967\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__8972\,
            I => \N__8964\
        );

    \I__1733\ : Span4Mux_v
    port map (
            O => \N__8967\,
            I => \N__8961\
        );

    \I__1732\ : Span4Mux_h
    port map (
            O => \N__8964\,
            I => \N__8958\
        );

    \I__1731\ : Span4Mux_v
    port map (
            O => \N__8961\,
            I => \N__8955\
        );

    \I__1730\ : Span4Mux_v
    port map (
            O => \N__8958\,
            I => \N__8952\
        );

    \I__1729\ : Odrv4
    port map (
            O => \N__8955\,
            I => \rTxByteZ0Z_1\
        );

    \I__1728\ : Odrv4
    port map (
            O => \N__8952\,
            I => \rTxByteZ0Z_1\
        );

    \I__1727\ : InMux
    port map (
            O => \N__8947\,
            I => \N__8944\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__8944\,
            I => \N__8941\
        );

    \I__1725\ : Odrv4
    port map (
            O => \N__8941\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_1\
        );

    \I__1724\ : InMux
    port map (
            O => \N__8938\,
            I => \N__8934\
        );

    \I__1723\ : InMux
    port map (
            O => \N__8937\,
            I => \N__8930\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__8934\,
            I => \N__8926\
        );

    \I__1721\ : InMux
    port map (
            O => \N__8933\,
            I => \N__8923\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__8930\,
            I => \N__8920\
        );

    \I__1719\ : InMux
    port map (
            O => \N__8929\,
            I => \N__8917\
        );

    \I__1718\ : Span4Mux_v
    port map (
            O => \N__8926\,
            I => \N__8914\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__8923\,
            I => \N__8911\
        );

    \I__1716\ : Span4Mux_v
    port map (
            O => \N__8920\,
            I => \N__8906\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__8917\,
            I => \N__8906\
        );

    \I__1714\ : Span4Mux_v
    port map (
            O => \N__8914\,
            I => \N__8903\
        );

    \I__1713\ : Span12Mux_v
    port map (
            O => \N__8911\,
            I => \N__8900\
        );

    \I__1712\ : Span4Mux_v
    port map (
            O => \N__8906\,
            I => \N__8897\
        );

    \I__1711\ : Odrv4
    port map (
            O => \N__8903\,
            I => \rTxByteZ0Z_0\
        );

    \I__1710\ : Odrv12
    port map (
            O => \N__8900\,
            I => \rTxByteZ0Z_0\
        );

    \I__1709\ : Odrv4
    port map (
            O => \N__8897\,
            I => \rTxByteZ0Z_0\
        );

    \I__1708\ : InMux
    port map (
            O => \N__8890\,
            I => \N__8887\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__8887\,
            I => \N__8884\
        );

    \I__1706\ : Span4Mux_v
    port map (
            O => \N__8884\,
            I => \N__8881\
        );

    \I__1705\ : Odrv4
    port map (
            O => \N__8881\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_0\
        );

    \I__1704\ : InMux
    port map (
            O => \N__8878\,
            I => \N__8873\
        );

    \I__1703\ : InMux
    port map (
            O => \N__8877\,
            I => \N__8870\
        );

    \I__1702\ : InMux
    port map (
            O => \N__8876\,
            I => \N__8867\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__8873\,
            I => \N__8863\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8870\,
            I => \N__8858\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__8867\,
            I => \N__8858\
        );

    \I__1698\ : InMux
    port map (
            O => \N__8866\,
            I => \N__8855\
        );

    \I__1697\ : Span4Mux_v
    port map (
            O => \N__8863\,
            I => \N__8852\
        );

    \I__1696\ : Span4Mux_h
    port map (
            O => \N__8858\,
            I => \N__8847\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__8855\,
            I => \N__8847\
        );

    \I__1694\ : Span4Mux_v
    port map (
            O => \N__8852\,
            I => \N__8844\
        );

    \I__1693\ : Span4Mux_v
    port map (
            O => \N__8847\,
            I => \N__8841\
        );

    \I__1692\ : Odrv4
    port map (
            O => \N__8844\,
            I => \rTxByteZ0Z_6\
        );

    \I__1691\ : Odrv4
    port map (
            O => \N__8841\,
            I => \rTxByteZ0Z_6\
        );

    \I__1690\ : InMux
    port map (
            O => \N__8836\,
            I => \N__8833\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__8833\,
            I => \N__8830\
        );

    \I__1688\ : Odrv4
    port map (
            O => \N__8830\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_6\
        );

    \I__1687\ : InMux
    port map (
            O => \N__8827\,
            I => \N__8824\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__8824\,
            I => \DUT.uart_inst0.tx_data_8_321_a2_0\
        );

    \I__1685\ : CascadeMux
    port map (
            O => \N__8821\,
            I => \DUT.uart_inst0.tx_countdown_0_1_5_cascade_\
        );

    \I__1684\ : InMux
    port map (
            O => \N__8818\,
            I => \N__8815\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__8815\,
            I => \DUT.uart_inst0.g0_i_o4_0_5\
        );

    \I__1682\ : CascadeMux
    port map (
            O => \N__8812\,
            I => \DUT.uart_inst0.N_14_cascade_\
        );

    \I__1681\ : IoInMux
    port map (
            O => \N__8809\,
            I => \N__8806\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__8806\,
            I => \N__8803\
        );

    \I__1679\ : Span4Mux_s1_v
    port map (
            O => \N__8803\,
            I => \N__8800\
        );

    \I__1678\ : Sp12to4
    port map (
            O => \N__8800\,
            I => \N__8797\
        );

    \I__1677\ : Span12Mux_h
    port map (
            O => \N__8797\,
            I => \N__8793\
        );

    \I__1676\ : CascadeMux
    port map (
            O => \N__8796\,
            I => \N__8790\
        );

    \I__1675\ : Span12Mux_v
    port map (
            O => \N__8793\,
            I => \N__8787\
        );

    \I__1674\ : InMux
    port map (
            O => \N__8790\,
            I => \N__8784\
        );

    \I__1673\ : Odrv12
    port map (
            O => \N__8787\,
            I => \P1A7_c\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__8784\,
            I => \P1A7_c\
        );

    \I__1671\ : InMux
    port map (
            O => \N__8779\,
            I => \N__8776\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__8776\,
            I => \DUT.uart_inst0.N_6\
        );

    \I__1669\ : InMux
    port map (
            O => \N__8773\,
            I => \N__8770\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__8770\,
            I => \N__8767\
        );

    \I__1667\ : Odrv4
    port map (
            O => \N__8767\,
            I => \DUT.uart_inst0.un1_tx_bits_remaining_axbxc2_N_4L5_1_0\
        );

    \I__1666\ : InMux
    port map (
            O => \N__8764\,
            I => \N__8761\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__8761\,
            I => \N__8758\
        );

    \I__1664\ : Odrv4
    port map (
            O => \N__8758\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1\
        );

    \I__1663\ : CascadeMux
    port map (
            O => \N__8755\,
            I => \N__8752\
        );

    \I__1662\ : InMux
    port map (
            O => \N__8752\,
            I => \N__8749\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__8749\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_1\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__8746\,
            I => \N__8743\
        );

    \I__1659\ : InMux
    port map (
            O => \N__8743\,
            I => \N__8740\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__8740\,
            I => \N__8736\
        );

    \I__1657\ : InMux
    port map (
            O => \N__8739\,
            I => \N__8733\
        );

    \I__1656\ : Odrv4
    port map (
            O => \N__8736\,
            I => \DUT.uart_inst0.tx_dataZ0Z_2\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__8733\,
            I => \DUT.uart_inst0.tx_dataZ0Z_2\
        );

    \I__1654\ : CascadeMux
    port map (
            O => \N__8728\,
            I => \DUT.rFifoDatarx_1_cascade_\
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__8725\,
            I => \DUT.uart_inst0.tx_data_RNO_0Z0Z_1_cascade_\
        );

    \I__1652\ : InMux
    port map (
            O => \N__8722\,
            I => \N__8719\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__8719\,
            I => \N__8715\
        );

    \I__1650\ : InMux
    port map (
            O => \N__8718\,
            I => \N__8712\
        );

    \I__1649\ : Odrv4
    port map (
            O => \N__8715\,
            I => \DUT.uart_inst0.tx_dataZ0Z_1\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__8712\,
            I => \DUT.uart_inst0.tx_dataZ0Z_1\
        );

    \I__1647\ : InMux
    port map (
            O => \N__8707\,
            I => \N__8704\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__8704\,
            I => \DUT.uart_inst0.tx_data_RNO_0Z0Z_0\
        );

    \I__1645\ : CascadeMux
    port map (
            O => \N__8701\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_6_cascade_\
        );

    \I__1644\ : InMux
    port map (
            O => \N__8698\,
            I => \N__8695\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__8695\,
            I => \DUT.uart_inst0.un1_tx_bits_remaining_axbxc2_N_4L5_1_1\
        );

    \I__1642\ : CascadeMux
    port map (
            O => \N__8692\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_0_cascade_\
        );

    \I__1641\ : InMux
    port map (
            O => \N__8689\,
            I => \N__8686\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__8686\,
            I => \DUT.uart_inst0.un1_tx_bits_remaining_axbxc2_N_4L5_1\
        );

    \I__1639\ : InMux
    port map (
            O => \N__8683\,
            I => \N__8677\
        );

    \I__1638\ : InMux
    port map (
            O => \N__8682\,
            I => \N__8670\
        );

    \I__1637\ : CascadeMux
    port map (
            O => \N__8681\,
            I => \N__8667\
        );

    \I__1636\ : CascadeMux
    port map (
            O => \N__8680\,
            I => \N__8664\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__8677\,
            I => \N__8661\
        );

    \I__1634\ : InMux
    port map (
            O => \N__8676\,
            I => \N__8658\
        );

    \I__1633\ : InMux
    port map (
            O => \N__8675\,
            I => \N__8651\
        );

    \I__1632\ : InMux
    port map (
            O => \N__8674\,
            I => \N__8651\
        );

    \I__1631\ : InMux
    port map (
            O => \N__8673\,
            I => \N__8651\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__8670\,
            I => \N__8648\
        );

    \I__1629\ : InMux
    port map (
            O => \N__8667\,
            I => \N__8643\
        );

    \I__1628\ : InMux
    port map (
            O => \N__8664\,
            I => \N__8643\
        );

    \I__1627\ : Span4Mux_h
    port map (
            O => \N__8661\,
            I => \N__8636\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__8658\,
            I => \N__8636\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__8651\,
            I => \N__8636\
        );

    \I__1624\ : Odrv4
    port map (
            O => \N__8648\,
            I => \rRxReadZ0\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__8643\,
            I => \rRxReadZ0\
        );

    \I__1622\ : Odrv4
    port map (
            O => \N__8636\,
            I => \rRxReadZ0\
        );

    \I__1621\ : CascadeMux
    port map (
            O => \N__8629\,
            I => \N__8626\
        );

    \I__1620\ : InMux
    port map (
            O => \N__8626\,
            I => \N__8623\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__8623\,
            I => \N__8617\
        );

    \I__1618\ : InMux
    port map (
            O => \N__8622\,
            I => \N__8614\
        );

    \I__1617\ : InMux
    port map (
            O => \N__8621\,
            I => \N__8609\
        );

    \I__1616\ : InMux
    port map (
            O => \N__8620\,
            I => \N__8609\
        );

    \I__1615\ : Odrv4
    port map (
            O => \N__8617\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_1\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__8614\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_1\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__8609\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_1\
        );

    \I__1612\ : CascadeMux
    port map (
            O => \N__8602\,
            I => \N__8599\
        );

    \I__1611\ : InMux
    port map (
            O => \N__8599\,
            I => \N__8596\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__8596\,
            I => \N__8593\
        );

    \I__1609\ : Odrv4
    port map (
            O => \N__8593\,
            I => \DUT.fifo_tx_inst.rFifoCount_RNIBPFMZ0Z_1\
        );

    \I__1608\ : CascadeMux
    port map (
            O => \N__8590\,
            I => \DUT.uart_inst0.g0_0_0_a3_3_cascade_\
        );

    \I__1607\ : CascadeMux
    port map (
            O => \N__8587\,
            I => \DUT.uart_inst0.g0_0_0_a3_5_cascade_\
        );

    \I__1606\ : InMux
    port map (
            O => \N__8584\,
            I => \N__8581\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__8581\,
            I => \DUT.uart_inst0.N_159_0_0\
        );

    \I__1604\ : InMux
    port map (
            O => \N__8578\,
            I => \N__8570\
        );

    \I__1603\ : InMux
    port map (
            O => \N__8577\,
            I => \N__8570\
        );

    \I__1602\ : InMux
    port map (
            O => \N__8576\,
            I => \N__8565\
        );

    \I__1601\ : InMux
    port map (
            O => \N__8575\,
            I => \N__8565\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__8570\,
            I => \N__8562\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__8565\,
            I => \N__8559\
        );

    \I__1598\ : Odrv12
    port map (
            O => \N__8562\,
            I => \DUT.N_37\
        );

    \I__1597\ : Odrv4
    port map (
            O => \N__8559\,
            I => \DUT.N_37\
        );

    \I__1596\ : InMux
    port map (
            O => \N__8554\,
            I => \N__8551\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__8551\,
            I => \N__8548\
        );

    \I__1594\ : Odrv4
    port map (
            O => \N__8548\,
            I => \DUT.uart_inst0.N_105\
        );

    \I__1593\ : InMux
    port map (
            O => \N__8545\,
            I => \N__8541\
        );

    \I__1592\ : CascadeMux
    port map (
            O => \N__8544\,
            I => \N__8537\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__8541\,
            I => \N__8534\
        );

    \I__1590\ : InMux
    port map (
            O => \N__8540\,
            I => \N__8531\
        );

    \I__1589\ : InMux
    port map (
            O => \N__8537\,
            I => \N__8528\
        );

    \I__1588\ : Odrv4
    port map (
            O => \N__8534\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_1\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__8531\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_1\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__8528\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_1\
        );

    \I__1585\ : InMux
    port map (
            O => \N__8521\,
            I => \N__8518\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__8518\,
            I => \N__8515\
        );

    \I__1583\ : Odrv4
    port map (
            O => \N__8515\,
            I => \DUT.uart_inst0.N_102\
        );

    \I__1582\ : CascadeMux
    port map (
            O => \N__8512\,
            I => \N__8509\
        );

    \I__1581\ : InMux
    port map (
            O => \N__8509\,
            I => \N__8505\
        );

    \I__1580\ : CascadeMux
    port map (
            O => \N__8508\,
            I => \N__8501\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__8505\,
            I => \N__8498\
        );

    \I__1578\ : InMux
    port map (
            O => \N__8504\,
            I => \N__8495\
        );

    \I__1577\ : InMux
    port map (
            O => \N__8501\,
            I => \N__8492\
        );

    \I__1576\ : Odrv4
    port map (
            O => \N__8498\,
            I => \DUT.uart_inst0.rx_countdownZ1Z_3\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__8495\,
            I => \DUT.uart_inst0.rx_countdownZ1Z_3\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__8492\,
            I => \DUT.uart_inst0.rx_countdownZ1Z_3\
        );

    \I__1573\ : InMux
    port map (
            O => \N__8485\,
            I => \N__8482\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__8482\,
            I => \N__8479\
        );

    \I__1571\ : Odrv4
    port map (
            O => \N__8479\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_1_1_2\
        );

    \I__1570\ : InMux
    port map (
            O => \N__8476\,
            I => \N__8472\
        );

    \I__1569\ : InMux
    port map (
            O => \N__8475\,
            I => \N__8469\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__8472\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_4\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__8469\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_4\
        );

    \I__1566\ : CascadeMux
    port map (
            O => \N__8464\,
            I => \N__8460\
        );

    \I__1565\ : CascadeMux
    port map (
            O => \N__8463\,
            I => \N__8456\
        );

    \I__1564\ : InMux
    port map (
            O => \N__8460\,
            I => \N__8451\
        );

    \I__1563\ : InMux
    port map (
            O => \N__8459\,
            I => \N__8451\
        );

    \I__1562\ : InMux
    port map (
            O => \N__8456\,
            I => \N__8448\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__8451\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_4\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__8448\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_4\
        );

    \I__1559\ : InMux
    port map (
            O => \N__8443\,
            I => \N__8440\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__8440\,
            I => \N__8437\
        );

    \I__1557\ : Span4Mux_h
    port map (
            O => \N__8437\,
            I => \N__8434\
        );

    \I__1556\ : Odrv4
    port map (
            O => \N__8434\,
            I => \DUT.uart_inst0.rx_countdown_RNO_0Z0Z_2\
        );

    \I__1555\ : InMux
    port map (
            O => \N__8431\,
            I => \N__8427\
        );

    \I__1554\ : InMux
    port map (
            O => \N__8430\,
            I => \N__8423\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__8427\,
            I => \N__8420\
        );

    \I__1552\ : InMux
    port map (
            O => \N__8426\,
            I => \N__8412\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__8423\,
            I => \N__8409\
        );

    \I__1550\ : Span4Mux_h
    port map (
            O => \N__8420\,
            I => \N__8406\
        );

    \I__1549\ : InMux
    port map (
            O => \N__8419\,
            I => \N__8401\
        );

    \I__1548\ : InMux
    port map (
            O => \N__8418\,
            I => \N__8401\
        );

    \I__1547\ : InMux
    port map (
            O => \N__8417\,
            I => \N__8394\
        );

    \I__1546\ : InMux
    port map (
            O => \N__8416\,
            I => \N__8394\
        );

    \I__1545\ : InMux
    port map (
            O => \N__8415\,
            I => \N__8394\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__8412\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_1_2\
        );

    \I__1543\ : Odrv4
    port map (
            O => \N__8409\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_1_2\
        );

    \I__1542\ : Odrv4
    port map (
            O => \N__8406\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_1_2\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__8401\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_1_2\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__8394\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_1_2\
        );

    \I__1539\ : CascadeMux
    port map (
            O => \N__8383\,
            I => \N__8380\
        );

    \I__1538\ : InMux
    port map (
            O => \N__8380\,
            I => \N__8377\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__8377\,
            I => \N__8374\
        );

    \I__1536\ : Odrv4
    port map (
            O => \N__8374\,
            I => \DUT.uart_inst0.rx_countdown_RNO_1Z0Z_2\
        );

    \I__1535\ : InMux
    port map (
            O => \N__8371\,
            I => \N__8363\
        );

    \I__1534\ : InMux
    port map (
            O => \N__8370\,
            I => \N__8360\
        );

    \I__1533\ : CascadeMux
    port map (
            O => \N__8369\,
            I => \N__8356\
        );

    \I__1532\ : CascadeMux
    port map (
            O => \N__8368\,
            I => \N__8352\
        );

    \I__1531\ : CascadeMux
    port map (
            O => \N__8367\,
            I => \N__8349\
        );

    \I__1530\ : InMux
    port map (
            O => \N__8366\,
            I => \N__8346\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__8363\,
            I => \N__8343\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__8360\,
            I => \N__8340\
        );

    \I__1527\ : InMux
    port map (
            O => \N__8359\,
            I => \N__8337\
        );

    \I__1526\ : InMux
    port map (
            O => \N__8356\,
            I => \N__8332\
        );

    \I__1525\ : InMux
    port map (
            O => \N__8355\,
            I => \N__8332\
        );

    \I__1524\ : InMux
    port map (
            O => \N__8352\,
            I => \N__8327\
        );

    \I__1523\ : InMux
    port map (
            O => \N__8349\,
            I => \N__8327\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__8346\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_2_2\
        );

    \I__1521\ : Odrv4
    port map (
            O => \N__8343\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_2_2\
        );

    \I__1520\ : Odrv4
    port map (
            O => \N__8340\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_2_2\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__8337\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_2_2\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__8332\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_2_2\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__8327\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_2_2\
        );

    \I__1516\ : InMux
    port map (
            O => \N__8314\,
            I => \N__8310\
        );

    \I__1515\ : CascadeMux
    port map (
            O => \N__8313\,
            I => \N__8307\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__8310\,
            I => \N__8304\
        );

    \I__1513\ : InMux
    port map (
            O => \N__8307\,
            I => \N__8301\
        );

    \I__1512\ : Span4Mux_h
    port map (
            O => \N__8304\,
            I => \N__8296\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__8301\,
            I => \N__8296\
        );

    \I__1510\ : Odrv4
    port map (
            O => \N__8296\,
            I => \DUT.uart_inst0.rx_countdownZ0Z_2\
        );

    \I__1509\ : CascadeMux
    port map (
            O => \N__8293\,
            I => \N__8285\
        );

    \I__1508\ : InMux
    port map (
            O => \N__8292\,
            I => \N__8280\
        );

    \I__1507\ : InMux
    port map (
            O => \N__8291\,
            I => \N__8280\
        );

    \I__1506\ : InMux
    port map (
            O => \N__8290\,
            I => \N__8275\
        );

    \I__1505\ : InMux
    port map (
            O => \N__8289\,
            I => \N__8275\
        );

    \I__1504\ : InMux
    port map (
            O => \N__8288\,
            I => \N__8270\
        );

    \I__1503\ : InMux
    port map (
            O => \N__8285\,
            I => \N__8270\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__8280\,
            I => \DUT.uart_inst0.recv_stateZ0Z_5\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__8275\,
            I => \DUT.uart_inst0.recv_stateZ0Z_5\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__8270\,
            I => \DUT.uart_inst0.recv_stateZ0Z_5\
        );

    \I__1499\ : InMux
    port map (
            O => \N__8263\,
            I => \N__8258\
        );

    \I__1498\ : InMux
    port map (
            O => \N__8262\,
            I => \N__8255\
        );

    \I__1497\ : InMux
    port map (
            O => \N__8261\,
            I => \N__8252\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__8258\,
            I => \N__8249\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__8255\,
            I => \DUT.uart_inst0.recv_stateZ0Z_3\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__8252\,
            I => \DUT.uart_inst0.recv_stateZ0Z_3\
        );

    \I__1493\ : Odrv4
    port map (
            O => \N__8249\,
            I => \DUT.uart_inst0.recv_stateZ0Z_3\
        );

    \I__1492\ : InMux
    port map (
            O => \N__8242\,
            I => \N__8233\
        );

    \I__1491\ : InMux
    port map (
            O => \N__8241\,
            I => \N__8233\
        );

    \I__1490\ : CascadeMux
    port map (
            O => \N__8240\,
            I => \N__8230\
        );

    \I__1489\ : CascadeMux
    port map (
            O => \N__8239\,
            I => \N__8225\
        );

    \I__1488\ : InMux
    port map (
            O => \N__8238\,
            I => \N__8220\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__8233\,
            I => \N__8217\
        );

    \I__1486\ : InMux
    port map (
            O => \N__8230\,
            I => \N__8214\
        );

    \I__1485\ : InMux
    port map (
            O => \N__8229\,
            I => \N__8211\
        );

    \I__1484\ : InMux
    port map (
            O => \N__8228\,
            I => \N__8206\
        );

    \I__1483\ : InMux
    port map (
            O => \N__8225\,
            I => \N__8206\
        );

    \I__1482\ : InMux
    port map (
            O => \N__8224\,
            I => \N__8203\
        );

    \I__1481\ : InMux
    port map (
            O => \N__8223\,
            I => \N__8200\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__8220\,
            I => \N__8197\
        );

    \I__1479\ : Span4Mux_h
    port map (
            O => \N__8217\,
            I => \N__8184\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__8214\,
            I => \N__8184\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__8211\,
            I => \N__8184\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__8206\,
            I => \N__8184\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__8203\,
            I => \N__8184\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__8200\,
            I => \N__8184\
        );

    \I__1473\ : Span4Mux_v
    port map (
            O => \N__8197\,
            I => \N__8180\
        );

    \I__1472\ : Span4Mux_v
    port map (
            O => \N__8184\,
            I => \N__8177\
        );

    \I__1471\ : InMux
    port map (
            O => \N__8183\,
            I => \N__8174\
        );

    \I__1470\ : Sp12to4
    port map (
            O => \N__8180\,
            I => \N__8167\
        );

    \I__1469\ : Sp12to4
    port map (
            O => \N__8177\,
            I => \N__8167\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__8174\,
            I => \N__8167\
        );

    \I__1467\ : Span12Mux_h
    port map (
            O => \N__8167\,
            I => \N__8164\
        );

    \I__1466\ : Span12Mux_v
    port map (
            O => \N__8164\,
            I => \N__8161\
        );

    \I__1465\ : Odrv12
    port map (
            O => \N__8161\,
            I => \P1A1_c\
        );

    \I__1464\ : InMux
    port map (
            O => \N__8158\,
            I => \N__8147\
        );

    \I__1463\ : InMux
    port map (
            O => \N__8157\,
            I => \N__8142\
        );

    \I__1462\ : InMux
    port map (
            O => \N__8156\,
            I => \N__8142\
        );

    \I__1461\ : InMux
    port map (
            O => \N__8155\,
            I => \N__8139\
        );

    \I__1460\ : InMux
    port map (
            O => \N__8154\,
            I => \N__8132\
        );

    \I__1459\ : InMux
    port map (
            O => \N__8153\,
            I => \N__8132\
        );

    \I__1458\ : InMux
    port map (
            O => \N__8152\,
            I => \N__8132\
        );

    \I__1457\ : InMux
    port map (
            O => \N__8151\,
            I => \N__8127\
        );

    \I__1456\ : InMux
    port map (
            O => \N__8150\,
            I => \N__8127\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__8147\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__8142\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__8139\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__8132\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__8127\,
            I => \DUT.uart_inst0.recv_stateZ0Z_1\
        );

    \I__1450\ : InMux
    port map (
            O => \N__8116\,
            I => \N__8113\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__8113\,
            I => \N__8110\
        );

    \I__1448\ : Odrv4
    port map (
            O => \N__8110\,
            I => \DUT.uart_inst0.recv_state_srsts_1_5\
        );

    \I__1447\ : InMux
    port map (
            O => \N__8107\,
            I => \N__8104\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__8104\,
            I => \N__8100\
        );

    \I__1445\ : InMux
    port map (
            O => \N__8103\,
            I => \N__8097\
        );

    \I__1444\ : Odrv4
    port map (
            O => \N__8100\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_1\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__8097\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_1\
        );

    \I__1442\ : InMux
    port map (
            O => \N__8092\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_0_s1\
        );

    \I__1441\ : InMux
    port map (
            O => \N__8089\,
            I => \N__8086\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__8086\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_1_s1_THRU_CO\
        );

    \I__1439\ : InMux
    port map (
            O => \N__8083\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_1_s1\
        );

    \I__1438\ : InMux
    port map (
            O => \N__8080\,
            I => \N__8074\
        );

    \I__1437\ : InMux
    port map (
            O => \N__8079\,
            I => \N__8074\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__8074\,
            I => \DUT.uart_inst0.rx_countdown_3_s1_3\
        );

    \I__1435\ : InMux
    port map (
            O => \N__8071\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_2_s1\
        );

    \I__1434\ : InMux
    port map (
            O => \N__8068\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_3_s1\
        );

    \I__1433\ : InMux
    port map (
            O => \N__8065\,
            I => \DUT.uart_inst0.rx_countdown_3_cry_4_s1\
        );

    \I__1432\ : CascadeMux
    port map (
            O => \N__8062\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_10_cascade_\
        );

    \I__1431\ : CascadeMux
    port map (
            O => \N__8059\,
            I => \N__8056\
        );

    \I__1430\ : InMux
    port map (
            O => \N__8056\,
            I => \N__8053\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__8053\,
            I => \DUT.uart_inst0.rx_clk_divider_RNIKU472Z0Z_10\
        );

    \I__1428\ : InMux
    port map (
            O => \N__8050\,
            I => \N__8047\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__8047\,
            I => \DUT.uart_inst0.recv_state_RNO_0Z0Z_0\
        );

    \I__1426\ : CascadeMux
    port map (
            O => \N__8044\,
            I => \DUT.uart_inst0.recv_state_RNO_1Z0Z_0_cascade_\
        );

    \I__1425\ : InMux
    port map (
            O => \N__8041\,
            I => \N__8031\
        );

    \I__1424\ : InMux
    port map (
            O => \N__8040\,
            I => \N__8031\
        );

    \I__1423\ : InMux
    port map (
            O => \N__8039\,
            I => \N__8031\
        );

    \I__1422\ : InMux
    port map (
            O => \N__8038\,
            I => \N__8028\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__8031\,
            I => \DUT.uart_inst0.recv_stateZ0Z_0\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__8028\,
            I => \DUT.uart_inst0.recv_stateZ0Z_0\
        );

    \I__1419\ : InMux
    port map (
            O => \N__8023\,
            I => \N__8020\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__8020\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_a_10\
        );

    \I__1417\ : CascadeMux
    port map (
            O => \N__8017\,
            I => \DUT.uart_inst0.un2_rx_clk_divider_0_cascade_\
        );

    \I__1416\ : InMux
    port map (
            O => \N__8014\,
            I => \N__8004\
        );

    \I__1415\ : InMux
    port map (
            O => \N__8013\,
            I => \N__8001\
        );

    \I__1414\ : InMux
    port map (
            O => \N__8012\,
            I => \N__7998\
        );

    \I__1413\ : InMux
    port map (
            O => \N__8011\,
            I => \N__7993\
        );

    \I__1412\ : InMux
    port map (
            O => \N__8010\,
            I => \N__7993\
        );

    \I__1411\ : InMux
    port map (
            O => \N__8009\,
            I => \N__7986\
        );

    \I__1410\ : InMux
    port map (
            O => \N__8008\,
            I => \N__7986\
        );

    \I__1409\ : InMux
    port map (
            O => \N__8007\,
            I => \N__7986\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__8004\,
            I => \DUT.uart_inst0.rx_countdown_3_2\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__8001\,
            I => \DUT.uart_inst0.rx_countdown_3_2\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__7998\,
            I => \DUT.uart_inst0.rx_countdown_3_2\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__7993\,
            I => \DUT.uart_inst0.rx_countdown_3_2\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__7986\,
            I => \DUT.uart_inst0.rx_countdown_3_2\
        );

    \I__1403\ : CascadeMux
    port map (
            O => \N__7975\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_1_2_cascade_\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__7972\,
            I => \DUT.uart_inst0.recv_state_RNO_0Z0Z_4_cascade_\
        );

    \I__1401\ : InMux
    port map (
            O => \N__7969\,
            I => \N__7966\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__7966\,
            I => \N__7962\
        );

    \I__1399\ : InMux
    port map (
            O => \N__7965\,
            I => \N__7959\
        );

    \I__1398\ : Odrv4
    port map (
            O => \N__7962\,
            I => \DUT.uart_inst0.recv_stateZ0Z_4\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__7959\,
            I => \DUT.uart_inst0.recv_stateZ0Z_4\
        );

    \I__1396\ : InMux
    port map (
            O => \N__7954\,
            I => \N__7951\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__7951\,
            I => \N__7948\
        );

    \I__1394\ : Odrv4
    port map (
            O => \N__7948\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_6\
        );

    \I__1393\ : InMux
    port map (
            O => \N__7945\,
            I => \N__7941\
        );

    \I__1392\ : InMux
    port map (
            O => \N__7944\,
            I => \N__7938\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__7941\,
            I => \N__7933\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__7938\,
            I => \N__7930\
        );

    \I__1389\ : InMux
    port map (
            O => \N__7937\,
            I => \N__7927\
        );

    \I__1388\ : InMux
    port map (
            O => \N__7936\,
            I => \N__7924\
        );

    \I__1387\ : Span4Mux_h
    port map (
            O => \N__7933\,
            I => \N__7915\
        );

    \I__1386\ : Span4Mux_h
    port map (
            O => \N__7930\,
            I => \N__7915\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__7927\,
            I => \N__7915\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__7924\,
            I => \N__7915\
        );

    \I__1383\ : Sp12to4
    port map (
            O => \N__7915\,
            I => \N__7912\
        );

    \I__1382\ : Odrv12
    port map (
            O => \N__7912\,
            I => \rTxByteZ0Z_7\
        );

    \I__1381\ : InMux
    port map (
            O => \N__7909\,
            I => \N__7906\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__7906\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_7\
        );

    \I__1379\ : CEMux
    port map (
            O => \N__7903\,
            I => \N__7900\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__7900\,
            I => \N__7897\
        );

    \I__1377\ : Span4Mux_h
    port map (
            O => \N__7897\,
            I => \N__7893\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7896\,
            I => \N__7890\
        );

    \I__1375\ : Odrv4
    port map (
            O => \N__7893\,
            I => \DUT.fifo_tx_inst.rFifoData_awe3\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__7890\,
            I => \DUT.fifo_tx_inst.rFifoData_awe3\
        );

    \I__1373\ : InMux
    port map (
            O => \N__7885\,
            I => \N__7882\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__7882\,
            I => \DUT.rFifoDatarx_7\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__7879\,
            I => \G_152_cascade_\
        );

    \I__1370\ : CascadeMux
    port map (
            O => \N__7876\,
            I => \N__7873\
        );

    \I__1369\ : InMux
    port map (
            O => \N__7873\,
            I => \N__7870\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__7870\,
            I => \N__7865\
        );

    \I__1367\ : InMux
    port map (
            O => \N__7869\,
            I => \N__7860\
        );

    \I__1366\ : InMux
    port map (
            O => \N__7868\,
            I => \N__7860\
        );

    \I__1365\ : Odrv12
    port map (
            O => \N__7865\,
            I => \G_151\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__7860\,
            I => \G_151\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__7855\,
            I => \N__7852\
        );

    \I__1362\ : InMux
    port map (
            O => \N__7852\,
            I => \N__7849\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__7849\,
            I => \N__7844\
        );

    \I__1360\ : InMux
    port map (
            O => \N__7848\,
            I => \N__7839\
        );

    \I__1359\ : InMux
    port map (
            O => \N__7847\,
            I => \N__7839\
        );

    \I__1358\ : Odrv12
    port map (
            O => \N__7844\,
            I => \G_150\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__7839\,
            I => \G_150\
        );

    \I__1356\ : InMux
    port map (
            O => \N__7834\,
            I => \N__7829\
        );

    \I__1355\ : InMux
    port map (
            O => \N__7833\,
            I => \N__7824\
        );

    \I__1354\ : InMux
    port map (
            O => \N__7832\,
            I => \N__7824\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__7829\,
            I => \fifo_inst.ftdi_input_inst.un1_rWrStateZ0Z_1\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__7824\,
            I => \fifo_inst.ftdi_input_inst.un1_rWrStateZ0Z_1\
        );

    \I__1351\ : CascadeMux
    port map (
            O => \N__7819\,
            I => \N__7816\
        );

    \I__1350\ : InMux
    port map (
            O => \N__7816\,
            I => \N__7813\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__7813\,
            I => \N__7807\
        );

    \I__1348\ : InMux
    port map (
            O => \N__7812\,
            I => \N__7800\
        );

    \I__1347\ : InMux
    port map (
            O => \N__7811\,
            I => \N__7800\
        );

    \I__1346\ : InMux
    port map (
            O => \N__7810\,
            I => \N__7800\
        );

    \I__1345\ : Odrv12
    port map (
            O => \N__7807\,
            I => \G_149\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__7800\,
            I => \G_149\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7795\,
            I => \N__7792\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__7792\,
            I => \fifo_inst.ftdi_input_inst.un2_oPacketAvail_iZ0\
        );

    \I__1341\ : CascadeMux
    port map (
            O => \N__7789\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_\
        );

    \I__1340\ : InMux
    port map (
            O => \N__7786\,
            I => \N__7783\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__7783\,
            I => \DUT.uart_inst0.tx_data_RNO_0Z0Z_2\
        );

    \I__1338\ : InMux
    port map (
            O => \N__7780\,
            I => \N__7777\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__7777\,
            I => \N__7774\
        );

    \I__1336\ : Odrv4
    port map (
            O => \N__7774\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_0\
        );

    \I__1335\ : InMux
    port map (
            O => \N__7771\,
            I => \N__7768\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__7768\,
            I => \N__7763\
        );

    \I__1333\ : InMux
    port map (
            O => \N__7767\,
            I => \N__7760\
        );

    \I__1332\ : InMux
    port map (
            O => \N__7766\,
            I => \N__7757\
        );

    \I__1331\ : Span4Mux_h
    port map (
            O => \N__7763\,
            I => \N__7751\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__7760\,
            I => \N__7751\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__7757\,
            I => \N__7748\
        );

    \I__1328\ : InMux
    port map (
            O => \N__7756\,
            I => \N__7745\
        );

    \I__1327\ : Span4Mux_v
    port map (
            O => \N__7751\,
            I => \N__7742\
        );

    \I__1326\ : Span4Mux_v
    port map (
            O => \N__7748\,
            I => \N__7737\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__7745\,
            I => \N__7737\
        );

    \I__1324\ : Span4Mux_v
    port map (
            O => \N__7742\,
            I => \N__7734\
        );

    \I__1323\ : Span4Mux_v
    port map (
            O => \N__7737\,
            I => \N__7731\
        );

    \I__1322\ : Odrv4
    port map (
            O => \N__7734\,
            I => \rTxByteZ0Z_2\
        );

    \I__1321\ : Odrv4
    port map (
            O => \N__7731\,
            I => \rTxByteZ0Z_2\
        );

    \I__1320\ : InMux
    port map (
            O => \N__7726\,
            I => \N__7723\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__7723\,
            I => \N__7720\
        );

    \I__1318\ : Odrv4
    port map (
            O => \N__7720\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_2\
        );

    \I__1317\ : InMux
    port map (
            O => \N__7717\,
            I => \N__7712\
        );

    \I__1316\ : InMux
    port map (
            O => \N__7716\,
            I => \N__7709\
        );

    \I__1315\ : InMux
    port map (
            O => \N__7715\,
            I => \N__7706\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__7712\,
            I => \N__7702\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__7709\,
            I => \N__7697\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__7706\,
            I => \N__7697\
        );

    \I__1311\ : InMux
    port map (
            O => \N__7705\,
            I => \N__7694\
        );

    \I__1310\ : Span4Mux_v
    port map (
            O => \N__7702\,
            I => \N__7691\
        );

    \I__1309\ : Span4Mux_v
    port map (
            O => \N__7697\,
            I => \N__7686\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__7694\,
            I => \N__7686\
        );

    \I__1307\ : Span4Mux_v
    port map (
            O => \N__7691\,
            I => \N__7683\
        );

    \I__1306\ : Span4Mux_v
    port map (
            O => \N__7686\,
            I => \N__7680\
        );

    \I__1305\ : Odrv4
    port map (
            O => \N__7683\,
            I => \rTxByteZ0Z_4\
        );

    \I__1304\ : Odrv4
    port map (
            O => \N__7680\,
            I => \rTxByteZ0Z_4\
        );

    \I__1303\ : CascadeMux
    port map (
            O => \N__7675\,
            I => \N__7672\
        );

    \I__1302\ : InMux
    port map (
            O => \N__7672\,
            I => \N__7669\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__7669\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_4\
        );

    \I__1300\ : InMux
    port map (
            O => \N__7666\,
            I => \N__7663\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__7663\,
            I => \N__7657\
        );

    \I__1298\ : InMux
    port map (
            O => \N__7662\,
            I => \N__7654\
        );

    \I__1297\ : InMux
    port map (
            O => \N__7661\,
            I => \N__7651\
        );

    \I__1296\ : InMux
    port map (
            O => \N__7660\,
            I => \N__7648\
        );

    \I__1295\ : Span4Mux_h
    port map (
            O => \N__7657\,
            I => \N__7639\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__7654\,
            I => \N__7639\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__7651\,
            I => \N__7639\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__7648\,
            I => \N__7639\
        );

    \I__1291\ : Span4Mux_v
    port map (
            O => \N__7639\,
            I => \N__7636\
        );

    \I__1290\ : Odrv4
    port map (
            O => \N__7636\,
            I => \rTxByteZ0Z_5\
        );

    \I__1289\ : InMux
    port map (
            O => \N__7633\,
            I => \N__7630\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__7630\,
            I => \N__7627\
        );

    \I__1287\ : Odrv4
    port map (
            O => \N__7627\,
            I => \DUT.fifo_tx_inst.rFifoData_ram3_5\
        );

    \I__1286\ : CascadeMux
    port map (
            O => \N__7624\,
            I => \DUT.uart_inst0.g0_i_o4_0_4_cascade_\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__7621\,
            I => \N__7616\
        );

    \I__1284\ : InMux
    port map (
            O => \N__7620\,
            I => \N__7613\
        );

    \I__1283\ : InMux
    port map (
            O => \N__7619\,
            I => \N__7605\
        );

    \I__1282\ : InMux
    port map (
            O => \N__7616\,
            I => \N__7602\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__7613\,
            I => \N__7599\
        );

    \I__1280\ : InMux
    port map (
            O => \N__7612\,
            I => \N__7596\
        );

    \I__1279\ : InMux
    port map (
            O => \N__7611\,
            I => \N__7591\
        );

    \I__1278\ : InMux
    port map (
            O => \N__7610\,
            I => \N__7591\
        );

    \I__1277\ : InMux
    port map (
            O => \N__7609\,
            I => \N__7588\
        );

    \I__1276\ : InMux
    port map (
            O => \N__7608\,
            I => \N__7585\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__7605\,
            I => \N__7582\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__7602\,
            I => \N__7575\
        );

    \I__1273\ : Span4Mux_v
    port map (
            O => \N__7599\,
            I => \N__7575\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__7596\,
            I => \N__7575\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__7591\,
            I => \N__7569\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__7588\,
            I => \N__7569\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__7585\,
            I => \N__7564\
        );

    \I__1268\ : Span4Mux_v
    port map (
            O => \N__7582\,
            I => \N__7564\
        );

    \I__1267\ : Span4Mux_v
    port map (
            O => \N__7575\,
            I => \N__7561\
        );

    \I__1266\ : InMux
    port map (
            O => \N__7574\,
            I => \N__7558\
        );

    \I__1265\ : Odrv12
    port map (
            O => \N__7569\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_1\
        );

    \I__1264\ : Odrv4
    port map (
            O => \N__7564\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_1\
        );

    \I__1263\ : Odrv4
    port map (
            O => \N__7561\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_1\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__7558\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_1\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__7549\,
            I => \N__7542\
        );

    \I__1260\ : InMux
    port map (
            O => \N__7548\,
            I => \N__7538\
        );

    \I__1259\ : CascadeMux
    port map (
            O => \N__7547\,
            I => \N__7535\
        );

    \I__1258\ : CascadeMux
    port map (
            O => \N__7546\,
            I => \N__7532\
        );

    \I__1257\ : InMux
    port map (
            O => \N__7545\,
            I => \N__7529\
        );

    \I__1256\ : InMux
    port map (
            O => \N__7542\,
            I => \N__7525\
        );

    \I__1255\ : InMux
    port map (
            O => \N__7541\,
            I => \N__7522\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__7538\,
            I => \N__7519\
        );

    \I__1253\ : InMux
    port map (
            O => \N__7535\,
            I => \N__7514\
        );

    \I__1252\ : InMux
    port map (
            O => \N__7532\,
            I => \N__7514\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__7529\,
            I => \N__7511\
        );

    \I__1250\ : InMux
    port map (
            O => \N__7528\,
            I => \N__7508\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__7525\,
            I => \N__7505\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__7522\,
            I => \N__7497\
        );

    \I__1247\ : Span4Mux_v
    port map (
            O => \N__7519\,
            I => \N__7497\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__7514\,
            I => \N__7488\
        );

    \I__1245\ : Span4Mux_v
    port map (
            O => \N__7511\,
            I => \N__7488\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__7508\,
            I => \N__7488\
        );

    \I__1243\ : Span4Mux_h
    port map (
            O => \N__7505\,
            I => \N__7488\
        );

    \I__1242\ : InMux
    port map (
            O => \N__7504\,
            I => \N__7481\
        );

    \I__1241\ : InMux
    port map (
            O => \N__7503\,
            I => \N__7481\
        );

    \I__1240\ : InMux
    port map (
            O => \N__7502\,
            I => \N__7481\
        );

    \I__1239\ : Odrv4
    port map (
            O => \N__7497\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_0\
        );

    \I__1238\ : Odrv4
    port map (
            O => \N__7488\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_0\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__7481\,
            I => \DUT.fifo_tx_inst.rWritePtrZ0Z_0\
        );

    \I__1236\ : InMux
    port map (
            O => \N__7474\,
            I => \N__7467\
        );

    \I__1235\ : InMux
    port map (
            O => \N__7473\,
            I => \N__7464\
        );

    \I__1234\ : InMux
    port map (
            O => \N__7472\,
            I => \N__7457\
        );

    \I__1233\ : InMux
    port map (
            O => \N__7471\,
            I => \N__7457\
        );

    \I__1232\ : InMux
    port map (
            O => \N__7470\,
            I => \N__7457\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__7467\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_2\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__7464\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_2\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__7457\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_2\
        );

    \I__1228\ : InMux
    port map (
            O => \N__7450\,
            I => \N__7447\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__7447\,
            I => \DUT.rFifoDatarxZ0Z_0\
        );

    \I__1226\ : InMux
    port map (
            O => \N__7444\,
            I => \N__7441\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__7441\,
            I => \N__7438\
        );

    \I__1224\ : Span4Mux_h
    port map (
            O => \N__7438\,
            I => \N__7435\
        );

    \I__1223\ : Odrv4
    port map (
            O => \N__7435\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_4\
        );

    \I__1222\ : InMux
    port map (
            O => \N__7432\,
            I => \N__7429\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__7429\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4\
        );

    \I__1220\ : CascadeMux
    port map (
            O => \N__7426\,
            I => \DUT.rFifoDatarx_4_cascade_\
        );

    \I__1219\ : InMux
    port map (
            O => \N__7423\,
            I => \N__7420\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__7420\,
            I => \DUT.uart_inst0.tx_data_RNO_0Z0Z_4\
        );

    \I__1217\ : InMux
    port map (
            O => \N__7417\,
            I => \N__7414\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__7414\,
            I => \N__7411\
        );

    \I__1215\ : Span4Mux_v
    port map (
            O => \N__7411\,
            I => \N__7408\
        );

    \I__1214\ : Odrv4
    port map (
            O => \N__7408\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_6\
        );

    \I__1213\ : CascadeMux
    port map (
            O => \N__7405\,
            I => \N__7402\
        );

    \I__1212\ : InMux
    port map (
            O => \N__7402\,
            I => \N__7399\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__7399\,
            I => \N__7396\
        );

    \I__1210\ : Odrv4
    port map (
            O => \N__7396\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_6\
        );

    \I__1209\ : CascadeMux
    port map (
            O => \N__7393\,
            I => \N__7387\
        );

    \I__1208\ : InMux
    port map (
            O => \N__7392\,
            I => \N__7377\
        );

    \I__1207\ : InMux
    port map (
            O => \N__7391\,
            I => \N__7374\
        );

    \I__1206\ : InMux
    port map (
            O => \N__7390\,
            I => \N__7367\
        );

    \I__1205\ : InMux
    port map (
            O => \N__7387\,
            I => \N__7367\
        );

    \I__1204\ : InMux
    port map (
            O => \N__7386\,
            I => \N__7367\
        );

    \I__1203\ : InMux
    port map (
            O => \N__7385\,
            I => \N__7362\
        );

    \I__1202\ : InMux
    port map (
            O => \N__7384\,
            I => \N__7362\
        );

    \I__1201\ : InMux
    port map (
            O => \N__7383\,
            I => \N__7353\
        );

    \I__1200\ : InMux
    port map (
            O => \N__7382\,
            I => \N__7353\
        );

    \I__1199\ : InMux
    port map (
            O => \N__7381\,
            I => \N__7353\
        );

    \I__1198\ : InMux
    port map (
            O => \N__7380\,
            I => \N__7353\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__7377\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__7374\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__7367\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__7362\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__7353\,
            I => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\
        );

    \I__1192\ : InMux
    port map (
            O => \N__7342\,
            I => \N__7339\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__7339\,
            I => \DUT.uart_inst0.tx_countdown_0_c3\
        );

    \I__1190\ : InMux
    port map (
            O => \N__7336\,
            I => \N__7333\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__7333\,
            I => \DUT.uart_inst0.un1_m7_3\
        );

    \I__1188\ : CascadeMux
    port map (
            O => \N__7330\,
            I => \DUT.uart_inst0.un1_tx_state_0_a4_1_cascade_\
        );

    \I__1187\ : CascadeMux
    port map (
            O => \N__7327\,
            I => \DUT.uart_inst0.un1_tx_clk_divider_s1_sn_0_cascade_\
        );

    \I__1186\ : InMux
    port map (
            O => \N__7324\,
            I => \N__7321\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__7321\,
            I => \DUT.uart_inst0.tx_countdown_7_1_0_3\
        );

    \I__1184\ : CascadeMux
    port map (
            O => \N__7318\,
            I => \DUT.uart_inst0.tx_countdown_RNO_0Z0Z_1_cascade_\
        );

    \I__1183\ : CascadeMux
    port map (
            O => \N__7315\,
            I => \DUT.uart_inst0.N_98_4_cascade_\
        );

    \I__1182\ : InMux
    port map (
            O => \N__7312\,
            I => \N__7308\
        );

    \I__1181\ : InMux
    port map (
            O => \N__7311\,
            I => \N__7305\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__7308\,
            I => \N__7302\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__7305\,
            I => \DUT.uart_inst0.rx_m2_e_0\
        );

    \I__1178\ : Odrv4
    port map (
            O => \N__7302\,
            I => \DUT.uart_inst0.rx_m2_e_0\
        );

    \I__1177\ : CascadeMux
    port map (
            O => \N__7297\,
            I => \DUT.uart_inst0.r_N_5_mux_cascade_\
        );

    \I__1176\ : InMux
    port map (
            O => \N__7294\,
            I => \N__7281\
        );

    \I__1175\ : InMux
    port map (
            O => \N__7293\,
            I => \N__7281\
        );

    \I__1174\ : InMux
    port map (
            O => \N__7292\,
            I => \N__7281\
        );

    \I__1173\ : InMux
    port map (
            O => \N__7291\,
            I => \N__7281\
        );

    \I__1172\ : InMux
    port map (
            O => \N__7290\,
            I => \N__7278\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__7281\,
            I => \DUT.uart_inst0.recv_stateZ0Z_2\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__7278\,
            I => \DUT.uart_inst0.recv_stateZ0Z_2\
        );

    \I__1169\ : InMux
    port map (
            O => \N__7273\,
            I => \N__7270\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__7270\,
            I => \DUT.uart_inst0.N_98_4\
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__7267\,
            I => \DUT.uart_inst0.r_N_3_mux_cascade_\
        );

    \I__1166\ : InMux
    port map (
            O => \N__7264\,
            I => \N__7258\
        );

    \I__1165\ : InMux
    port map (
            O => \N__7263\,
            I => \N__7258\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__7258\,
            I => \DUT.uart_inst0.recv_N_5_mux\
        );

    \I__1163\ : CascadeMux
    port map (
            O => \N__7255\,
            I => \DUT.uart_inst0.g3_cascade_\
        );

    \I__1162\ : CascadeMux
    port map (
            O => \N__7252\,
            I => \N__7249\
        );

    \I__1161\ : InMux
    port map (
            O => \N__7249\,
            I => \N__7246\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__7246\,
            I => \DUT.uart_inst0.g3_1\
        );

    \I__1159\ : CascadeMux
    port map (
            O => \N__7243\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_2_2_cascade_\
        );

    \I__1158\ : CascadeMux
    port map (
            O => \N__7240\,
            I => \DUT.uart_inst0.recv_state_RNO_0Z0Z_1_cascade_\
        );

    \I__1157\ : CascadeMux
    port map (
            O => \N__7237\,
            I => \DUT.uart_inst0.un1_m2_e_0_cascade_\
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__7234\,
            I => \N__7230\
        );

    \I__1155\ : InMux
    port map (
            O => \N__7233\,
            I => \N__7227\
        );

    \I__1154\ : InMux
    port map (
            O => \N__7230\,
            I => \N__7224\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__7227\,
            I => \N__7221\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__7224\,
            I => \DUT.uart_inst0.N_69\
        );

    \I__1151\ : Odrv4
    port map (
            O => \N__7221\,
            I => \DUT.uart_inst0.N_69\
        );

    \I__1150\ : CascadeMux
    port map (
            O => \N__7216\,
            I => \DUT.uart_inst0.recv_state_RNITN8GJZ0Z_2_cascade_\
        );

    \I__1149\ : CEMux
    port map (
            O => \N__7213\,
            I => \N__7210\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__7210\,
            I => \N__7207\
        );

    \I__1147\ : Span4Mux_h
    port map (
            O => \N__7207\,
            I => \N__7203\
        );

    \I__1146\ : InMux
    port map (
            O => \N__7206\,
            I => \N__7200\
        );

    \I__1145\ : Odrv4
    port map (
            O => \N__7203\,
            I => \DUT.uart_inst0.recv_state_RNITN8GJZ0Z_2\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__7200\,
            I => \DUT.uart_inst0.recv_state_RNITN8GJZ0Z_2\
        );

    \I__1143\ : InMux
    port map (
            O => \N__7195\,
            I => \N__7190\
        );

    \I__1142\ : InMux
    port map (
            O => \N__7194\,
            I => \N__7187\
        );

    \I__1141\ : InMux
    port map (
            O => \N__7193\,
            I => \N__7184\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__7190\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_2\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__7187\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_2\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__7184\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_2\
        );

    \I__1137\ : InMux
    port map (
            O => \N__7177\,
            I => \N__7173\
        );

    \I__1136\ : CascadeMux
    port map (
            O => \N__7176\,
            I => \N__7170\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__7173\,
            I => \N__7166\
        );

    \I__1134\ : InMux
    port map (
            O => \N__7170\,
            I => \N__7161\
        );

    \I__1133\ : InMux
    port map (
            O => \N__7169\,
            I => \N__7161\
        );

    \I__1132\ : Odrv4
    port map (
            O => \N__7166\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_1\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__7161\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_1\
        );

    \I__1130\ : CascadeMux
    port map (
            O => \N__7156\,
            I => \N__7153\
        );

    \I__1129\ : InMux
    port map (
            O => \N__7153\,
            I => \N__7149\
        );

    \I__1128\ : InMux
    port map (
            O => \N__7152\,
            I => \N__7146\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__7149\,
            I => \N__7143\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__7146\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_3\
        );

    \I__1125\ : Odrv4
    port map (
            O => \N__7143\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_3\
        );

    \I__1124\ : InMux
    port map (
            O => \N__7138\,
            I => \N__7132\
        );

    \I__1123\ : InMux
    port map (
            O => \N__7137\,
            I => \N__7127\
        );

    \I__1122\ : InMux
    port map (
            O => \N__7136\,
            I => \N__7127\
        );

    \I__1121\ : InMux
    port map (
            O => \N__7135\,
            I => \N__7124\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__7132\,
            I => \N__7119\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__7127\,
            I => \N__7119\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__7124\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_0\
        );

    \I__1117\ : Odrv4
    port map (
            O => \N__7119\,
            I => \DUT.uart_inst0.rx_bits_remainingZ0Z_0\
        );

    \I__1116\ : CEMux
    port map (
            O => \N__7114\,
            I => \N__7111\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__7111\,
            I => \N__7108\
        );

    \I__1114\ : Odrv12
    port map (
            O => \N__7108\,
            I => \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa\
        );

    \I__1113\ : CascadeMux
    port map (
            O => \N__7105\,
            I => \DUT.uart_inst0.rx_countdown_3_2_cascade_\
        );

    \I__1112\ : CascadeMux
    port map (
            O => \N__7102\,
            I => \N__7097\
        );

    \I__1111\ : InMux
    port map (
            O => \N__7101\,
            I => \N__7094\
        );

    \I__1110\ : InMux
    port map (
            O => \N__7100\,
            I => \N__7088\
        );

    \I__1109\ : InMux
    port map (
            O => \N__7097\,
            I => \N__7085\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__7094\,
            I => \N__7082\
        );

    \I__1107\ : InMux
    port map (
            O => \N__7093\,
            I => \N__7079\
        );

    \I__1106\ : InMux
    port map (
            O => \N__7092\,
            I => \N__7074\
        );

    \I__1105\ : InMux
    port map (
            O => \N__7091\,
            I => \N__7074\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__7088\,
            I => \DUT.wRcvd\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__7085\,
            I => \DUT.wRcvd\
        );

    \I__1102\ : Odrv4
    port map (
            O => \N__7082\,
            I => \DUT.wRcvd\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__7079\,
            I => \DUT.wRcvd\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__7074\,
            I => \DUT.wRcvd\
        );

    \I__1099\ : CascadeMux
    port map (
            O => \N__7063\,
            I => \DUT.uart_inst0.rx_countdown_8_i_o2_2_1_2_cascade_\
        );

    \I__1098\ : CascadeMux
    port map (
            O => \N__7060\,
            I => \N__7057\
        );

    \I__1097\ : InMux
    port map (
            O => \N__7057\,
            I => \N__7054\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__7054\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_7\
        );

    \I__1095\ : CEMux
    port map (
            O => \N__7051\,
            I => \N__7048\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__7048\,
            I => \N__7045\
        );

    \I__1093\ : Span4Mux_h
    port map (
            O => \N__7045\,
            I => \N__7042\
        );

    \I__1092\ : Span4Mux_h
    port map (
            O => \N__7042\,
            I => \N__7039\
        );

    \I__1091\ : Odrv4
    port map (
            O => \N__7039\,
            I => \DUT.fifo_rx_inst.rFifoData_awe1\
        );

    \I__1090\ : InMux
    port map (
            O => \N__7036\,
            I => \N__7033\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__7033\,
            I => \N__7028\
        );

    \I__1088\ : InMux
    port map (
            O => \N__7032\,
            I => \N__7025\
        );

    \I__1087\ : InMux
    port map (
            O => \N__7031\,
            I => \N__7021\
        );

    \I__1086\ : Span4Mux_v
    port map (
            O => \N__7028\,
            I => \N__7016\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__7025\,
            I => \N__7016\
        );

    \I__1084\ : InMux
    port map (
            O => \N__7024\,
            I => \N__7013\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__7021\,
            I => \DUT.wRxByte_0\
        );

    \I__1082\ : Odrv4
    port map (
            O => \N__7016\,
            I => \DUT.wRxByte_0\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__7013\,
            I => \DUT.wRxByte_0\
        );

    \I__1080\ : InMux
    port map (
            O => \N__7006\,
            I => \N__7003\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__7003\,
            I => \N__6998\
        );

    \I__1078\ : InMux
    port map (
            O => \N__7002\,
            I => \N__6995\
        );

    \I__1077\ : InMux
    port map (
            O => \N__7001\,
            I => \N__6990\
        );

    \I__1076\ : Span4Mux_v
    port map (
            O => \N__6998\,
            I => \N__6985\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__6995\,
            I => \N__6985\
        );

    \I__1074\ : InMux
    port map (
            O => \N__6994\,
            I => \N__6982\
        );

    \I__1073\ : InMux
    port map (
            O => \N__6993\,
            I => \N__6979\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__6990\,
            I => \DUT.wRxByte_1\
        );

    \I__1071\ : Odrv4
    port map (
            O => \N__6985\,
            I => \DUT.wRxByte_1\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__6982\,
            I => \DUT.wRxByte_1\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__6979\,
            I => \DUT.wRxByte_1\
        );

    \I__1068\ : InMux
    port map (
            O => \N__6970\,
            I => \N__6967\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__6967\,
            I => \N__6962\
        );

    \I__1066\ : InMux
    port map (
            O => \N__6966\,
            I => \N__6959\
        );

    \I__1065\ : InMux
    port map (
            O => \N__6965\,
            I => \N__6956\
        );

    \I__1064\ : Span4Mux_h
    port map (
            O => \N__6962\,
            I => \N__6951\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__6959\,
            I => \N__6946\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__6956\,
            I => \N__6946\
        );

    \I__1061\ : InMux
    port map (
            O => \N__6955\,
            I => \N__6943\
        );

    \I__1060\ : InMux
    port map (
            O => \N__6954\,
            I => \N__6940\
        );

    \I__1059\ : Odrv4
    port map (
            O => \N__6951\,
            I => \DUT.wRxByte_2\
        );

    \I__1058\ : Odrv4
    port map (
            O => \N__6946\,
            I => \DUT.wRxByte_2\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__6943\,
            I => \DUT.wRxByte_2\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__6940\,
            I => \DUT.wRxByte_2\
        );

    \I__1055\ : InMux
    port map (
            O => \N__6931\,
            I => \N__6927\
        );

    \I__1054\ : InMux
    port map (
            O => \N__6930\,
            I => \N__6924\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__6927\,
            I => \N__6920\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__6924\,
            I => \N__6917\
        );

    \I__1051\ : InMux
    port map (
            O => \N__6923\,
            I => \N__6914\
        );

    \I__1050\ : Span4Mux_h
    port map (
            O => \N__6920\,
            I => \N__6909\
        );

    \I__1049\ : Span4Mux_v
    port map (
            O => \N__6917\,
            I => \N__6904\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__6914\,
            I => \N__6904\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6913\,
            I => \N__6901\
        );

    \I__1046\ : InMux
    port map (
            O => \N__6912\,
            I => \N__6898\
        );

    \I__1045\ : Odrv4
    port map (
            O => \N__6909\,
            I => \DUT.wRxByte_3\
        );

    \I__1044\ : Odrv4
    port map (
            O => \N__6904\,
            I => \DUT.wRxByte_3\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__6901\,
            I => \DUT.wRxByte_3\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__6898\,
            I => \DUT.wRxByte_3\
        );

    \I__1041\ : InMux
    port map (
            O => \N__6889\,
            I => \N__6885\
        );

    \I__1040\ : InMux
    port map (
            O => \N__6888\,
            I => \N__6882\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__6885\,
            I => \N__6878\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__6882\,
            I => \N__6875\
        );

    \I__1037\ : InMux
    port map (
            O => \N__6881\,
            I => \N__6872\
        );

    \I__1036\ : Span4Mux_v
    port map (
            O => \N__6878\,
            I => \N__6863\
        );

    \I__1035\ : Span4Mux_v
    port map (
            O => \N__6875\,
            I => \N__6863\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__6872\,
            I => \N__6863\
        );

    \I__1033\ : InMux
    port map (
            O => \N__6871\,
            I => \N__6860\
        );

    \I__1032\ : InMux
    port map (
            O => \N__6870\,
            I => \N__6857\
        );

    \I__1031\ : Odrv4
    port map (
            O => \N__6863\,
            I => \DUT.wRxByte_4\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__6860\,
            I => \DUT.wRxByte_4\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__6857\,
            I => \DUT.wRxByte_4\
        );

    \I__1028\ : InMux
    port map (
            O => \N__6850\,
            I => \N__6846\
        );

    \I__1027\ : InMux
    port map (
            O => \N__6849\,
            I => \N__6843\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__6846\,
            I => \N__6839\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__6843\,
            I => \N__6836\
        );

    \I__1024\ : InMux
    port map (
            O => \N__6842\,
            I => \N__6833\
        );

    \I__1023\ : Span4Mux_v
    port map (
            O => \N__6839\,
            I => \N__6824\
        );

    \I__1022\ : Span4Mux_v
    port map (
            O => \N__6836\,
            I => \N__6824\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__6833\,
            I => \N__6824\
        );

    \I__1020\ : InMux
    port map (
            O => \N__6832\,
            I => \N__6821\
        );

    \I__1019\ : InMux
    port map (
            O => \N__6831\,
            I => \N__6818\
        );

    \I__1018\ : Odrv4
    port map (
            O => \N__6824\,
            I => \DUT.wRxByte_5\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__6821\,
            I => \DUT.wRxByte_5\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__6818\,
            I => \DUT.wRxByte_5\
        );

    \I__1015\ : InMux
    port map (
            O => \N__6811\,
            I => \N__6807\
        );

    \I__1014\ : InMux
    port map (
            O => \N__6810\,
            I => \N__6804\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__6807\,
            I => \N__6800\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__6804\,
            I => \N__6797\
        );

    \I__1011\ : InMux
    port map (
            O => \N__6803\,
            I => \N__6794\
        );

    \I__1010\ : Span4Mux_v
    port map (
            O => \N__6800\,
            I => \N__6785\
        );

    \I__1009\ : Span4Mux_v
    port map (
            O => \N__6797\,
            I => \N__6785\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__6794\,
            I => \N__6785\
        );

    \I__1007\ : InMux
    port map (
            O => \N__6793\,
            I => \N__6782\
        );

    \I__1006\ : InMux
    port map (
            O => \N__6792\,
            I => \N__6779\
        );

    \I__1005\ : Odrv4
    port map (
            O => \N__6785\,
            I => \DUT.wRxByte_6\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__6782\,
            I => \DUT.wRxByte_6\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__6779\,
            I => \DUT.wRxByte_6\
        );

    \I__1002\ : InMux
    port map (
            O => \N__6772\,
            I => \N__6769\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__6769\,
            I => \N__6765\
        );

    \I__1000\ : InMux
    port map (
            O => \N__6768\,
            I => \N__6761\
        );

    \I__999\ : Span4Mux_h
    port map (
            O => \N__6765\,
            I => \N__6756\
        );

    \I__998\ : InMux
    port map (
            O => \N__6764\,
            I => \N__6753\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__6761\,
            I => \N__6750\
        );

    \I__996\ : InMux
    port map (
            O => \N__6760\,
            I => \N__6747\
        );

    \I__995\ : InMux
    port map (
            O => \N__6759\,
            I => \N__6744\
        );

    \I__994\ : Odrv4
    port map (
            O => \N__6756\,
            I => \DUT.wRxByte_7\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__6753\,
            I => \DUT.wRxByte_7\
        );

    \I__992\ : Odrv4
    port map (
            O => \N__6750\,
            I => \DUT.wRxByte_7\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__6747\,
            I => \DUT.wRxByte_7\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__6744\,
            I => \DUT.wRxByte_7\
        );

    \I__989\ : CascadeMux
    port map (
            O => \N__6733\,
            I => \G_141_cascade_\
        );

    \I__988\ : CascadeMux
    port map (
            O => \N__6730\,
            I => \N__6726\
        );

    \I__987\ : CascadeMux
    port map (
            O => \N__6729\,
            I => \N__6722\
        );

    \I__986\ : InMux
    port map (
            O => \N__6726\,
            I => \N__6715\
        );

    \I__985\ : InMux
    port map (
            O => \N__6725\,
            I => \N__6715\
        );

    \I__984\ : InMux
    port map (
            O => \N__6722\,
            I => \N__6708\
        );

    \I__983\ : InMux
    port map (
            O => \N__6721\,
            I => \N__6708\
        );

    \I__982\ : InMux
    port map (
            O => \N__6720\,
            I => \N__6708\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__6715\,
            I => \G_140\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__6708\,
            I => \G_140\
        );

    \I__979\ : InMux
    port map (
            O => \N__6703\,
            I => \N__6700\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__6700\,
            I => \fifo_inst_ftdi_input_inst_oTxFull_0\
        );

    \I__977\ : CascadeMux
    port map (
            O => \N__6697\,
            I => \G_140_cascade_\
        );

    \I__976\ : InMux
    port map (
            O => \N__6694\,
            I => \N__6684\
        );

    \I__975\ : InMux
    port map (
            O => \N__6693\,
            I => \N__6684\
        );

    \I__974\ : InMux
    port map (
            O => \N__6692\,
            I => \N__6684\
        );

    \I__973\ : InMux
    port map (
            O => \N__6691\,
            I => \N__6681\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__6684\,
            I => \G_143\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__6681\,
            I => \G_143\
        );

    \I__970\ : InMux
    port map (
            O => \N__6676\,
            I => \N__6667\
        );

    \I__969\ : InMux
    port map (
            O => \N__6675\,
            I => \N__6667\
        );

    \I__968\ : InMux
    port map (
            O => \N__6674\,
            I => \N__6667\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__6667\,
            I => \G_146\
        );

    \I__966\ : InMux
    port map (
            O => \N__6664\,
            I => \N__6661\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__6661\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_0\
        );

    \I__964\ : CascadeMux
    port map (
            O => \N__6658\,
            I => \N__6655\
        );

    \I__963\ : InMux
    port map (
            O => \N__6655\,
            I => \N__6652\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__6652\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_1\
        );

    \I__961\ : CascadeMux
    port map (
            O => \N__6649\,
            I => \N__6646\
        );

    \I__960\ : InMux
    port map (
            O => \N__6646\,
            I => \N__6643\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__6643\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_2\
        );

    \I__958\ : CascadeMux
    port map (
            O => \N__6640\,
            I => \N__6637\
        );

    \I__957\ : InMux
    port map (
            O => \N__6637\,
            I => \N__6634\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__6634\,
            I => \N__6631\
        );

    \I__955\ : Span4Mux_v
    port map (
            O => \N__6631\,
            I => \N__6628\
        );

    \I__954\ : Odrv4
    port map (
            O => \N__6628\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_3\
        );

    \I__953\ : CascadeMux
    port map (
            O => \N__6625\,
            I => \N__6622\
        );

    \I__952\ : InMux
    port map (
            O => \N__6622\,
            I => \N__6619\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__6619\,
            I => \N__6616\
        );

    \I__950\ : Span4Mux_h
    port map (
            O => \N__6616\,
            I => \N__6613\
        );

    \I__949\ : Odrv4
    port map (
            O => \N__6613\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_4\
        );

    \I__948\ : CascadeMux
    port map (
            O => \N__6610\,
            I => \N__6607\
        );

    \I__947\ : InMux
    port map (
            O => \N__6607\,
            I => \N__6604\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__6604\,
            I => \N__6601\
        );

    \I__945\ : Span4Mux_h
    port map (
            O => \N__6601\,
            I => \N__6598\
        );

    \I__944\ : Odrv4
    port map (
            O => \N__6598\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_5\
        );

    \I__943\ : CascadeMux
    port map (
            O => \N__6595\,
            I => \N__6592\
        );

    \I__942\ : InMux
    port map (
            O => \N__6592\,
            I => \N__6589\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__6589\,
            I => \N__6586\
        );

    \I__940\ : Span4Mux_h
    port map (
            O => \N__6586\,
            I => \N__6583\
        );

    \I__939\ : Odrv4
    port map (
            O => \N__6583\,
            I => \DUT.fifo_rx_inst.rFifoData_ram1_6\
        );

    \I__938\ : CEMux
    port map (
            O => \N__6580\,
            I => \N__6576\
        );

    \I__937\ : CEMux
    port map (
            O => \N__6579\,
            I => \N__6573\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__6576\,
            I => \DUT.fifo_tx_inst.N_40\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__6573\,
            I => \DUT.fifo_tx_inst.N_40\
        );

    \I__934\ : CascadeMux
    port map (
            O => \N__6568\,
            I => \G_145_cascade_\
        );

    \I__933\ : InMux
    port map (
            O => \N__6565\,
            I => \N__6559\
        );

    \I__932\ : InMux
    port map (
            O => \N__6564\,
            I => \N__6559\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__6559\,
            I => \G_145\
        );

    \I__930\ : CascadeMux
    port map (
            O => \N__6556\,
            I => \G_142_cascade_\
        );

    \I__929\ : InMux
    port map (
            O => \N__6553\,
            I => \N__6542\
        );

    \I__928\ : InMux
    port map (
            O => \N__6552\,
            I => \N__6542\
        );

    \I__927\ : InMux
    port map (
            O => \N__6551\,
            I => \N__6542\
        );

    \I__926\ : InMux
    port map (
            O => \N__6550\,
            I => \N__6539\
        );

    \I__925\ : InMux
    port map (
            O => \N__6549\,
            I => \N__6536\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__6542\,
            I => \G_144\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__6539\,
            I => \G_144\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__6536\,
            I => \G_144\
        );

    \I__921\ : InMux
    port map (
            O => \N__6529\,
            I => \N__6526\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__6526\,
            I => \fifo_inst.ftdi_input_inst.SUMZ0Z_3\
        );

    \I__919\ : SRMux
    port map (
            O => \N__6523\,
            I => \N__6520\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__6520\,
            I => \N__6517\
        );

    \I__917\ : Span4Mux_h
    port map (
            O => \N__6517\,
            I => \N__6512\
        );

    \I__916\ : InMux
    port map (
            O => \N__6516\,
            I => \N__6509\
        );

    \I__915\ : InMux
    port map (
            O => \N__6515\,
            I => \N__6506\
        );

    \I__914\ : Odrv4
    port map (
            O => \N__6512\,
            I => \G_147\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__6509\,
            I => \G_147\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__6506\,
            I => \G_147\
        );

    \I__911\ : CascadeMux
    port map (
            O => \N__6499\,
            I => \N__6493\
        );

    \I__910\ : InMux
    port map (
            O => \N__6498\,
            I => \N__6484\
        );

    \I__909\ : InMux
    port map (
            O => \N__6497\,
            I => \N__6484\
        );

    \I__908\ : InMux
    port map (
            O => \N__6496\,
            I => \N__6484\
        );

    \I__907\ : InMux
    port map (
            O => \N__6493\,
            I => \N__6484\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__6484\,
            I => \G_142\
        );

    \I__905\ : InMux
    port map (
            O => \N__6481\,
            I => \N__6474\
        );

    \I__904\ : InMux
    port map (
            O => \N__6480\,
            I => \N__6474\
        );

    \I__903\ : InMux
    port map (
            O => \N__6479\,
            I => \N__6471\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__6474\,
            I => \G_141\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__6471\,
            I => \G_141\
        );

    \I__900\ : InMux
    port map (
            O => \N__6466\,
            I => \N__6463\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__6463\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_5\
        );

    \I__898\ : CascadeMux
    port map (
            O => \N__6460\,
            I => \N__6457\
        );

    \I__897\ : InMux
    port map (
            O => \N__6457\,
            I => \N__6454\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__6454\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_5\
        );

    \I__895\ : CascadeMux
    port map (
            O => \N__6451\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_\
        );

    \I__894\ : InMux
    port map (
            O => \N__6448\,
            I => \N__6445\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__6445\,
            I => \N__6442\
        );

    \I__892\ : Odrv4
    port map (
            O => \N__6442\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_5\
        );

    \I__891\ : InMux
    port map (
            O => \N__6439\,
            I => \N__6436\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__6436\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_7\
        );

    \I__889\ : InMux
    port map (
            O => \N__6433\,
            I => \N__6430\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__6430\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_7\
        );

    \I__887\ : CascadeMux
    port map (
            O => \N__6427\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_\
        );

    \I__886\ : InMux
    port map (
            O => \N__6424\,
            I => \N__6421\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__6421\,
            I => \N__6418\
        );

    \I__884\ : Odrv4
    port map (
            O => \N__6418\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_7\
        );

    \I__883\ : InMux
    port map (
            O => \N__6415\,
            I => \N__6404\
        );

    \I__882\ : InMux
    port map (
            O => \N__6414\,
            I => \N__6401\
        );

    \I__881\ : InMux
    port map (
            O => \N__6413\,
            I => \N__6393\
        );

    \I__880\ : InMux
    port map (
            O => \N__6412\,
            I => \N__6393\
        );

    \I__879\ : InMux
    port map (
            O => \N__6411\,
            I => \N__6393\
        );

    \I__878\ : InMux
    port map (
            O => \N__6410\,
            I => \N__6389\
        );

    \I__877\ : InMux
    port map (
            O => \N__6409\,
            I => \N__6386\
        );

    \I__876\ : InMux
    port map (
            O => \N__6408\,
            I => \N__6381\
        );

    \I__875\ : InMux
    port map (
            O => \N__6407\,
            I => \N__6381\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__6404\,
            I => \N__6378\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__6401\,
            I => \N__6375\
        );

    \I__872\ : InMux
    port map (
            O => \N__6400\,
            I => \N__6372\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__6393\,
            I => \N__6369\
        );

    \I__870\ : InMux
    port map (
            O => \N__6392\,
            I => \N__6366\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__6389\,
            I => \DUT.fifo_tx_inst.N_33\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__6386\,
            I => \DUT.fifo_tx_inst.N_33\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__6381\,
            I => \DUT.fifo_tx_inst.N_33\
        );

    \I__866\ : Odrv4
    port map (
            O => \N__6378\,
            I => \DUT.fifo_tx_inst.N_33\
        );

    \I__865\ : Odrv12
    port map (
            O => \N__6375\,
            I => \DUT.fifo_tx_inst.N_33\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__6372\,
            I => \DUT.fifo_tx_inst.N_33\
        );

    \I__863\ : Odrv4
    port map (
            O => \N__6369\,
            I => \DUT.fifo_tx_inst.N_33\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__6366\,
            I => \DUT.fifo_tx_inst.N_33\
        );

    \I__861\ : CEMux
    port map (
            O => \N__6349\,
            I => \N__6346\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__6346\,
            I => \DUT.fifo_tx_inst.N_41\
        );

    \I__859\ : InMux
    port map (
            O => \N__6343\,
            I => \N__6340\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__6340\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_4\
        );

    \I__857\ : InMux
    port map (
            O => \N__6337\,
            I => \N__6334\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__6334\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_4\
        );

    \I__855\ : InMux
    port map (
            O => \N__6331\,
            I => \N__6328\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__6328\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_2\
        );

    \I__853\ : InMux
    port map (
            O => \N__6325\,
            I => \N__6322\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__6322\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_2\
        );

    \I__851\ : CascadeMux
    port map (
            O => \N__6319\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_\
        );

    \I__850\ : InMux
    port map (
            O => \N__6316\,
            I => \N__6313\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__6313\,
            I => \N__6310\
        );

    \I__848\ : Odrv4
    port map (
            O => \N__6310\,
            I => \DUT.fifo_tx_inst.rFifoData_ram2_2\
        );

    \I__847\ : CascadeMux
    port map (
            O => \N__6307\,
            I => \DUT.rFifoDatarx_2_cascade_\
        );

    \I__846\ : InMux
    port map (
            O => \N__6304\,
            I => \N__6300\
        );

    \I__845\ : InMux
    port map (
            O => \N__6303\,
            I => \N__6297\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__6300\,
            I => \DUT.fifo_tx_inst.rFifoDataro_1\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__6297\,
            I => \DUT.fifo_tx_inst.rFifoDataro_1\
        );

    \I__842\ : InMux
    port map (
            O => \N__6292\,
            I => \N__6288\
        );

    \I__841\ : InMux
    port map (
            O => \N__6291\,
            I => \N__6285\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__6288\,
            I => \DUT.fifo_tx_inst.rFifoDataro_0\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__6285\,
            I => \DUT.fifo_tx_inst.rFifoDataro_0\
        );

    \I__838\ : CascadeMux
    port map (
            O => \N__6280\,
            I => \DUT.fifo_tx_inst.rFifoDataror_1_0_cascade_\
        );

    \I__837\ : InMux
    port map (
            O => \N__6277\,
            I => \N__6274\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__6274\,
            I => \N__6271\
        );

    \I__835\ : Odrv4
    port map (
            O => \N__6271\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_0\
        );

    \I__834\ : InMux
    port map (
            O => \N__6268\,
            I => \N__6265\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__6265\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_0\
        );

    \I__832\ : CascadeMux
    port map (
            O => \N__6262\,
            I => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_\
        );

    \I__831\ : CascadeMux
    port map (
            O => \N__6259\,
            I => \DUT.fifo_tx_inst.un1_i11_2_i_cascade_\
        );

    \I__830\ : InMux
    port map (
            O => \N__6256\,
            I => \N__6253\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__6253\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_1\
        );

    \I__828\ : CascadeMux
    port map (
            O => \N__6250\,
            I => \N__6247\
        );

    \I__827\ : InMux
    port map (
            O => \N__6247\,
            I => \N__6244\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__6244\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_1\
        );

    \I__825\ : InMux
    port map (
            O => \N__6241\,
            I => \N__6238\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__6238\,
            I => \DUT.fifo_tx_inst.rFifoData_ram1_3\
        );

    \I__823\ : InMux
    port map (
            O => \N__6235\,
            I => \N__6232\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__6232\,
            I => \DUT.fifo_tx_inst.rFifoData_ram0_3\
        );

    \I__821\ : InMux
    port map (
            O => \N__6229\,
            I => \N__6226\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__6226\,
            I => \DUT.fifo_tx_inst.CO0\
        );

    \I__819\ : CascadeMux
    port map (
            O => \N__6223\,
            I => \DUT.fifo_tx_inst.CO0_cascade_\
        );

    \I__818\ : InMux
    port map (
            O => \N__6220\,
            I => \N__6217\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__6217\,
            I => \DUT.fifo_tx_inst.un1_i11_2_i\
        );

    \I__816\ : IoInMux
    port map (
            O => \N__6214\,
            I => \N__6211\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__6211\,
            I => \N__6208\
        );

    \I__814\ : Span4Mux_s1_v
    port map (
            O => \N__6208\,
            I => \N__6205\
        );

    \I__813\ : Span4Mux_v
    port map (
            O => \N__6205\,
            I => \N__6201\
        );

    \I__812\ : InMux
    port map (
            O => \N__6204\,
            I => \N__6198\
        );

    \I__811\ : Span4Mux_v
    port map (
            O => \N__6201\,
            I => \N__6193\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__6198\,
            I => \N__6193\
        );

    \I__809\ : Span4Mux_v
    port map (
            O => \N__6193\,
            I => \N__6189\
        );

    \I__808\ : InMux
    port map (
            O => \N__6192\,
            I => \N__6186\
        );

    \I__807\ : Odrv4
    port map (
            O => \N__6189\,
            I => \oTx_n_c\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__6186\,
            I => \oTx_n_c\
        );

    \I__805\ : IoInMux
    port map (
            O => \N__6181\,
            I => \N__6178\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__6178\,
            I => \N__6175\
        );

    \I__803\ : Span4Mux_s3_v
    port map (
            O => \N__6175\,
            I => \N__6172\
        );

    \I__802\ : Span4Mux_h
    port map (
            O => \N__6172\,
            I => \N__6169\
        );

    \I__801\ : Sp12to4
    port map (
            O => \N__6169\,
            I => \N__6166\
        );

    \I__800\ : Span12Mux_v
    port map (
            O => \N__6166\,
            I => \N__6162\
        );

    \I__799\ : InMux
    port map (
            O => \N__6165\,
            I => \N__6159\
        );

    \I__798\ : Odrv12
    port map (
            O => \N__6162\,
            I => \P1A2_c\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__6159\,
            I => \P1A2_c\
        );

    \I__796\ : InMux
    port map (
            O => \N__6154\,
            I => \N__6150\
        );

    \I__795\ : InMux
    port map (
            O => \N__6153\,
            I => \N__6147\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__6150\,
            I => \N__6139\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__6147\,
            I => \N__6139\
        );

    \I__792\ : InMux
    port map (
            O => \N__6146\,
            I => \N__6132\
        );

    \I__791\ : InMux
    port map (
            O => \N__6145\,
            I => \N__6132\
        );

    \I__790\ : InMux
    port map (
            O => \N__6144\,
            I => \N__6132\
        );

    \I__789\ : Odrv4
    port map (
            O => \N__6139\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_0\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__6132\,
            I => \DUT.fifo_tx_inst.rFifoCountZ0Z_0\
        );

    \I__787\ : CascadeMux
    port map (
            O => \N__6127\,
            I => \N__6124\
        );

    \I__786\ : InMux
    port map (
            O => \N__6124\,
            I => \N__6121\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__6121\,
            I => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0\
        );

    \I__784\ : InMux
    port map (
            O => \N__6118\,
            I => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0\
        );

    \I__783\ : CascadeMux
    port map (
            O => \N__6115\,
            I => \N__6111\
        );

    \I__782\ : CascadeMux
    port map (
            O => \N__6114\,
            I => \N__6108\
        );

    \I__781\ : InMux
    port map (
            O => \N__6111\,
            I => \N__6105\
        );

    \I__780\ : InMux
    port map (
            O => \N__6108\,
            I => \N__6102\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__6105\,
            I => \DUT.fifo_tx_inst.N_35\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__6102\,
            I => \DUT.fifo_tx_inst.N_35\
        );

    \I__777\ : InMux
    port map (
            O => \N__6097\,
            I => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1\
        );

    \I__776\ : InMux
    port map (
            O => \N__6094\,
            I => \N__6088\
        );

    \I__775\ : InMux
    port map (
            O => \N__6093\,
            I => \N__6088\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__6088\,
            I => \DUT.fifo_tx_inst.rFifoDataro_3\
        );

    \I__773\ : InMux
    port map (
            O => \N__6085\,
            I => \N__6079\
        );

    \I__772\ : InMux
    port map (
            O => \N__6084\,
            I => \N__6079\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__6079\,
            I => \DUT.fifo_tx_inst.rFifoDataro_2\
        );

    \I__770\ : InMux
    port map (
            O => \N__6076\,
            I => \N__6073\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__6073\,
            I => \DUT.fifo_rx_inst.rTxByte_42_0\
        );

    \I__768\ : CascadeMux
    port map (
            O => \N__6070\,
            I => \DUT.fifo_rx_inst.rTxByte_42_1_cascade_\
        );

    \I__767\ : InMux
    port map (
            O => \N__6067\,
            I => \N__6063\
        );

    \I__766\ : CascadeMux
    port map (
            O => \N__6066\,
            I => \N__6059\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__6063\,
            I => \N__6055\
        );

    \I__764\ : InMux
    port map (
            O => \N__6062\,
            I => \N__6050\
        );

    \I__763\ : InMux
    port map (
            O => \N__6059\,
            I => \N__6050\
        );

    \I__762\ : InMux
    port map (
            O => \N__6058\,
            I => \N__6047\
        );

    \I__761\ : Odrv4
    port map (
            O => \N__6055\,
            I => \wRxBufferEmpty_i_0\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__6050\,
            I => \wRxBufferEmpty_i_0\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__6047\,
            I => \wRxBufferEmpty_i_0\
        );

    \I__758\ : SRMux
    port map (
            O => \N__6040\,
            I => \N__6037\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__6037\,
            I => \N__6033\
        );

    \I__756\ : SRMux
    port map (
            O => \N__6036\,
            I => \N__6030\
        );

    \I__755\ : Span4Mux_v
    port map (
            O => \N__6033\,
            I => \N__6025\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__6030\,
            I => \N__6025\
        );

    \I__753\ : Sp12to4
    port map (
            O => \N__6025\,
            I => \N__6021\
        );

    \I__752\ : InMux
    port map (
            O => \N__6024\,
            I => \N__6018\
        );

    \I__751\ : Odrv12
    port map (
            O => \N__6021\,
            I => \rFifoDatarff_0_RNIHJV05\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__6018\,
            I => \rFifoDatarff_0_RNIHJV05\
        );

    \I__749\ : CascadeMux
    port map (
            O => \N__6013\,
            I => \N__6004\
        );

    \I__748\ : InMux
    port map (
            O => \N__6012\,
            I => \N__5976\
        );

    \I__747\ : InMux
    port map (
            O => \N__6011\,
            I => \N__5976\
        );

    \I__746\ : InMux
    port map (
            O => \N__6010\,
            I => \N__5976\
        );

    \I__745\ : InMux
    port map (
            O => \N__6009\,
            I => \N__5976\
        );

    \I__744\ : InMux
    port map (
            O => \N__6008\,
            I => \N__5976\
        );

    \I__743\ : InMux
    port map (
            O => \N__6007\,
            I => \N__5976\
        );

    \I__742\ : InMux
    port map (
            O => \N__6004\,
            I => \N__5976\
        );

    \I__741\ : InMux
    port map (
            O => \N__6003\,
            I => \N__5976\
        );

    \I__740\ : CascadeMux
    port map (
            O => \N__6002\,
            I => \N__5971\
        );

    \I__739\ : CascadeMux
    port map (
            O => \N__6001\,
            I => \N__5968\
        );

    \I__738\ : InMux
    port map (
            O => \N__6000\,
            I => \N__5951\
        );

    \I__737\ : InMux
    port map (
            O => \N__5999\,
            I => \N__5951\
        );

    \I__736\ : InMux
    port map (
            O => \N__5998\,
            I => \N__5951\
        );

    \I__735\ : InMux
    port map (
            O => \N__5997\,
            I => \N__5951\
        );

    \I__734\ : InMux
    port map (
            O => \N__5996\,
            I => \N__5951\
        );

    \I__733\ : InMux
    port map (
            O => \N__5995\,
            I => \N__5951\
        );

    \I__732\ : InMux
    port map (
            O => \N__5994\,
            I => \N__5951\
        );

    \I__731\ : InMux
    port map (
            O => \N__5993\,
            I => \N__5951\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__5976\,
            I => \N__5948\
        );

    \I__729\ : InMux
    port map (
            O => \N__5975\,
            I => \N__5941\
        );

    \I__728\ : InMux
    port map (
            O => \N__5974\,
            I => \N__5941\
        );

    \I__727\ : InMux
    port map (
            O => \N__5971\,
            I => \N__5941\
        );

    \I__726\ : InMux
    port map (
            O => \N__5968\,
            I => \N__5938\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__5951\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__724\ : Odrv4
    port map (
            O => \N__5948\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__5941\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__5938\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\
        );

    \I__721\ : InMux
    port map (
            O => \N__5929\,
            I => \N__5926\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__5926\,
            I => \DUT.fifo_rx_inst.rReadPtr_RNI4NC92Z0Z_0\
        );

    \I__719\ : CascadeMux
    port map (
            O => \N__5923\,
            I => \N__5920\
        );

    \I__718\ : InMux
    port map (
            O => \N__5920\,
            I => \N__5911\
        );

    \I__717\ : InMux
    port map (
            O => \N__5919\,
            I => \N__5911\
        );

    \I__716\ : InMux
    port map (
            O => \N__5918\,
            I => \N__5911\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__5911\,
            I => \DUT.fifo_rx_inst.N_73\
        );

    \I__714\ : CascadeMux
    port map (
            O => \N__5908\,
            I => \DUT.fifo_rx_inst.rReadPtr_RNI4NC92Z0Z_0_cascade_\
        );

    \I__713\ : InMux
    port map (
            O => \N__5905\,
            I => \N__5889\
        );

    \I__712\ : InMux
    port map (
            O => \N__5904\,
            I => \N__5889\
        );

    \I__711\ : InMux
    port map (
            O => \N__5903\,
            I => \N__5889\
        );

    \I__710\ : InMux
    port map (
            O => \N__5902\,
            I => \N__5889\
        );

    \I__709\ : InMux
    port map (
            O => \N__5901\,
            I => \N__5875\
        );

    \I__708\ : InMux
    port map (
            O => \N__5900\,
            I => \N__5875\
        );

    \I__707\ : InMux
    port map (
            O => \N__5899\,
            I => \N__5875\
        );

    \I__706\ : InMux
    port map (
            O => \N__5898\,
            I => \N__5875\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__5889\,
            I => \N__5872\
        );

    \I__704\ : InMux
    port map (
            O => \N__5888\,
            I => \N__5863\
        );

    \I__703\ : InMux
    port map (
            O => \N__5887\,
            I => \N__5863\
        );

    \I__702\ : InMux
    port map (
            O => \N__5886\,
            I => \N__5863\
        );

    \I__701\ : InMux
    port map (
            O => \N__5885\,
            I => \N__5863\
        );

    \I__700\ : InMux
    port map (
            O => \N__5884\,
            I => \N__5860\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__5875\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__698\ : Odrv4
    port map (
            O => \N__5872\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__5863\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__5860\,
            I => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\
        );

    \I__695\ : CascadeMux
    port map (
            O => \N__5851\,
            I => \DUT.uart_inst0.recv_state_srsts_1_0_6_cascade_\
        );

    \I__694\ : InMux
    port map (
            O => \N__5848\,
            I => \N__5844\
        );

    \I__693\ : InMux
    port map (
            O => \N__5847\,
            I => \N__5841\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__5844\,
            I => \DUT.fifo_rx_inst.un1_rFifoCount16_0_0\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__5841\,
            I => \DUT.fifo_rx_inst.un1_rFifoCount16_0_0\
        );

    \I__690\ : InMux
    port map (
            O => \N__5836\,
            I => \N__5833\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__5833\,
            I => \N__5828\
        );

    \I__688\ : CascadeMux
    port map (
            O => \N__5832\,
            I => \N__5825\
        );

    \I__687\ : InMux
    port map (
            O => \N__5831\,
            I => \N__5820\
        );

    \I__686\ : Span4Mux_h
    port map (
            O => \N__5828\,
            I => \N__5817\
        );

    \I__685\ : InMux
    port map (
            O => \N__5825\,
            I => \N__5814\
        );

    \I__684\ : InMux
    port map (
            O => \N__5824\,
            I => \N__5809\
        );

    \I__683\ : InMux
    port map (
            O => \N__5823\,
            I => \N__5809\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__5820\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_0\
        );

    \I__681\ : Odrv4
    port map (
            O => \N__5817\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_0\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__5814\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_0\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__5809\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_0\
        );

    \I__678\ : CEMux
    port map (
            O => \N__5800\,
            I => \N__5797\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__5797\,
            I => \N__5794\
        );

    \I__676\ : Sp12to4
    port map (
            O => \N__5794\,
            I => \N__5790\
        );

    \I__675\ : InMux
    port map (
            O => \N__5793\,
            I => \N__5787\
        );

    \I__674\ : Odrv12
    port map (
            O => \N__5790\,
            I => \DUT.fifo_rx_inst.rFifoData_awe0\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__5787\,
            I => \DUT.fifo_rx_inst.rFifoData_awe0\
        );

    \I__672\ : InMux
    port map (
            O => \N__5782\,
            I => \N__5778\
        );

    \I__671\ : InMux
    port map (
            O => \N__5781\,
            I => \N__5775\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__5778\,
            I => \DUT.fifo_rx_inst.rFifoDataro_0\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__5775\,
            I => \DUT.fifo_rx_inst.rFifoDataro_0\
        );

    \I__668\ : InMux
    port map (
            O => \N__5770\,
            I => \N__5767\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__5767\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_1\
        );

    \I__666\ : InMux
    port map (
            O => \N__5764\,
            I => \N__5761\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__5761\,
            I => \N__5758\
        );

    \I__664\ : Odrv4
    port map (
            O => \N__5758\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_1\
        );

    \I__663\ : CascadeMux
    port map (
            O => \N__5755\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1_cascade_\
        );

    \I__662\ : InMux
    port map (
            O => \N__5752\,
            I => \N__5749\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__5749\,
            I => \N__5746\
        );

    \I__660\ : Odrv4
    port map (
            O => \N__5746\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_1\
        );

    \I__659\ : InMux
    port map (
            O => \N__5743\,
            I => \N__5740\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__5740\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_7\
        );

    \I__657\ : InMux
    port map (
            O => \N__5737\,
            I => \N__5734\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__5734\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7\
        );

    \I__655\ : InMux
    port map (
            O => \N__5731\,
            I => \N__5728\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__5728\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_0\
        );

    \I__653\ : InMux
    port map (
            O => \N__5725\,
            I => \N__5722\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__5722\,
            I => \N__5719\
        );

    \I__651\ : Odrv4
    port map (
            O => \N__5719\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_0\
        );

    \I__650\ : InMux
    port map (
            O => \N__5716\,
            I => \N__5713\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__5713\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_0\
        );

    \I__648\ : CascadeMux
    port map (
            O => \N__5710\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_\
        );

    \I__647\ : CEMux
    port map (
            O => \N__5707\,
            I => \N__5703\
        );

    \I__646\ : CEMux
    port map (
            O => \N__5706\,
            I => \N__5700\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__5703\,
            I => \N__5697\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__5700\,
            I => \N__5694\
        );

    \I__643\ : Odrv4
    port map (
            O => \N__5697\,
            I => \wRxBufferEmpty_i_0_0\
        );

    \I__642\ : Odrv4
    port map (
            O => \N__5694\,
            I => \wRxBufferEmpty_i_0_0\
        );

    \I__641\ : InMux
    port map (
            O => \N__5689\,
            I => \N__5685\
        );

    \I__640\ : InMux
    port map (
            O => \N__5688\,
            I => \N__5682\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__5685\,
            I => \DUT.fifo_rx_inst.rFifoDataro_1\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__5682\,
            I => \DUT.fifo_rx_inst.rFifoDataro_1\
        );

    \I__637\ : CascadeMux
    port map (
            O => \N__5677\,
            I => \G_143_cascade_\
        );

    \I__636\ : CascadeMux
    port map (
            O => \N__5674\,
            I => \fifo_inst.ftdi_input_inst.SUMZ0Z_2_cascade_\
        );

    \I__635\ : CEMux
    port map (
            O => \N__5671\,
            I => \N__5667\
        );

    \I__634\ : CEMux
    port map (
            O => \N__5670\,
            I => \N__5664\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__5667\,
            I => \N__5660\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__5664\,
            I => \N__5657\
        );

    \I__631\ : CEMux
    port map (
            O => \N__5663\,
            I => \N__5654\
        );

    \I__630\ : Span4Mux_v
    port map (
            O => \N__5660\,
            I => \N__5651\
        );

    \I__629\ : Span4Mux_h
    port map (
            O => \N__5657\,
            I => \N__5647\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__5654\,
            I => \N__5642\
        );

    \I__627\ : Span4Mux_h
    port map (
            O => \N__5651\,
            I => \N__5642\
        );

    \I__626\ : InMux
    port map (
            O => \N__5650\,
            I => \N__5639\
        );

    \I__625\ : Odrv4
    port map (
            O => \N__5647\,
            I => \DUT.fifo_rx_inst.N_86\
        );

    \I__624\ : Odrv4
    port map (
            O => \N__5642\,
            I => \DUT.fifo_rx_inst.N_86\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__5639\,
            I => \DUT.fifo_rx_inst.N_86\
        );

    \I__622\ : InMux
    port map (
            O => \N__5632\,
            I => \N__5629\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__5629\,
            I => \N__5626\
        );

    \I__620\ : Odrv4
    port map (
            O => \N__5626\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_7\
        );

    \I__619\ : CascadeMux
    port map (
            O => \N__5623\,
            I => \N__5620\
        );

    \I__618\ : InMux
    port map (
            O => \N__5620\,
            I => \N__5617\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__5617\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_7\
        );

    \I__616\ : InMux
    port map (
            O => \N__5614\,
            I => \N__5611\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__5611\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_2\
        );

    \I__614\ : InMux
    port map (
            O => \N__5608\,
            I => \N__5605\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__5605\,
            I => \N__5602\
        );

    \I__612\ : Odrv12
    port map (
            O => \N__5602\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_2\
        );

    \I__611\ : CascadeMux
    port map (
            O => \N__5599\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2_cascade_\
        );

    \I__610\ : InMux
    port map (
            O => \N__5596\,
            I => \N__5593\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__5593\,
            I => \N__5590\
        );

    \I__608\ : Odrv4
    port map (
            O => \N__5590\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_2\
        );

    \I__607\ : CascadeMux
    port map (
            O => \N__5587\,
            I => \wRxBufferEmpty_i_0_cascade_\
        );

    \I__606\ : InMux
    port map (
            O => \N__5584\,
            I => \N__5581\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__5581\,
            I => \DUT.fifo_rx_inst.un1_rFifoCount16_0_i_0\
        );

    \I__604\ : CascadeMux
    port map (
            O => \N__5578\,
            I => \N__5575\
        );

    \I__603\ : InMux
    port map (
            O => \N__5575\,
            I => \N__5572\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__5572\,
            I => \DUT.fifo_rx_inst.rFifoCount_RNIK3G92Z0Z_1\
        );

    \I__601\ : InMux
    port map (
            O => \N__5569\,
            I => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0\
        );

    \I__600\ : InMux
    port map (
            O => \N__5566\,
            I => \N__5563\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__5563\,
            I => \DUT.fifo_rx_inst.un1_rFifoCount_1_axb_2\
        );

    \I__598\ : InMux
    port map (
            O => \N__5560\,
            I => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1\
        );

    \I__597\ : InMux
    port map (
            O => \N__5557\,
            I => \N__5552\
        );

    \I__596\ : InMux
    port map (
            O => \N__5556\,
            I => \N__5549\
        );

    \I__595\ : InMux
    port map (
            O => \N__5555\,
            I => \N__5542\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__5552\,
            I => \N__5537\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__5549\,
            I => \N__5537\
        );

    \I__592\ : InMux
    port map (
            O => \N__5548\,
            I => \N__5528\
        );

    \I__591\ : InMux
    port map (
            O => \N__5547\,
            I => \N__5528\
        );

    \I__590\ : InMux
    port map (
            O => \N__5546\,
            I => \N__5528\
        );

    \I__589\ : InMux
    port map (
            O => \N__5545\,
            I => \N__5528\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__5542\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\
        );

    \I__587\ : Odrv4
    port map (
            O => \N__5537\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__5528\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\
        );

    \I__585\ : CascadeMux
    port map (
            O => \N__5521\,
            I => \N__5515\
        );

    \I__584\ : InMux
    port map (
            O => \N__5520\,
            I => \N__5511\
        );

    \I__583\ : InMux
    port map (
            O => \N__5519\,
            I => \N__5508\
        );

    \I__582\ : InMux
    port map (
            O => \N__5518\,
            I => \N__5501\
        );

    \I__581\ : InMux
    port map (
            O => \N__5515\,
            I => \N__5501\
        );

    \I__580\ : InMux
    port map (
            O => \N__5514\,
            I => \N__5501\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__5511\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_1\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__5508\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_1\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__5501\,
            I => \DUT.fifo_rx_inst.rFifoCountZ0Z_1\
        );

    \I__576\ : CascadeMux
    port map (
            O => \N__5494\,
            I => \DUT.fifo_tx_inst.N_35_cascade_\
        );

    \I__575\ : InMux
    port map (
            O => \N__5491\,
            I => \N__5485\
        );

    \I__574\ : InMux
    port map (
            O => \N__5490\,
            I => \N__5485\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__5485\,
            I => \DUT.fifo_rx_inst.rFifoDataro_3\
        );

    \I__572\ : InMux
    port map (
            O => \N__5482\,
            I => \N__5476\
        );

    \I__571\ : InMux
    port map (
            O => \N__5481\,
            I => \N__5476\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__5476\,
            I => \DUT.fifo_rx_inst.rFifoDataro_2\
        );

    \I__569\ : InMux
    port map (
            O => \N__5473\,
            I => \N__5465\
        );

    \I__568\ : InMux
    port map (
            O => \N__5472\,
            I => \N__5465\
        );

    \I__567\ : InMux
    port map (
            O => \N__5471\,
            I => \N__5460\
        );

    \I__566\ : InMux
    port map (
            O => \N__5470\,
            I => \N__5460\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__5465\,
            I => \DUT.fifo_rx_inst.N_42\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__5460\,
            I => \DUT.fifo_rx_inst.N_42\
        );

    \I__563\ : CascadeMux
    port map (
            O => \N__5455\,
            I => \N__5447\
        );

    \I__562\ : InMux
    port map (
            O => \N__5454\,
            I => \N__5440\
        );

    \I__561\ : InMux
    port map (
            O => \N__5453\,
            I => \N__5440\
        );

    \I__560\ : InMux
    port map (
            O => \N__5452\,
            I => \N__5440\
        );

    \I__559\ : InMux
    port map (
            O => \N__5451\,
            I => \N__5433\
        );

    \I__558\ : InMux
    port map (
            O => \N__5450\,
            I => \N__5433\
        );

    \I__557\ : InMux
    port map (
            O => \N__5447\,
            I => \N__5433\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__5440\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_0\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__5433\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_0\
        );

    \I__554\ : CascadeMux
    port map (
            O => \N__5428\,
            I => \DUT.fifo_rx_inst.N_42_cascade_\
        );

    \I__553\ : CascadeMux
    port map (
            O => \N__5425\,
            I => \N__5419\
        );

    \I__552\ : InMux
    port map (
            O => \N__5424\,
            I => \N__5411\
        );

    \I__551\ : InMux
    port map (
            O => \N__5423\,
            I => \N__5411\
        );

    \I__550\ : InMux
    port map (
            O => \N__5422\,
            I => \N__5411\
        );

    \I__549\ : InMux
    port map (
            O => \N__5419\,
            I => \N__5406\
        );

    \I__548\ : InMux
    port map (
            O => \N__5418\,
            I => \N__5406\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__5411\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_1\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__5406\,
            I => \DUT.fifo_rx_inst.rWritePtrZ0Z_1\
        );

    \I__545\ : CascadeMux
    port map (
            O => \N__5401\,
            I => \DUT.fifo_rx_inst.rFifoData_awe1_cascade_\
        );

    \I__544\ : CascadeMux
    port map (
            O => \N__5398\,
            I => \N__5395\
        );

    \I__543\ : InMux
    port map (
            O => \N__5395\,
            I => \N__5392\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__5392\,
            I => \DUT.fifo_tx_inst.un1_i11_i\
        );

    \I__541\ : CascadeMux
    port map (
            O => \N__5389\,
            I => \DUT.fifo_tx_inst.un1_i11_i_cascade_\
        );

    \I__540\ : InMux
    port map (
            O => \N__5386\,
            I => \N__5383\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__5383\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_5\
        );

    \I__538\ : InMux
    port map (
            O => \N__5380\,
            I => \N__5377\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__5377\,
            I => \N__5374\
        );

    \I__536\ : Odrv4
    port map (
            O => \N__5374\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_6\
        );

    \I__535\ : InMux
    port map (
            O => \N__5371\,
            I => \N__5368\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__5368\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_6\
        );

    \I__533\ : CascadeMux
    port map (
            O => \N__5365\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6_cascade_\
        );

    \I__532\ : InMux
    port map (
            O => \N__5362\,
            I => \N__5359\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__5359\,
            I => \N__5356\
        );

    \I__530\ : Odrv4
    port map (
            O => \N__5356\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_6\
        );

    \I__529\ : InMux
    port map (
            O => \N__5353\,
            I => \N__5350\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__5350\,
            I => \N__5347\
        );

    \I__527\ : Odrv4
    port map (
            O => \N__5347\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_4\
        );

    \I__526\ : InMux
    port map (
            O => \N__5344\,
            I => \N__5341\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__5341\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4\
        );

    \I__524\ : InMux
    port map (
            O => \N__5338\,
            I => \N__5335\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__5335\,
            I => \N__5332\
        );

    \I__522\ : Odrv4
    port map (
            O => \N__5332\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_3\
        );

    \I__521\ : InMux
    port map (
            O => \N__5329\,
            I => \N__5326\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__5326\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_3\
        );

    \I__519\ : InMux
    port map (
            O => \N__5323\,
            I => \N__5320\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__5320\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_3\
        );

    \I__517\ : CascadeMux
    port map (
            O => \N__5317\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_\
        );

    \I__516\ : CEMux
    port map (
            O => \N__5314\,
            I => \N__5311\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__5311\,
            I => \N__5308\
        );

    \I__514\ : Span4Mux_v
    port map (
            O => \N__5308\,
            I => \N__5305\
        );

    \I__513\ : Odrv4
    port map (
            O => \N__5305\,
            I => \DUT.fifo_rx_inst.rFifoData_awe2\
        );

    \I__512\ : CascadeMux
    port map (
            O => \N__5302\,
            I => \DUT.fifo_rx_inst.rFifoData_awe2_cascade_\
        );

    \I__511\ : InMux
    port map (
            O => \N__5299\,
            I => \N__5296\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__5296\,
            I => \DUT.fifo_rx_inst.rFifoData_ram2_4\
        );

    \I__509\ : CascadeMux
    port map (
            O => \N__5293\,
            I => \N__5290\
        );

    \I__508\ : InMux
    port map (
            O => \N__5290\,
            I => \N__5287\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__5287\,
            I => \N__5284\
        );

    \I__506\ : Odrv4
    port map (
            O => \N__5284\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_4\
        );

    \I__505\ : InMux
    port map (
            O => \N__5281\,
            I => \N__5278\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__5278\,
            I => \N__5275\
        );

    \I__503\ : Odrv4
    port map (
            O => \N__5275\,
            I => \DUT.fifo_rx_inst.rFifoData_ram0_5\
        );

    \I__502\ : InMux
    port map (
            O => \N__5272\,
            I => \N__5269\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__5269\,
            I => \DUT.fifo_rx_inst.rFifoData_ram3_5\
        );

    \I__500\ : CascadeMux
    port map (
            O => \N__5266\,
            I => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_\
        );

    \I__499\ : CascadeMux
    port map (
            O => \N__5263\,
            I => \DUT.fifo_rx_inst.N_86_cascade_\
        );

    \I__498\ : InMux
    port map (
            O => \N__5260\,
            I => \N__5257\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__5257\,
            I => \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1\
        );

    \I__496\ : CascadeMux
    port map (
            O => \N__5254\,
            I => \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1_cascade_\
        );

    \I__495\ : IoInMux
    port map (
            O => \N__5251\,
            I => \N__5247\
        );

    \I__494\ : IoInMux
    port map (
            O => \N__5250\,
            I => \N__5244\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__5247\,
            I => \N__5239\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__5244\,
            I => \N__5236\
        );

    \I__491\ : IoInMux
    port map (
            O => \N__5243\,
            I => \N__5233\
        );

    \I__490\ : IoInMux
    port map (
            O => \N__5242\,
            I => \N__5230\
        );

    \I__489\ : IoSpan4Mux
    port map (
            O => \N__5239\,
            I => \N__5220\
        );

    \I__488\ : IoSpan4Mux
    port map (
            O => \N__5236\,
            I => \N__5220\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__5233\,
            I => \N__5220\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__5230\,
            I => \N__5220\
        );

    \I__485\ : IoInMux
    port map (
            O => \N__5229\,
            I => \N__5217\
        );

    \I__484\ : IoSpan4Mux
    port map (
            O => \N__5220\,
            I => \N__5209\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__5217\,
            I => \N__5209\
        );

    \I__482\ : IoInMux
    port map (
            O => \N__5216\,
            I => \N__5206\
        );

    \I__481\ : IoInMux
    port map (
            O => \N__5215\,
            I => \N__5203\
        );

    \I__480\ : IoInMux
    port map (
            O => \N__5214\,
            I => \N__5200\
        );

    \I__479\ : IoSpan4Mux
    port map (
            O => \N__5209\,
            I => \N__5197\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__5206\,
            I => \N__5194\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__5203\,
            I => \N__5189\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__5200\,
            I => \N__5189\
        );

    \I__475\ : Span4Mux_s2_v
    port map (
            O => \N__5197\,
            I => \N__5184\
        );

    \I__474\ : Span4Mux_s2_v
    port map (
            O => \N__5194\,
            I => \N__5184\
        );

    \I__473\ : IoSpan4Mux
    port map (
            O => \N__5189\,
            I => \N__5181\
        );

    \I__472\ : Span4Mux_v
    port map (
            O => \N__5184\,
            I => \N__5178\
        );

    \I__471\ : Sp12to4
    port map (
            O => \N__5181\,
            I => \N__5175\
        );

    \I__470\ : Span4Mux_v
    port map (
            O => \N__5178\,
            I => \N__5172\
        );

    \I__469\ : Span12Mux_v
    port map (
            O => \N__5175\,
            I => \N__5169\
        );

    \I__468\ : Span4Mux_v
    port map (
            O => \N__5172\,
            I => \N__5166\
        );

    \I__467\ : Odrv12
    port map (
            O => \N__5169\,
            I => \oTx_n_c_i\
        );

    \I__466\ : Odrv4
    port map (
            O => \N__5166\,
            I => \oTx_n_c_i\
        );

    \I__465\ : IoInMux
    port map (
            O => \N__5161\,
            I => \N__5158\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__5158\,
            I => \N__5155\
        );

    \I__463\ : Span4Mux_s3_v
    port map (
            O => \N__5155\,
            I => \N__5152\
        );

    \I__462\ : Span4Mux_v
    port map (
            O => \N__5152\,
            I => \N__5149\
        );

    \I__461\ : Span4Mux_h
    port map (
            O => \N__5149\,
            I => \N__5146\
        );

    \I__460\ : Odrv4
    port map (
            O => \N__5146\,
            I => \wRamRdData_1\
        );

    \I__459\ : InMux
    port map (
            O => \N__5143\,
            I => \N__5140\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__5140\,
            I => \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO\
        );

    \I__457\ : IoInMux
    port map (
            O => \N__5137\,
            I => \N__5134\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__5134\,
            I => \N__5131\
        );

    \I__455\ : Span12Mux_s9_v
    port map (
            O => \N__5131\,
            I => \N__5128\
        );

    \I__454\ : Span12Mux_v
    port map (
            O => \N__5128\,
            I => \N__5125\
        );

    \I__453\ : Odrv12
    port map (
            O => \N__5125\,
            I => \BTN_N_c\
        );

    \I__452\ : IoInMux
    port map (
            O => \N__5122\,
            I => \N__5119\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__5119\,
            I => \N__5116\
        );

    \I__450\ : Sp12to4
    port map (
            O => \N__5116\,
            I => \N__5113\
        );

    \I__449\ : Span12Mux_v
    port map (
            O => \N__5113\,
            I => \N__5110\
        );

    \I__448\ : Odrv12
    port map (
            O => \N__5110\,
            I => \wRamRdData_7\
        );

    \I__447\ : IoInMux
    port map (
            O => \N__5107\,
            I => \N__5104\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__5104\,
            I => \N__5101\
        );

    \I__445\ : Span4Mux_s1_v
    port map (
            O => \N__5101\,
            I => \N__5098\
        );

    \I__444\ : Span4Mux_v
    port map (
            O => \N__5098\,
            I => \N__5095\
        );

    \I__443\ : Span4Mux_v
    port map (
            O => \N__5095\,
            I => \N__5092\
        );

    \I__442\ : Span4Mux_h
    port map (
            O => \N__5092\,
            I => \N__5089\
        );

    \I__441\ : Odrv4
    port map (
            O => \N__5089\,
            I => \wRamRdData_0\
        );

    \I__440\ : IoInMux
    port map (
            O => \N__5086\,
            I => \N__5083\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__5083\,
            I => \N__5080\
        );

    \I__438\ : Span12Mux_s3_v
    port map (
            O => \N__5080\,
            I => \N__5077\
        );

    \I__437\ : Odrv12
    port map (
            O => \N__5077\,
            I => \wRamRdData_4\
        );

    \I__436\ : IoInMux
    port map (
            O => \N__5074\,
            I => \N__5071\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__5071\,
            I => \N__5068\
        );

    \I__434\ : Span12Mux_s10_v
    port map (
            O => \N__5068\,
            I => \N__5065\
        );

    \I__433\ : Odrv12
    port map (
            O => \N__5065\,
            I => \wRamRdData_6\
        );

    \I__432\ : IoInMux
    port map (
            O => \N__5062\,
            I => \N__5059\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__5059\,
            I => \N__5056\
        );

    \I__430\ : Span4Mux_s1_v
    port map (
            O => \N__5056\,
            I => \N__5053\
        );

    \I__429\ : Span4Mux_v
    port map (
            O => \N__5053\,
            I => \N__5050\
        );

    \I__428\ : Span4Mux_v
    port map (
            O => \N__5050\,
            I => \N__5047\
        );

    \I__427\ : Odrv4
    port map (
            O => \N__5047\,
            I => \wRamRdData_2\
        );

    \I__426\ : IoInMux
    port map (
            O => \N__5044\,
            I => \N__5041\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__5041\,
            I => \N__5038\
        );

    \I__424\ : Span4Mux_s1_v
    port map (
            O => \N__5038\,
            I => \N__5035\
        );

    \I__423\ : Span4Mux_v
    port map (
            O => \N__5035\,
            I => \N__5032\
        );

    \I__422\ : Span4Mux_v
    port map (
            O => \N__5032\,
            I => \N__5029\
        );

    \I__421\ : Odrv4
    port map (
            O => \N__5029\,
            I => \wRamRdData_3\
        );

    \I__420\ : IoInMux
    port map (
            O => \N__5026\,
            I => \N__5023\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__5023\,
            I => \N__5020\
        );

    \I__418\ : Span12Mux_s8_v
    port map (
            O => \N__5020\,
            I => \N__5017\
        );

    \I__417\ : Odrv12
    port map (
            O => \N__5017\,
            I => \wRamRdData_5\
        );

    \IN_MUX_bfv_18_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_19_0_\
        );

    \IN_MUX_bfv_18_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DUT.uart_inst0.tx_clk_divider_cry_7\,
            carryinitout => \bfn_18_20_0_\
        );

    \IN_MUX_bfv_16_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_16_0_\
        );

    \IN_MUX_bfv_18_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_13_0_\
        );

    \IN_MUX_bfv_18_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DUT.uart_inst0.rx_clk_divider_1_cry_7\,
            carryinitout => \bfn_18_14_0_\
        );

    \IN_MUX_bfv_18_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DUT.uart_inst0.rx_clk_divider_1_cry_15\,
            carryinitout => \bfn_18_15_0_\
        );

    \IN_MUX_bfv_14_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_19_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_18_0_\
        );

    \top_pll_inst.top_pll_inst_RNISDA2_1\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__10830\,
            GLOBALBUFFEROUTPUT => \wPllLocked_iso_i_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \top_pll_inst.top_pll_inst_RNISDA2\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__11536\,
            GLOBALBUFFEROUTPUT => \wPllLocked_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5143\,
            lcout => \wPllLocked\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6966\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12109\,
            ce => \N__5663\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6850\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12102\,
            ce => \N__5671\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6889\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12102\,
            ce => \N__5671\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6930\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12102\,
            ce => \N__5671\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6811\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12102\,
            ce => \N__5671\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_1_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010110100"
        )
    port map (
            in0 => \N__5473\,
            in1 => \N__5451\,
            in2 => \N__5425\,
            in3 => \N__5260\,
            lcout => \DUT.fifo_rx_inst.rWritePtrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI96D91_2_1_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__5557\,
            in1 => \N__5418\,
            in2 => \N__5455\,
            in3 => \N__7101\,
            lcout => \DUT.fifo_rx_inst.N_86\,
            ltout => \DUT.fifo_rx_inst.N_86_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1_1_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5263\,
            in3 => \N__11506\,
            lcout => \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1\,
            ltout => \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_0_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000101"
        )
    port map (
            in0 => \N__5450\,
            in1 => \_gnd_net_\,
            in2 => \N__5254\,
            in3 => \N__5472\,
            lcout => \DUT.fifo_rx_inst.rWritePtrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \oTx_n_c_sbtinv_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6204\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \oTx_n_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_0_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010000011011"
        )
    port map (
            in0 => \N__11619\,
            in1 => \N__6410\,
            in2 => \N__6115\,
            in3 => \N__6154\,
            lcout => \DUT.fifo_tx_inst.rFifoCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12080\,
            ce => 'H',
            sr => \N__12484\
        );

    \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__7528\,
            in1 => \N__7619\,
            in2 => \_gnd_net_\,
            in3 => \N__6400\,
            lcout => \DUT.fifo_tx_inst.N_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \top_pll_inst.top_pll_inst_RNISDA2_0_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11924\,
            lcout => \wPllLocked_iso_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7662\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12076\,
            ce => \N__10211\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7945\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12075\,
            ce => \N__10229\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7716\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12075\,
            ce => \N__10229\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7771\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12075\,
            ce => \N__10229\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7036\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12121\,
            ce => \N__5800\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7006\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12121\,
            ce => \N__5800\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6970\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12121\,
            ce => \N__5800\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6931\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12121\,
            ce => \N__5800\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6888\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12121\,
            ce => \N__5800\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6849\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12121\,
            ce => \N__5800\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6810\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12121\,
            ce => \N__5800\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6772\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12121\,
            ce => \N__5800\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7032\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12115\,
            ce => \N__5314\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7002\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12115\,
            ce => \N__5314\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6965\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12115\,
            ce => \N__5314\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6923\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12115\,
            ce => \N__5314\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6881\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12115\,
            ce => \N__5314\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6842\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12115\,
            ce => \N__5314\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6803\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12115\,
            ce => \N__5314\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6768\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12115\,
            ce => \N__5314\,
            sr => \_gnd_net_\
        );

    \rTxByte_esr_4_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110101"
        )
    port map (
            in0 => \N__5998\,
            in1 => \N__5299\,
            in2 => \N__5293\,
            in3 => \N__5344\,
            lcout => \rTxByteZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12110\,
            ce => \N__5706\,
            sr => \N__6040\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__5900\,
            in1 => \N__5281\,
            in2 => \N__6610\,
            in3 => \N__5995\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rTxByte_esr_5_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__5999\,
            in1 => \N__5272\,
            in2 => \N__5266\,
            in3 => \N__5386\,
            lcout => \rTxByteZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12110\,
            ce => \N__5706\,
            sr => \N__6040\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__5901\,
            in1 => \N__5380\,
            in2 => \N__6595\,
            in3 => \N__5996\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rTxByte_esr_6_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__6000\,
            in1 => \N__5371\,
            in2 => \N__5365\,
            in3 => \N__5362\,
            lcout => \rTxByteZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12110\,
            ce => \N__5706\,
            sr => \N__6040\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100011011"
        )
    port map (
            in0 => \N__5898\,
            in1 => \N__5353\,
            in2 => \N__6625\,
            in3 => \N__5993\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__5994\,
            in1 => \N__5338\,
            in2 => \N__6640\,
            in3 => \N__5899\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rTxByte_esr_3_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__5329\,
            in1 => \N__5323\,
            in2 => \N__5317\,
            in3 => \N__5997\,
            lcout => \rTxByteZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12110\,
            ce => \N__5706\,
            sr => \N__6040\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__5454\,
            in1 => \N__5424\,
            in2 => \_gnd_net_\,
            in3 => \N__5471\,
            lcout => \DUT.fifo_rx_inst.rFifoData_awe2\,
            ltout => \DUT.fifo_rx_inst.rFifoData_awe2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_2_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5302\,
            in3 => \N__5482\,
            lcout => \DUT.fifo_rx_inst.rFifoDataro_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12103\,
            ce => 'H',
            sr => \N__12491\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_3_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011101110"
        )
    port map (
            in0 => \N__5491\,
            in1 => \N__5650\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_rx_inst.rFifoDataro_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12103\,
            ce => 'H',
            sr => \N__12491\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111101111111"
        )
    port map (
            in0 => \N__5884\,
            in1 => \N__5490\,
            in2 => \N__6001\,
            in3 => \N__5481\,
            lcout => \DUT.fifo_rx_inst.rTxByte_42_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5452\,
            in1 => \N__5422\,
            in2 => \_gnd_net_\,
            in3 => \N__5470\,
            lcout => \DUT.fifo_rx_inst.rFifoData_awe0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7093\,
            in2 => \_gnd_net_\,
            in3 => \N__5556\,
            lcout => \DUT.fifo_rx_inst.N_42\,
            ltout => \DUT.fifo_rx_inst.N_42_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__5453\,
            in1 => \_gnd_net_\,
            in2 => \N__5428\,
            in3 => \N__5423\,
            lcout => \DUT.fifo_rx_inst.rFifoData_awe1\,
            ltout => \DUT.fifo_rx_inst.rFifoData_awe1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_1_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5401\,
            in3 => \N__5689\,
            lcout => \DUT.fifo_rx_inst.rFifoDataro_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12103\,
            ce => 'H',
            sr => \N__12491\
        );

    \DUT.fifo_tx_inst.rWritePtr_1_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100000100"
        )
    port map (
            in0 => \N__6413\,
            in1 => \N__7504\,
            in2 => \N__5398\,
            in3 => \N__7608\,
            lcout => \DUT.fifo_tx_inst.rWritePtrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12098\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_RNIJLJC_1_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110001111"
        )
    port map (
            in0 => \N__7502\,
            in1 => \N__7574\,
            in2 => \N__11520\,
            in3 => \N__6411\,
            lcout => \DUT.fifo_tx_inst.un1_i11_i\,
            ltout => \DUT.fifo_tx_inst.un1_i11_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_0_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000101"
        )
    port map (
            in0 => \N__6412\,
            in1 => \_gnd_net_\,
            in2 => \N__5389\,
            in3 => \N__7503\,
            lcout => \DUT.fifo_tx_inst.rWritePtrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12098\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNI9EGD1_0_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110111"
        )
    port map (
            in0 => \N__5824\,
            in1 => \N__8676\,
            in2 => \N__5521\,
            in3 => \N__5547\,
            lcout => \DUT.fifo_rx_inst.N_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNIK3G92_1_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__7092\,
            in1 => \N__5518\,
            in2 => \N__6066\,
            in3 => \N__8674\,
            lcout => \DUT.fifo_rx_inst.rFifoCount_RNIK3G92Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNO_0_2_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100011011001100"
        )
    port map (
            in0 => \N__8675\,
            in1 => \N__5548\,
            in2 => \N__7102\,
            in3 => \N__6062\,
            lcout => \DUT.fifo_rx_inst.un1_rFifoCount_1_axb_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__5545\,
            in1 => \N__5514\,
            in2 => \_gnd_net_\,
            in3 => \N__5823\,
            lcout => \wRxBufferEmpty_i_0\,
            ltout => \wRxBufferEmpty_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNIL4G92_2_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110011011"
        )
    port map (
            in0 => \N__8673\,
            in1 => \N__7091\,
            in2 => \N__5587\,
            in3 => \N__5546\,
            lcout => \DUT.fifo_rx_inst.un1_rFifoCount16_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_inv_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5584\,
            in2 => \N__5832\,
            in3 => \N__5847\,
            lcout => \DUT.fifo_rx_inst.un1_rFifoCount16_0_i_0\,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_1_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5519\,
            in2 => \N__5578\,
            in3 => \N__5569\,
            lcout => \DUT.fifo_rx_inst.rFifoCountZ0Z_1\,
            ltout => OPEN,
            carryin => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0\,
            carryout => \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1\,
            clk => \N__12091\,
            ce => 'H',
            sr => \N__12488\
        );

    \DUT.fifo_rx_inst.rFifoCount_2_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5566\,
            in2 => \_gnd_net_\,
            in3 => \N__5560\,
            lcout => \DUT.fifo_rx_inst.rFifoCountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12091\,
            ce => 'H',
            sr => \N__12488\
        );

    \rRxRead_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__5555\,
            in1 => \N__5520\,
            in2 => \_gnd_net_\,
            in3 => \N__5836\,
            lcout => \rRxReadZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12086\,
            ce => 'H',
            sr => \N__12486\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNIF689_0_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__7472\,
            in1 => \N__6145\,
            in2 => \N__8681\,
            in3 => \N__8621\,
            lcout => \DUT.fifo_tx_inst.N_35\,
            ltout => \DUT.fifo_tx_inst.N_35_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000111111"
        )
    port map (
            in0 => \N__6146\,
            in1 => \N__11617\,
            in2 => \N__5494\,
            in3 => \N__6392\,
            lcout => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNIMBD3_2_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__7471\,
            in1 => \_gnd_net_\,
            in2 => \N__8680\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_tx_inst.N_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNIN9O8_0_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__7470\,
            in1 => \N__6144\,
            in2 => \_gnd_net_\,
            in3 => \N__8620\,
            lcout => \DUT.N_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_1_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__7611\,
            in1 => \N__6304\,
            in2 => \N__7547\,
            in3 => \N__6408\,
            lcout => \DUT.fifo_tx_inst.rFifoDataro_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12081\,
            ce => 'H',
            sr => \N__12485\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_0_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001101"
        )
    port map (
            in0 => \N__7610\,
            in1 => \N__6292\,
            in2 => \N__7546\,
            in3 => \N__6407\,
            lcout => \DUT.fifo_tx_inst.rFifoDataro_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12081\,
            ce => 'H',
            sr => \N__12485\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8929\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12079\,
            ce => \N__6349\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8983\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12079\,
            ce => \N__6349\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7756\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12079\,
            ce => \N__6349\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_13_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10267\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12079\,
            ce => \N__6349\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7705\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12079\,
            ce => \N__6349\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7660\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12079\,
            ce => \N__6349\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8866\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12079\,
            ce => \N__6349\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7936\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12079\,
            ce => \N__6349\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7937\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12077\,
            ce => \N__6579\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7766\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12077\,
            ce => \N__6579\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10268\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12077\,
            ce => \N__6579\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8937\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12077\,
            ce => \N__6579\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7661\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12077\,
            ce => \N__6579\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8984\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12077\,
            ce => \N__6579\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7715\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12077\,
            ce => \N__6579\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_RNIN79A_0_1_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__7545\,
            in1 => \N__7609\,
            in2 => \_gnd_net_\,
            in3 => \N__6414\,
            lcout => \DUT.fifo_tx_inst.N_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.rPacketCount_latch_1_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010001000100"
        )
    port map (
            in0 => \N__12528\,
            in1 => \N__6691\,
            in2 => \N__6730\,
            in3 => \N__6480\,
            lcout => \G_143\,
            ltout => \G_143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.SUM_2_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6549\,
            in2 => \N__5677\,
            in3 => \N__6725\,
            lcout => OPEN,
            ltout => \fifo_inst.ftdi_input_inst.SUMZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.rPacketCount_latch_2_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__12529\,
            in1 => \N__6550\,
            in2 => \N__5674\,
            in3 => \N__6481\,
            lcout => \G_144\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7031\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12127\,
            ce => \N__5670\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7001\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12127\,
            ce => \N__5670\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6764\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12127\,
            ce => \N__5670\,
            sr => \_gnd_net_\
        );

    \rTxByte_esr_7_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011011101"
        )
    port map (
            in0 => \N__6012\,
            in1 => \N__5632\,
            in2 => \N__5623\,
            in3 => \N__5737\,
            lcout => \rTxByteZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12122\,
            ce => \N__5707\,
            sr => \N__6036\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__5614\,
            in1 => \N__6008\,
            in2 => \N__6649\,
            in3 => \N__5905\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rTxByte_esr_2_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__6011\,
            in1 => \N__5608\,
            in2 => \N__5599\,
            in3 => \N__5596\,
            lcout => \rTxByteZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12122\,
            ce => \N__5707\,
            sr => \N__6036\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__5770\,
            in1 => \N__6007\,
            in2 => \N__6658\,
            in3 => \N__5904\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rTxByte_esr_1_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__6010\,
            in1 => \N__5764\,
            in2 => \N__5755\,
            in3 => \N__5752\,
            lcout => \rTxByteZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12122\,
            ce => \N__5707\,
            sr => \N__6036\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__5743\,
            in1 => \N__6003\,
            in2 => \N__7060\,
            in3 => \N__5902\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__5903\,
            in1 => \N__6664\,
            in2 => \N__6013\,
            in3 => \N__5731\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rTxByte_esr_0_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__5725\,
            in1 => \N__5716\,
            in2 => \N__5710\,
            in3 => \N__6009\,
            lcout => \rTxByteZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12122\,
            ce => \N__5707\,
            sr => \N__6036\
        );

    \DUT.uart_inst0.rx_bits_remaining_3_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011101101"
        )
    port map (
            in0 => \N__7152\,
            in1 => \N__8157\,
            in2 => \N__7234\,
            in3 => \N__7194\,
            lcout => \DUT.uart_inst0.rx_bits_remainingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12116\,
            ce => \N__7213\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_0_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8156\,
            in2 => \_gnd_net_\,
            in3 => \N__7135\,
            lcout => \DUT.uart_inst0.rx_bits_remainingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12116\,
            ce => \N__7213\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_RNI250E6_0_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6067\,
            in2 => \_gnd_net_\,
            in3 => \N__6024\,
            lcout => \wRxBufferEmpty_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_0_RNI0AQO1_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110011"
        )
    port map (
            in0 => \N__5688\,
            in1 => \N__5781\,
            in2 => \N__6002\,
            in3 => \N__5885\,
            lcout => OPEN,
            ltout => \DUT.fifo_rx_inst.rTxByte_42_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_0_RNIHJV05_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010101010101"
        )
    port map (
            in0 => \N__11502\,
            in1 => \N__6076\,
            in2 => \N__6070\,
            in3 => \N__6058\,
            lcout => \rFifoDatarff_0_RNIHJV05\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rReadPtr_1_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000100100010"
        )
    port map (
            in0 => \N__5975\,
            in1 => \N__5929\,
            in2 => \N__5923\,
            in3 => \N__5888\,
            lcout => \DUT.fifo_rx_inst.rReadPtrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12111\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rReadPtr_RNI4NC92_0_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100001111"
        )
    port map (
            in0 => \N__5886\,
            in1 => \N__5918\,
            in2 => \N__11524\,
            in3 => \N__5974\,
            lcout => \DUT.fifo_rx_inst.rReadPtr_RNI4NC92Z0Z_0\,
            ltout => \DUT.fifo_rx_inst.rReadPtr_RNI4NC92Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rReadPtr_0_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000101"
        )
    port map (
            in0 => \N__5919\,
            in1 => \_gnd_net_\,
            in2 => \N__5908\,
            in3 => \N__5887\,
            lcout => \DUT.fifo_rx_inst.rReadPtrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12111\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_6_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__8238\,
            in1 => \N__11922\,
            in2 => \_gnd_net_\,
            in3 => \N__8261\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.recv_state_srsts_1_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_6_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8014\,
            in1 => \N__8431\,
            in2 => \N__5851\,
            in3 => \N__8366\,
            lcout => \DUT.wRcvd\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12111\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoCount_0_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5831\,
            in2 => \_gnd_net_\,
            in3 => \N__5848\,
            lcout => \DUT.fifo_rx_inst.rFifoCountZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12104\,
            ce => 'H',
            sr => \N__12492\
        );

    \DUT.fifo_rx_inst.rFifoDatarff_0_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5793\,
            in2 => \_gnd_net_\,
            in3 => \N__5782\,
            lcout => \DUT.fifo_rx_inst.rFifoDataro_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12104\,
            ce => 'H',
            sr => \N__12492\
        );

    \fifo_inst.ftdi_output_inst.oTx_n_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6192\,
            in2 => \_gnd_net_\,
            in3 => \N__9250\,
            lcout => \oTx_n_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12104\,
            ce => 'H',
            sr => \N__12492\
        );

    \fifo_inst.ftdi_output_inst.rWrDelay_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11044\,
            in2 => \_gnd_net_\,
            in3 => \N__11005\,
            lcout => \fifo_inst.ftdi_output_inst.rWrDelayZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12104\,
            ce => 'H',
            sr => \N__12492\
        );

    \fifo_inst.ftdi_output_inst.oRxFlag_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__6165\,
            in1 => \N__11296\,
            in2 => \_gnd_net_\,
            in3 => \N__9235\,
            lcout => \P1A2_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12099\,
            ce => 'H',
            sr => \N__12490\
        );

    \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6153\,
            in2 => \N__6127\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_19_0_\,
            carryout => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_1_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8622\,
            in2 => \N__8602\,
            in3 => \N__6118\,
            lcout => \DUT.fifo_tx_inst.rFifoCountZ0Z_1\,
            ltout => OPEN,
            carryin => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0\,
            carryout => \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1\,
            clk => \N__12092\,
            ce => 'H',
            sr => \N__12489\
        );

    \DUT.fifo_tx_inst.rFifoCount_2_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011100111000110"
        )
    port map (
            in0 => \N__11618\,
            in1 => \N__7474\,
            in2 => \N__6114\,
            in3 => \N__6097\,
            lcout => \DUT.fifo_tx_inst.rFifoCountZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12092\,
            ce => 'H',
            sr => \N__12489\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_3_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7896\,
            in2 => \_gnd_net_\,
            in3 => \N__6094\,
            lcout => \DUT.fifo_tx_inst.rFifoDataro_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12087\,
            ce => 'H',
            sr => \N__12487\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_2_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010111010"
        )
    port map (
            in0 => \N__6085\,
            in1 => \N__7541\,
            in2 => \N__7621\,
            in3 => \N__6409\,
            lcout => \DUT.fifo_tx_inst.rFifoDataro_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12087\,
            ce => 'H',
            sr => \N__12487\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010101110101"
        )
    port map (
            in0 => \N__7384\,
            in1 => \N__6093\,
            in2 => \N__9670\,
            in3 => \N__6084\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoDataror_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoDatarff_0_RNIJBAM_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110101"
        )
    port map (
            in0 => \N__6303\,
            in1 => \N__6291\,
            in2 => \N__6280\,
            in3 => \N__9642\,
            lcout => \DUT.rFifoDataror_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__7385\,
            in1 => \N__6277\,
            in2 => \N__9671\,
            in3 => \N__6268\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__7780\,
            in1 => \N__8890\,
            in2 => \N__6262\,
            in3 => \N__9643\,
            lcout => \DUT.rFifoDatarxZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rReadPtr_RNILV421_1_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__11501\,
            in1 => \N__9650\,
            in2 => \_gnd_net_\,
            in3 => \N__6229\,
            lcout => \DUT.fifo_tx_inst.un1_i11_2_i\,
            ltout => \DUT.fifo_tx_inst.un1_i11_2_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rReadPtr_0_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100000100"
        )
    port map (
            in0 => \N__8576\,
            in1 => \N__11621\,
            in2 => \N__6259\,
            in3 => \N__7392\,
            lcout => \DUT.fifo_tx_inst.rReadPtrZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12082\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__6256\,
            in1 => \N__9647\,
            in2 => \N__6250\,
            in3 => \N__7382\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__7380\,
            in1 => \N__6241\,
            in2 => \N__9672\,
            in3 => \N__6235\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rReadPtr_RNINFEP_0_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__11620\,
            in1 => \N__7383\,
            in2 => \_gnd_net_\,
            in3 => \N__8575\,
            lcout => \DUT.fifo_tx_inst.CO0\,
            ltout => \DUT.fifo_tx_inst.CO0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rReadPtr_1_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__9651\,
            in1 => \_gnd_net_\,
            in2 => \N__6223\,
            in3 => \N__6220\,
            lcout => \DUT.fifo_tx_inst.rReadPtrZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12082\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111011101"
        )
    port map (
            in0 => \N__6466\,
            in1 => \N__9648\,
            in2 => \N__6460\,
            in3 => \N__7381\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__9649\,
            in1 => \N__7633\,
            in2 => \N__6451\,
            in3 => \N__6448\,
            lcout => \DUT.rFifoDatarx_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110000011111"
        )
    port map (
            in0 => \N__6439\,
            in1 => \N__9652\,
            in2 => \N__7393\,
            in3 => \N__6433\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_14_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__9656\,
            in1 => \N__7909\,
            in2 => \N__6427\,
            in3 => \N__6424\,
            lcout => \DUT.rFifoDatarx_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_1_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__7548\,
            in1 => \N__7620\,
            in2 => \_gnd_net_\,
            in3 => \N__6415\,
            lcout => \DUT.fifo_tx_inst.N_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010000110111"
        )
    port map (
            in0 => \N__6343\,
            in1 => \N__7386\,
            in2 => \N__9673\,
            in3 => \N__6337\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001001010111"
        )
    port map (
            in0 => \N__7390\,
            in1 => \N__6331\,
            in2 => \N__9674\,
            in3 => \N__6325\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__9657\,
            in1 => \N__7726\,
            in2 => \N__6319\,
            in3 => \N__6316\,
            lcout => OPEN,
            ltout => \DUT.rFifoDatarx_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_RNO_0_2_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111000"
        )
    port map (
            in0 => \N__9910\,
            in1 => \N__12674\,
            in2 => \N__6307\,
            in3 => \N__10041\,
            lcout => \DUT.uart_inst0.tx_data_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8878\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12078\,
            ce => \N__6580\,
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.rWrState_latch_1_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \N__11918\,
            in1 => \N__6675\,
            in2 => \_gnd_net_\,
            in3 => \N__6564\,
            lcout => \G_145\,
            ltout => \G_145_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.rRamWrEn_latch_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001010"
        )
    port map (
            in0 => \N__6674\,
            in1 => \N__6515\,
            in2 => \N__6568\,
            in3 => \N__12534\,
            lcout => \G_147\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.un1_rWrState_1_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6676\,
            in2 => \_gnd_net_\,
            in3 => \N__6565\,
            lcout => \fifo_inst.ftdi_input_inst.un1_rWrStateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.un2_oPacketAvail_i_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6553\,
            in1 => \N__6498\,
            in2 => \N__6729\,
            in3 => \N__6694\,
            lcout => \fifo_inst.ftdi_input_inst.un2_oPacketAvail_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.rPacketCount_latch_3_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__6497\,
            in1 => \N__6479\,
            in2 => \N__12540\,
            in3 => \N__6529\,
            lcout => \G_142\,
            ltout => \G_142_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.oTxFull_0_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__6552\,
            in1 => \_gnd_net_\,
            in2 => \N__6556\,
            in3 => \_gnd_net_\,
            lcout => \fifo_inst_ftdi_input_inst_oTxFull_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.SUM_3_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__6693\,
            in1 => \N__6551\,
            in2 => \N__6499\,
            in3 => \N__6720\,
            lcout => \fifo_inst.ftdi_input_inst.SUMZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.rPacketCount15_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__6516\,
            in1 => \N__6496\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \G_141\,
            ltout => \G_141_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.rPacketCount_latch_0_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__12530\,
            in1 => \_gnd_net_\,
            in2 => \N__6733\,
            in3 => \N__6721\,
            lcout => \G_140\,
            ltout => \G_140_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.wTxEn_1_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000100"
        )
    port map (
            in0 => \N__6703\,
            in1 => \N__11919\,
            in2 => \N__6697\,
            in3 => \N__6692\,
            lcout => \G_146\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7024\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12132\,
            ce => \N__7051\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6994\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12132\,
            ce => \N__7051\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6955\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12132\,
            ce => \N__7051\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6913\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12132\,
            ce => \N__7051\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6871\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12132\,
            ce => \N__7051\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6832\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12132\,
            ce => \N__7051\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6793\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12132\,
            ce => \N__7051\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6760\,
            lcout => \DUT.fifo_rx_inst.rFifoData_ram1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12132\,
            ce => \N__7051\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_0_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6993\,
            lcout => \DUT.wRxByte_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12128\,
            ce => \N__7114\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_1_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6954\,
            lcout => \DUT.wRxByte_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12128\,
            ce => \N__7114\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_2_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6912\,
            lcout => \DUT.wRxByte_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12128\,
            ce => \N__7114\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_3_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6870\,
            lcout => \DUT.wRxByte_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12128\,
            ce => \N__7114\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_4_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6831\,
            lcout => \DUT.wRxByte_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12128\,
            ce => \N__7114\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_5_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6792\,
            lcout => \DUT.wRxByte_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12128\,
            ce => \N__7114\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_6_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6759\,
            lcout => \DUT.wRxByte_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12128\,
            ce => \N__7114\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_data_7_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8223\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DUT.wRxByte_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12128\,
            ce => \N__7114\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNIQJ1OI_2_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__7312\,
            in1 => \N__8418\,
            in2 => \N__8367\,
            in3 => \N__8010\,
            lcout => \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNITG1J4_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001101010101010"
        )
    port map (
            in0 => \N__8314\,
            in1 => \N__8089\,
            in2 => \N__8059\,
            in3 => \N__9196\,
            lcout => \DUT.uart_inst0.rx_countdown_3_2\,
            ltout => \DUT.uart_inst0.rx_countdown_3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011010000"
        )
    port map (
            in0 => \N__8041\,
            in1 => \N__8228\,
            in2 => \N__7105\,
            in3 => \N__8289\,
            lcout => \DUT.uart_inst0.rx_countdown_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_0_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101010"
        )
    port map (
            in0 => \N__11921\,
            in1 => \N__8039\,
            in2 => \N__8239\,
            in3 => \N__7100\,
            lcout => \DUT.uart_inst0.recv_state_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNIT7PG_1_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__7138\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7177\,
            lcout => \DUT.uart_inst0.N_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_5_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8116\,
            in1 => \N__8011\,
            in2 => \N__8368\,
            in3 => \N__8419\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNIHH651_0_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__8290\,
            in1 => \N__8224\,
            in2 => \_gnd_net_\,
            in3 => \N__8040\,
            lcout => \DUT.uart_inst0.N_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNIEMU42_5_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000111001101"
        )
    port map (
            in0 => \N__8540\,
            in1 => \N__9069\,
            in2 => \N__9169\,
            in3 => \N__9180\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.rx_countdown_8_i_o2_2_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNIDB3D7_0_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111110101111"
        )
    port map (
            in0 => \N__9070\,
            in1 => \N__8103\,
            in2 => \N__7063\,
            in3 => \N__9127\,
            lcout => \DUT.uart_inst0.rx_countdown_8_i_o2_2_2\,
            ltout => \DUT.uart_inst0.rx_countdown_8_i_o2_2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNIIQN8I_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000001"
        )
    port map (
            in0 => \N__8416\,
            in1 => \N__8008\,
            in2 => \N__7243\,
            in3 => \_gnd_net_\,
            lcout => \DUT.uart_inst0.recv_N_5_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_1_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__8009\,
            in1 => \N__8417\,
            in2 => \N__8369\,
            in3 => \N__11194\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.recv_state_RNO_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_1_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000000100"
        )
    port map (
            in0 => \N__11195\,
            in1 => \N__11527\,
            in2 => \N__7240\,
            in3 => \N__8158\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNIBTG71_2_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000000"
        )
    port map (
            in0 => \N__8229\,
            in1 => \N__8150\,
            in2 => \N__11535\,
            in3 => \N__7290\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.un1_m2_e_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNITN8GJ_2_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__8415\,
            in1 => \N__8007\,
            in2 => \N__7237\,
            in3 => \N__8355\,
            lcout => \DUT.uart_inst0.recv_state_RNITN8GJZ0Z_2\,
            ltout => \DUT.uart_inst0.recv_state_RNITN8GJZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_2_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100010000"
        )
    port map (
            in0 => \N__7233\,
            in1 => \N__8151\,
            in2 => \N__7216\,
            in3 => \N__7195\,
            lcout => \DUT.uart_inst0.rx_bits_remainingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12117\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010101"
        )
    port map (
            in0 => \N__7292\,
            in1 => \N__8242\,
            in2 => \_gnd_net_\,
            in3 => \N__8152\,
            lcout => \DUT.uart_inst0.rx_countdown_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNI8P9F_2_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11925\,
            in2 => \_gnd_net_\,
            in3 => \N__7291\,
            lcout => \DUT.uart_inst0.rx_m2_e_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_1_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000111110000"
        )
    port map (
            in0 => \N__7137\,
            in1 => \N__8154\,
            in2 => \N__7176\,
            in3 => \N__7206\,
            lcout => \DUT.uart_inst0.rx_bits_remainingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_bits_remaining_RNIUJI11_3_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__7193\,
            in1 => \N__7169\,
            in2 => \N__7156\,
            in3 => \N__7136\,
            lcout => \DUT.uart_inst0.N_98_4\,
            ltout => \DUT.uart_inst0.N_98_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_2_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011110101"
        )
    port map (
            in0 => \N__7294\,
            in1 => \N__8241\,
            in2 => \N__7315\,
            in3 => \N__8153\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.r_N_5_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_2_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__11525\,
            in1 => \N__7311\,
            in2 => \N__7297\,
            in3 => \N__7263\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_3_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7293\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7273\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.r_N_3_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_3_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__11526\,
            in1 => \N__8262\,
            in2 => \N__7267\,
            in3 => \N__7264\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12112\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_0_4_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__9405\,
            in1 => \N__9513\,
            in2 => \N__7252\,
            in3 => \N__11396\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_4_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100100001011010"
        )
    port map (
            in0 => \N__9335\,
            in1 => \N__12323\,
            in2 => \N__7255\,
            in3 => \N__9986\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12105\,
            ce => \N__11844\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNO_4_2_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__9402\,
            in1 => \N__9333\,
            in2 => \_gnd_net_\,
            in3 => \N__9832\,
            lcout => \DUT.uart_inst0.un1_tx_bits_remaining_axbxc2_N_4L5_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_1_4_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000101"
        )
    port map (
            in0 => \N__9754\,
            in1 => \_gnd_net_\,
            in2 => \N__9850\,
            in3 => \_gnd_net_\,
            lcout => \DUT.uart_inst0.g3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_RNO_4_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9403\,
            in1 => \N__9334\,
            in2 => \N__9463\,
            in3 => \N__9509\,
            lcout => \DUT.uart_inst0.g0_i_a4_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_3_3_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9837\,
            in1 => \N__12322\,
            in2 => \N__9521\,
            in3 => \N__9461\,
            lcout => \DUT.uart_inst0.un1_m7_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_2_3_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__9404\,
            in1 => \N__9833\,
            in2 => \_gnd_net_\,
            in3 => \N__9753\,
            lcout => \DUT.uart_inst0.tx_countdown_0_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNIUUGK1_3_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9385\,
            in1 => \N__9831\,
            in2 => \N__9517\,
            in3 => \N__9740\,
            lcout => \DUT.uart_inst0.tx_countdown_0_c4_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011011101"
        )
    port map (
            in0 => \N__11392\,
            in1 => \N__7342\,
            in2 => \_gnd_net_\,
            in3 => \N__9503\,
            lcout => \DUT.uart_inst0.tx_countdown_7_1_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_4_3_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000010000"
        )
    port map (
            in0 => \N__9386\,
            in1 => \N__9741\,
            in2 => \N__12673\,
            in3 => \N__11393\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.un1_tx_state_0_a4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110011101100"
        )
    port map (
            in0 => \N__7336\,
            in1 => \N__10288\,
            in2 => \N__7330\,
            in3 => \N__9343\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.un1_tx_clk_divider_s1_sn_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_3_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000011011101"
        )
    port map (
            in0 => \N__9966\,
            in1 => \N__12339\,
            in2 => \N__7327\,
            in3 => \N__7324\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12100\,
            ce => \N__11848\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_0_1_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011110101"
        )
    port map (
            in0 => \N__11394\,
            in1 => \_gnd_net_\,
            in2 => \N__9764\,
            in3 => \N__9849\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_countdown_RNO_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_1_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100000101"
        )
    port map (
            in0 => \N__9965\,
            in1 => \_gnd_net_\,
            in2 => \N__7318\,
            in3 => \N__12338\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12100\,
            ce => \N__11848\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_0_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100100001011010"
        )
    port map (
            in0 => \N__11395\,
            in1 => \N__12340\,
            in2 => \N__9765\,
            in3 => \N__9964\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12100\,
            ce => \N__11848\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_4_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__10896\,
            in1 => \N__7423\,
            in2 => \N__10075\,
            in3 => \N__9989\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_RNO_6_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__9347\,
            in1 => \N__9505\,
            in2 => \N__9457\,
            in3 => \N__9399\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g0_i_o4_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_RNO_3_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__12317\,
            in1 => \N__12662\,
            in2 => \N__7624\,
            in3 => \N__9842\,
            lcout => \DUT.uart_inst0.g0_i_o4_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNIN79A_2_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__7612\,
            in1 => \N__8683\,
            in2 => \N__7549\,
            in3 => \N__7473\,
            lcout => \DUT.fifo_tx_inst.rFifoData_awe3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_RNO_0_0_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111000000"
        )
    port map (
            in0 => \N__10026\,
            in1 => \N__8718\,
            in2 => \N__12675\,
            in3 => \N__7450\,
            lcout => \DUT.uart_inst0.tx_data_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__7444\,
            in1 => \N__9660\,
            in2 => \N__7675\,
            in3 => \N__7432\,
            lcout => OPEN,
            ltout => \DUT.rFifoDatarx_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_RNO_0_4_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__12666\,
            in1 => \N__9007\,
            in2 => \N__7426\,
            in3 => \N__10030\,
            lcout => \DUT.uart_inst0.tx_data_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110101111"
        )
    port map (
            in0 => \N__9658\,
            in1 => \N__7417\,
            in2 => \N__7405\,
            in3 => \N__7391\,
            lcout => OPEN,
            ltout => \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__7954\,
            in1 => \N__8836\,
            in2 => \N__7789\,
            in3 => \N__9659\,
            lcout => \DUT.rFifoDatarx_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_2_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__7786\,
            in1 => \N__10904\,
            in2 => \N__8746\,
            in3 => \N__9993\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12088\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_0_2_LC_15_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__9855\,
            in1 => \N__9771\,
            in2 => \_gnd_net_\,
            in3 => \N__11398\,
            lcout => \DUT.uart_inst0.N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8933\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12083\,
            ce => \N__7903\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8991\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12083\,
            ce => \N__7903\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7767\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12083\,
            ce => \N__7903\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_15_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10275\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12083\,
            ce => \N__7903\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7717\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12083\,
            ce => \N__7903\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7666\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12083\,
            ce => \N__7903\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8876\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12083\,
            ce => \N__7903\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7944\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12083\,
            ce => \N__7903\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_RNO_0_7_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12672\,
            in2 => \_gnd_net_\,
            in3 => \N__7885\,
            lcout => \DUT.uart_inst0.tx_data_8_321_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.SUM_0_2_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__7847\,
            in1 => \N__7868\,
            in2 => \_gnd_net_\,
            in3 => \N__7810\,
            lcout => OPEN,
            ltout => \G_152_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_2_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011100010"
        )
    port map (
            in0 => \N__7869\,
            in1 => \N__7834\,
            in2 => \N__7879\,
            in3 => \N__12539\,
            lcout => \G_151\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_1_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000001010"
        )
    port map (
            in0 => \N__7848\,
            in1 => \N__7812\,
            in2 => \N__12541\,
            in3 => \N__7833\,
            lcout => \G_150\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_0_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__12535\,
            in1 => \N__7811\,
            in2 => \_gnd_net_\,
            in3 => \N__7832\,
            lcout => \G_149\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_input_inst.oPacketAvail_latch_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__11920\,
            in1 => \N__9264\,
            in2 => \_gnd_net_\,
            in3 => \N__7795\,
            lcout => \G_148\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNI237O_0_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__8183\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8038\,
            lcout => \DUT.uart_inst0.N_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNI6B671_5_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10397\,
            in1 => \N__10424\,
            in2 => \N__10372\,
            in3 => \N__10451\,
            lcout => \DUT.uart_inst0.un2_rx_clk_divider_a_10\,
            ltout => \DUT.uart_inst0.un2_rx_clk_divider_a_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIKU472_10_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__9030\,
            in1 => \_gnd_net_\,
            in2 => \N__8062\,
            in3 => \N__9045\,
            lcout => \DUT.uart_inst0.rx_clk_divider_RNIKU472Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_1_0_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__7965\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8013\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.recv_state_RNO_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_0_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101110101"
        )
    port map (
            in0 => \N__8050\,
            in1 => \N__8426\,
            in2 => \N__8044\,
            in3 => \N__8370\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12133\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_0_1_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__8107\,
            in1 => \N__9128\,
            in2 => \N__8293\,
            in3 => \N__8545\,
            lcout => \DUT.uart_inst0.N_105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNI7H9R3_10_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8023\,
            in1 => \N__9046\,
            in2 => \N__9034\,
            in3 => \N__9192\,
            lcout => \DUT.uart_inst0.un2_rx_clk_divider_0\,
            ltout => \DUT.uart_inst0.un2_rx_clk_divider_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNI8UI86_3_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111000101"
        )
    port map (
            in0 => \N__8485\,
            in1 => \N__8079\,
            in2 => \N__8017\,
            in3 => \N__8475\,
            lcout => \DUT.uart_inst0.rx_countdown_8_i_o2_1_2\,
            ltout => \DUT.uart_inst0.rx_countdown_8_i_o2_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_4_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8291\,
            in1 => \N__8012\,
            in2 => \N__7975\,
            in3 => \N__8359\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.recv_state_RNO_0Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_4_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__11531\,
            in1 => \N__7969\,
            in2 => \N__7972\,
            in3 => \N__8292\,
            lcout => \DUT.uart_inst0.recv_stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNO_0_3_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101000101"
        )
    port map (
            in0 => \N__8288\,
            in1 => \N__9129\,
            in2 => \N__8512\,
            in3 => \N__8080\,
            lcout => \DUT.uart_inst0.N_102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.recv_state_RNO_0_5_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011111110111"
        )
    port map (
            in0 => \N__8263\,
            in1 => \N__11923\,
            in2 => \N__8240\,
            in3 => \N__8155\,
            lcout => \DUT.uart_inst0.recv_state_srsts_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_0_s1_c_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9062\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_16_16_0_\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_0_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_0_s1_c_RNIKPDT_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12997\,
            in2 => \N__8544\,
            in3 => \N__8092\,
            lcout => \DUT.uart_inst0.rx_countdown_3_s1_1\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_countdown_3_cry_0_s1\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_1_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_1_s1_THRU_LUT4_0_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13000\,
            in2 => \N__8313\,
            in3 => \N__8083\,
            lcout => \DUT.uart_inst0.rx_countdown_3_cry_1_s1_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_countdown_3_cry_1_s1\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_2_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_2_s1_c_RNIO52I_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12998\,
            in2 => \N__8508\,
            in3 => \N__8071\,
            lcout => \DUT.uart_inst0.rx_countdown_3_s1_3\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_countdown_3_cry_2_s1\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_3_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_3_s1_c_RNIQBCS_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13001\,
            in2 => \N__8463\,
            in3 => \N__8068\,
            lcout => \DUT.uart_inst0.rx_countdown_3_s1_4\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_countdown_3_cry_3_s1\,
            carryout => \DUT.uart_inst0.rx_countdown_3_cry_4_s1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_cry_4_s1_c_RNISHMM_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__9161\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8065\,
            lcout => \DUT.uart_inst0.rx_countdown_3_s1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_0_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__12999\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11276\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12124\,
            ce => 'H',
            sr => \N__12730\
        );

    \DUT.uart_inst0.rx_clk_divider_3_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110110111"
        )
    port map (
            in0 => \N__10501\,
            in1 => \N__11177\,
            in2 => \N__10530\,
            in3 => \N__9142\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12118\,
            ce => \N__11845\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_1_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11175\,
            in2 => \_gnd_net_\,
            in3 => \N__8554\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12118\,
            ce => \N__11845\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_3_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__11176\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8521\,
            lcout => \DUT.uart_inst0.rx_countdownZ1Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12118\,
            ce => \N__11845\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_RNIFRQU_3_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8459\,
            in2 => \_gnd_net_\,
            in3 => \N__8504\,
            lcout => \DUT.uart_inst0.rx_countdown_8_i_o2_1_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_4_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__9143\,
            in1 => \N__9092\,
            in2 => \N__8464\,
            in3 => \N__8476\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12118\,
            ce => \N__11845\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_2_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110001"
        )
    port map (
            in0 => \N__8443\,
            in1 => \N__8430\,
            in2 => \N__8383\,
            in3 => \N__8371\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12113\,
            ce => \N__11849\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_3_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12435\,
            in1 => \N__12217\,
            in2 => \N__10333\,
            in3 => \N__12387\,
            lcout => \DUT.uart_inst0.N_159\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNO_1_2_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110111111101"
        )
    port map (
            in0 => \N__12388\,
            in1 => \N__8773\,
            in2 => \N__12676\,
            in3 => \N__8689\,
            lcout => \DUT.uart_inst0.tx_bits_remaining_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_RNIBPK2_0_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11277\,
            in2 => \_gnd_net_\,
            in3 => \N__11257\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.un1_tx_clk_divider_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_RNITC2S1_0_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9529\,
            in1 => \N__9535\,
            in2 => \N__8701\,
            in3 => \N__9541\,
            lcout => \DUT.uart_inst0.un1_tx_clk_divider_0\,
            ltout => \DUT.uart_inst0.un1_tx_clk_divider_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNO_2_2_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000010"
        )
    port map (
            in0 => \N__8698\,
            in1 => \N__9885\,
            in2 => \N__8692\,
            in3 => \N__9755\,
            lcout => \DUT.uart_inst0.un1_tx_bits_remaining_axbxc2_N_4L5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoCount_RNIBPFM_1_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__11602\,
            in1 => \N__8682\,
            in2 => \N__8629\,
            in3 => \N__8577\,
            lcout => \DUT.fifo_tx_inst.rFifoCount_RNIBPFMZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNI18BH1_5_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__9504\,
            in1 => \N__12654\,
            in2 => \N__9456\,
            in3 => \N__9838\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g0_0_0_a3_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNIP6303_4_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__9339\,
            in1 => \N__8584\,
            in2 => \N__8590\,
            in3 => \N__9400\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g0_0_0_a3_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNI1BIT5_0_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010111010"
        )
    port map (
            in0 => \N__9682\,
            in1 => \N__9759\,
            in2 => \N__8587\,
            in3 => \N__11388\,
            lcout => \DUT.uart_inst0.N_152_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_0_3_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12443\,
            in1 => \N__12216\,
            in2 => \N__10331\,
            in3 => \N__12389\,
            lcout => \DUT.uart_inst0.N_159_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.rTransmit_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__12655\,
            in1 => \N__12324\,
            in2 => \_gnd_net_\,
            in3 => \N__8578\,
            lcout => \DUT.rTransmitZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12106\,
            ce => 'H',
            sr => \N__12493\
        );

    \DUT.uart_inst0.tx_countdown_RNO_0_5_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001011110000"
        )
    port map (
            in0 => \N__11399\,
            in1 => \N__9348\,
            in2 => \N__9462\,
            in3 => \N__9291\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_countdown_0_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_5_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011110000"
        )
    port map (
            in0 => \N__12328\,
            in1 => \_gnd_net_\,
            in2 => \N__8821\,
            in3 => \N__9968\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12101\,
            ce => \N__11862\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_RNO_1_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001110"
        )
    port map (
            in0 => \N__8818\,
            in1 => \N__11400\,
            in2 => \N__8796\,
            in3 => \N__9763\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.N_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001101"
        )
    port map (
            in0 => \N__10294\,
            in1 => \N__12670\,
            in2 => \N__8812\,
            in3 => \N__9688\,
            lcout => \P1A7_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12101\,
            ce => \N__11862\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_2_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111001011101"
        )
    port map (
            in0 => \N__8779\,
            in1 => \N__9967\,
            in2 => \N__12337\,
            in3 => \N__9401\,
            lcout => \DUT.uart_inst0.tx_countdownZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12101\,
            ce => \N__11862\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNO_3_2_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001101000111"
        )
    port map (
            in0 => \N__9451\,
            in1 => \N__12645\,
            in2 => \N__11623\,
            in3 => \N__9522\,
            lcout => \DUT.uart_inst0.un1_tx_bits_remaining_axbxc2_N_4L5_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100000110011"
        )
    port map (
            in0 => \N__8947\,
            in1 => \N__8764\,
            in2 => \N__8755\,
            in3 => \N__9676\,
            lcout => OPEN,
            ltout => \DUT.rFifoDatarx_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_RNO_0_1_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111000"
        )
    port map (
            in0 => \N__8739\,
            in1 => \N__12646\,
            in2 => \N__8728\,
            in3 => \N__10052\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_data_RNO_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_1_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__9991\,
            in1 => \N__10900\,
            in2 => \N__8725\,
            in3 => \N__8722\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12094\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_0_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__9870\,
            in1 => \N__8707\,
            in2 => \N__10906\,
            in3 => \N__9990\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12094\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_RNO_0_5_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010111000000"
        )
    port map (
            in0 => \N__10053\,
            in1 => \N__10093\,
            in2 => \N__12671\,
            in3 => \N__9019\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_data_RNO_0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_5_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__10899\,
            in1 => \N__9006\,
            in2 => \N__9010\,
            in3 => \N__9992\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12094\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8992\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12089\,
            ce => \N__10237\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8938\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12089\,
            ce => \N__10237\,
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8877\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12089\,
            ce => \N__10237\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_7_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__10905\,
            in1 => \N__8827\,
            in2 => \N__10116\,
            in3 => \N__10054\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12084\,
            ce => \N__9997\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_0_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11145\,
            in2 => \_gnd_net_\,
            in3 => \N__10152\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12138\,
            ce => \N__11832\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_6_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110011111"
        )
    port map (
            in0 => \N__10408\,
            in1 => \N__10426\,
            in2 => \N__11179\,
            in3 => \N__9145\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12138\,
            ce => \N__11832\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_7_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__10399\,
            in1 => \N__10381\,
            in2 => \_gnd_net_\,
            in3 => \N__11146\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12138\,
            ce => \N__11832\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_5_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110011111"
        )
    port map (
            in0 => \N__10435\,
            in1 => \N__10453\,
            in2 => \N__11178\,
            in3 => \N__9144\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12138\,
            ce => \N__11832\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIB99J_10_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10796\,
            in1 => \N__10769\,
            in2 => \N__10723\,
            in3 => \N__10745\,
            lcout => \DUT.uart_inst0.un2_rx_clk_divider_a_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_9_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100001000100"
        )
    port map (
            in0 => \N__10798\,
            in1 => \N__11163\,
            in2 => \_gnd_net_\,
            in3 => \N__10780\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12136\,
            ce => \N__11836\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_10_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000001010000"
        )
    port map (
            in0 => \N__10756\,
            in1 => \_gnd_net_\,
            in2 => \N__11180\,
            in3 => \N__10770\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12136\,
            ce => \N__11836\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_11_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__10746\,
            in1 => \N__10732\,
            in2 => \_gnd_net_\,
            in3 => \N__11156\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12136\,
            ce => \N__11836\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_12_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000001010000"
        )
    port map (
            in0 => \N__10721\,
            in1 => \_gnd_net_\,
            in2 => \N__11181\,
            in3 => \N__10705\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12136\,
            ce => \N__11836\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100001000100"
        )
    port map (
            in0 => \N__10570\,
            in1 => \N__11161\,
            in2 => \_gnd_net_\,
            in3 => \N__10588\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12136\,
            ce => \N__11836\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_16_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__11160\,
            in1 => \N__10597\,
            in2 => \_gnd_net_\,
            in3 => \N__10615\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12136\,
            ce => \N__11836\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_4_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100001000100"
        )
    port map (
            in0 => \N__10462\,
            in1 => \N__11162\,
            in2 => \_gnd_net_\,
            in3 => \N__10484\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12136\,
            ce => \N__11836\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNI3ALC_17_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10667\,
            in1 => \N__10694\,
            in2 => \N__11083\,
            in3 => \N__10640\,
            lcout => \DUT.uart_inst0.un2_rx_clk_divider_a_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_13_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010100000000"
        )
    port map (
            in0 => \N__10695\,
            in1 => \_gnd_net_\,
            in2 => \N__10681\,
            in3 => \N__11196\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12134\,
            ce => \N__11843\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_14_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000001010000"
        )
    port map (
            in0 => \N__10651\,
            in1 => \_gnd_net_\,
            in2 => \N__11203\,
            in3 => \N__10669\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12134\,
            ce => \N__11843\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_15_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010100000000"
        )
    port map (
            in0 => \N__10641\,
            in1 => \_gnd_net_\,
            in2 => \N__10627\,
            in3 => \N__11200\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12134\,
            ce => \N__11843\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIIDCT_2_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10556\,
            in2 => \N__10485\,
            in3 => \N__10526\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.un2_rx_clk_divider_a_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_RNIJI4K1_16_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__10613\,
            in1 => \N__10153\,
            in2 => \N__9199\,
            in3 => \N__10586\,
            lcout => \DUT.uart_inst0.un2_rx_clk_divider_a_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_2_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__10557\,
            in1 => \N__10543\,
            in2 => \_gnd_net_\,
            in3 => \N__11201\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12134\,
            ce => \N__11843\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_5_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000010"
        )
    port map (
            in0 => \N__9165\,
            in1 => \N__9131\,
            in2 => \N__9097\,
            in3 => \N__9181\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12130\,
            ce => \N__11846\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_countdown_0_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__9130\,
            in1 => \N__9093\,
            in2 => \_gnd_net_\,
            in3 => \N__9068\,
            lcout => \DUT.uart_inst0.rx_countdownZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12130\,
            ce => \N__11846\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_8_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__11174\,
            in1 => \N__10345\,
            in2 => \_gnd_net_\,
            in3 => \N__10367\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12130\,
            ce => \N__11846\,
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rRxF_n_1_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__12165\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fifo_inst.ftdi_output_inst.rRxF_nZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12130\,
            ce => \N__11846\,
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rTxE_n_RNIJBK2_1_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__9271\,
            in1 => \N__10195\,
            in2 => \_gnd_net_\,
            in3 => \N__10171\,
            lcout => \fifo_inst.ftdi_output_inst.N_86_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_2_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11930\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11292\,
            lcout => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12125\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rRxF_n_RNIHPJ8_1_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__12164\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11307\,
            lcout => \fifo_inst.ftdi_output_inst.N_95\,
            ltout => \fifo_inst.ftdi_output_inst.N_95_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_3_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9208\,
            in1 => \N__11935\,
            in2 => \N__9253\,
            in3 => \N__11329\,
            lcout => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12125\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_4_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001000000"
        )
    port map (
            in0 => \N__11012\,
            in1 => \N__11931\,
            in2 => \N__11043\,
            in3 => \N__9249\,
            lcout => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12125\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_RNO_0_0_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__9228\,
            in1 => \N__11036\,
            in2 => \N__11941\,
            in3 => \N__11011\,
            lcout => OPEN,
            ltout => \fifo_inst.ftdi_output_inst.m14_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_0_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111110001111"
        )
    port map (
            in0 => \N__11328\,
            in1 => \N__9217\,
            in2 => \N__9211\,
            in3 => \N__9207\,
            lcout => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12125\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_1_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011100001000"
        )
    port map (
            in0 => \N__9983\,
            in1 => \N__10871\,
            in2 => \N__12405\,
            in3 => \N__12224\,
            lcout => \DUT.uart_inst0.tx_bits_remainingZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12119\,
            ce => 'H',
            sr => \N__11632\
        );

    \DUT.uart_inst0.tx_bits_remaining_0_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__10869\,
            in1 => \N__12396\,
            in2 => \_gnd_net_\,
            in3 => \N__9982\,
            lcout => \DUT.uart_inst0.tx_bits_remainingZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12119\,
            ce => 'H',
            sr => \N__11632\
        );

    \DUT.uart_inst0.tx_bits_remaining_3_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__9985\,
            in1 => \N__10870\,
            in2 => \N__12352\,
            in3 => \N__10327\,
            lcout => \DUT.uart_inst0.tx_bits_remainingZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12119\,
            ce => 'H',
            sr => \N__11632\
        );

    \DUT.uart_inst0.tx_bits_remaining_2_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010011010"
        )
    port map (
            in0 => \N__12442\,
            in1 => \N__9984\,
            in2 => \N__12190\,
            in3 => \N__9547\,
            lcout => \DUT.uart_inst0.tx_bits_remainingZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12119\,
            ce => 'H',
            sr => \N__11632\
        );

    \DUT.uart_inst0.tx_clk_divider_RNI2V95_2_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11739\,
            in1 => \N__11758\,
            in2 => \N__11236\,
            in3 => \N__11217\,
            lcout => \DUT.uart_inst0.un1_tx_clk_divider_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_13_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12762\,
            in1 => \N__11724\,
            in2 => \N__12745\,
            in3 => \N__11709\,
            lcout => \DUT.uart_inst0.un1_tx_clk_divider_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_8_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11694\,
            in1 => \N__11679\,
            in2 => \N__11650\,
            in3 => \N__11664\,
            lcout => \DUT.uart_inst0.un1_tx_clk_divider_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNIJ3F33_3_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000000011"
        )
    port map (
            in0 => \N__9767\,
            in1 => \N__9851\,
            in2 => \N__9523\,
            in3 => \N__11376\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_data_i_m_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNIHJJ88_5_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__9452\,
            in1 => \N__9409\,
            in2 => \N__9352\,
            in3 => \N__9277\,
            lcout => \DUT.uart_inst0.N_345_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNIBSRA4_4_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110111101110"
        )
    port map (
            in0 => \N__9766\,
            in1 => \N__9349\,
            in2 => \N__9295\,
            in3 => \N__11375\,
            lcout => \DUT.uart_inst0.tx_state_ns_0_o3_1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_RNO_0_6_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__12619\,
            in1 => \N__10132\,
            in2 => \N__10120\,
            in3 => \N__10043\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_data_RNO_0Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_6_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__10898\,
            in1 => \N__10089\,
            in2 => \N__10096\,
            in3 => \N__9988\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_RNO_0_3_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011100100"
        )
    port map (
            in0 => \N__12618\,
            in1 => \N__9553\,
            in2 => \N__10074\,
            in3 => \N__10042\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.tx_data_RNO_0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_data_3_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__10897\,
            in1 => \N__9903\,
            in2 => \N__10000\,
            in3 => \N__9987\,
            lcout => \DUT.uart_inst0.tx_dataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_RNO_5_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__12617\,
            in1 => \N__9889\,
            in2 => \N__9874\,
            in3 => \N__9856\,
            lcout => OPEN,
            ltout => \DUT.uart_inst0.g0_i_a4_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_RNO_2_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000100000"
        )
    port map (
            in0 => \N__9784\,
            in1 => \N__9772\,
            in2 => \N__9691\,
            in3 => \N__11401\,
            lcout => \DUT.uart_inst0.N_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNI5H8K_0_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11586\,
            in2 => \_gnd_net_\,
            in3 => \N__12591\,
            lcout => \DUT.uart_inst0.N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__10246\,
            in1 => \N__9675\,
            in2 => \N__9577\,
            in3 => \N__9562\,
            lcout => \DUT.rFifoDatarx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNIB46K_3_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__12614\,
            in1 => \N__10332\,
            in2 => \_gnd_net_\,
            in3 => \N__12444\,
            lcout => \DUT.uart_inst0.tx_state_ns_i_i_a2_0_0_0\,
            ltout => \DUT.uart_inst0.tx_state_ns_i_i_a2_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNICODU_1_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12235\,
            in2 => \N__10297\,
            in3 => \N__12404\,
            lcout => \DUT.uart_inst0.tx_state_ns_i_i_a2_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_RNO_0_0_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__12320\,
            in1 => \N__11610\,
            in2 => \_gnd_net_\,
            in3 => \N__12616\,
            lcout => \DUT.uart_inst0.tx_state_ns_i_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_out_RNO_0_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__11609\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12319\,
            lcout => \DUT.uart_inst0.g0_i_a4_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_countdown_RNO_5_3_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__12318\,
            in1 => \N__11608\,
            in2 => \_gnd_net_\,
            in3 => \N__12615\,
            lcout => \DUT.uart_inst0.d_N_5_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10276\,
            lcout => \DUT.fifo_tx_inst.rFifoData_ram2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12095\,
            ce => \N__10233\,
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rTxE_n_1_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10167\,
            lcout => \fifo_inst.ftdi_output_inst.rTxE_nZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12090\,
            ce => \N__11866\,
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rTxE_n_0_LC_17_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10183\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \fifo_inst.ftdi_output_inst.rTxE_nZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12085\,
            ce => \N__11867\,
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10151\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_13_0_\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10587\,
            in2 => \N__12991\,
            in3 => \N__10564\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_0\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10561\,
            in2 => \N__12995\,
            in3 => \N__10534\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_1\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_2_THRU_LUT4_0_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10531\,
            in2 => \N__12992\,
            in3 => \N__10489\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_2\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12947\,
            in2 => \N__10486\,
            in3 => \N__10456\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_3\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_4_THRU_LUT4_0_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10452\,
            in2 => \N__12993\,
            in3 => \N__10429\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_4\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_5_THRU_LUT4_0_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10425\,
            in2 => \N__12996\,
            in3 => \N__10402\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_5\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10398\,
            in2 => \N__12994\,
            in3 => \N__10375\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_6\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10371\,
            in2 => \N__12989\,
            in3 => \N__10336\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_18_14_0_\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10797\,
            in2 => \N__12986\,
            in3 => \N__10774\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_8\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_LUT4_0_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10771\,
            in2 => \N__12990\,
            in3 => \N__10750\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_9\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_LUT4_0_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10747\,
            in2 => \N__12983\,
            in3 => \N__10726\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_10\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_LUT4_0_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10722\,
            in2 => \N__12987\,
            in3 => \N__10699\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_11\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_LUT4_0_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10696\,
            in2 => \N__12984\,
            in3 => \N__10672\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_12\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_LUT4_0_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10668\,
            in2 => \N__12988\,
            in3 => \N__10645\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_13\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_LUT4_0_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10642\,
            in2 => \N__12985\,
            in3 => \N__10618\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.rx_clk_divider_1_cry_14\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_LUT4_0_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10614\,
            in2 => \N__12982\,
            in3 => \N__10591\,
            lcout => \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_18_15_0_\,
            carryout => \DUT.uart_inst0.rx_clk_divider_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.rx_clk_divider_17_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100001000100"
        )
    port map (
            in0 => \N__11082\,
            in1 => \N__11202\,
            in2 => \_gnd_net_\,
            in3 => \N__11086\,
            lcout => \DUT.uart_inst0.rx_clk_dividerZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12137\,
            ce => \N__11847\,
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.oRamRdAddr_0_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__10963\,
            in1 => \N__11035\,
            in2 => \N__11940\,
            in3 => \N__11014\,
            lcout => \fifo_inst.wRamRdAddr_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12135\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.oRamRdAddr_2_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__10931\,
            in1 => \N__10965\,
            in2 => \N__11061\,
            in3 => \N__10981\,
            lcout => \fifo_inst.wRamRdAddr_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12135\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_RNIBT9K_4_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__11929\,
            in1 => \N__11034\,
            in2 => \_gnd_net_\,
            in3 => \N__11013\,
            lcout => \fifo_inst.ftdi_output_inst.N_3_0\,
            ltout => \fifo_inst.ftdi_output_inst.N_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.oRamRdAddr_1_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110101001101010"
        )
    port map (
            in0 => \N__10932\,
            in1 => \N__10964\,
            in2 => \N__10948\,
            in3 => \_gnd_net_\,
            lcout => \fifo_inst.wRamRdAddr_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12135\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_esr_1_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__10918\,
            in1 => \N__12223\,
            in2 => \_gnd_net_\,
            in3 => \N__12400\,
            lcout => \DUT.tx_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12131\,
            ce => \N__10804\,
            sr => \N__12495\
        );

    \CONSTANT_ONE_LUT4_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_esr_RNICLU7_1_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11936\,
            in2 => \_gnd_net_\,
            in3 => \N__12266\,
            lcout => \DUT.uart_inst0.tx_state_0_sqmuxa_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_esr_RNO_1_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10831\,
            in2 => \_gnd_net_\,
            in3 => \N__12693\,
            lcout => \DUT.uart_inst0.N_345_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_esr_RNIH67S_1_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11937\,
            in2 => \_gnd_net_\,
            in3 => \N__11542\,
            lcout => \DUT.uart_inst0.tx_bits_remaining_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_esr_RNILOSP_1_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__12265\,
            in1 => \N__11622\,
            in2 => \_gnd_net_\,
            in3 => \N__12653\,
            lcout => \DUT.uart_inst0.tx_clk_divider_0_sqmuxa\,
            ltout => \DUT.uart_inst0.tx_clk_divider_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_state_esr_RNIEJ9O2_1_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__11494\,
            in1 => \_gnd_net_\,
            in2 => \N__11404\,
            in3 => \N__11397\,
            lcout => \DUT.uart_inst0.tx_clk_divider_1_sqmuxa_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rFifoState_1_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101000000000"
        )
    port map (
            in0 => \N__11322\,
            in1 => \N__11311\,
            in2 => \N__12166\,
            in3 => \N__11938\,
            lcout => \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12126\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11281\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_19_0_\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_clk_divider_1_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11253\,
            in2 => \N__12892\,
            in3 => \N__11239\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_1\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_0\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_1\,
            clk => \N__12120\,
            ce => 'H',
            sr => \N__12716\
        );

    \DUT.uart_inst0.tx_clk_divider_2_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11235\,
            in2 => \N__12896\,
            in3 => \N__11221\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_2\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_1\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_2\,
            clk => \N__12120\,
            ce => 'H',
            sr => \N__12716\
        );

    \DUT.uart_inst0.tx_clk_divider_3_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11218\,
            in2 => \N__12893\,
            in3 => \N__11206\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_3\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_2\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_3\,
            clk => \N__12120\,
            ce => 'H',
            sr => \N__12716\
        );

    \DUT.uart_inst0.tx_clk_divider_4_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11757\,
            in2 => \N__12897\,
            in3 => \N__11743\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_4\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_3\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_4\,
            clk => \N__12120\,
            ce => 'H',
            sr => \N__12716\
        );

    \DUT.uart_inst0.tx_clk_divider_5_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11740\,
            in2 => \N__12894\,
            in3 => \N__11728\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_5\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_4\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_5\,
            clk => \N__12120\,
            ce => 'H',
            sr => \N__12716\
        );

    \DUT.uart_inst0.tx_clk_divider_6_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11725\,
            in2 => \N__12898\,
            in3 => \N__11713\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_6\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_5\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_6\,
            clk => \N__12120\,
            ce => 'H',
            sr => \N__12716\
        );

    \DUT.uart_inst0.tx_clk_divider_7_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11710\,
            in2 => \N__12895\,
            in3 => \N__11698\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_7\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_6\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_7\,
            clk => \N__12120\,
            ce => 'H',
            sr => \N__12716\
        );

    \DUT.uart_inst0.tx_clk_divider_8_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11695\,
            in2 => \N__12979\,
            in3 => \N__11683\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_18_20_0_\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_8\,
            clk => \N__12114\,
            ce => 'H',
            sr => \N__12729\
        );

    \DUT.uart_inst0.tx_clk_divider_9_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11680\,
            in2 => \N__12981\,
            in3 => \N__11668\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_9\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_8\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_9\,
            clk => \N__12114\,
            ce => 'H',
            sr => \N__12729\
        );

    \DUT.uart_inst0.tx_clk_divider_10_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11665\,
            in2 => \N__12977\,
            in3 => \N__11653\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_10\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_9\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_10\,
            clk => \N__12114\,
            ce => 'H',
            sr => \N__12729\
        );

    \DUT.uart_inst0.tx_clk_divider_11_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11649\,
            in2 => \N__12980\,
            in3 => \N__11635\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_11\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_10\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_11\,
            clk => \N__12114\,
            ce => 'H',
            sr => \N__12729\
        );

    \DUT.uart_inst0.tx_clk_divider_12_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12763\,
            in2 => \N__12978\,
            in3 => \N__12751\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_12\,
            ltout => OPEN,
            carryin => \DUT.uart_inst0.tx_clk_divider_cry_11\,
            carryout => \DUT.uart_inst0.tx_clk_divider_cry_12\,
            clk => \N__12114\,
            ce => 'H',
            sr => \N__12729\
        );

    \DUT.uart_inst0.tx_clk_divider_13_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12744\,
            in2 => \_gnd_net_\,
            in3 => \N__12748\,
            lcout => \DUT.uart_inst0.tx_clk_dividerZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12114\,
            ce => 'H',
            sr => \N__12729\
        );

    \DUT.uart_inst0.tx_state_0_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__12703\,
            in1 => \N__12697\,
            in2 => \_gnd_net_\,
            in3 => \N__12682\,
            lcout => \DUT.tx_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12108\,
            ce => 'H',
            sr => \N__12494\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_18_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__12234\,
            in1 => \N__12445\,
            in2 => \_gnd_net_\,
            in3 => \N__12406\,
            lcout => \DUT.uart_inst0.tx_bits_remaining_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DUT.uart_inst0.tx_bits_remaining_RNO_0_2_LC_18_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__11939\,
            in1 => \N__12321\,
            in2 => \_gnd_net_\,
            in3 => \N__12233\,
            lcout => \DUT.uart_inst0.tx_bits_remaining_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \fifo_inst.ftdi_output_inst.rRxF_n_0_LC_18_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12175\,
            lcout => \fifo_inst.ftdi_output_inst.rRxF_nZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12096\,
            ce => \N__11868\,
            sr => \_gnd_net_\
        );
end \INTERFACE\;
