// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Mar 29 2020 02:25:19

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    ioFifoData,
    P1A9,
    P1A1,
    P1A8,
    oRx_n,
    P1A7,
    P1A3,
    iTxE_n,
    iRxF_n,
    iClk,
    P1A2,
    BTN_N,
    BTN1,
    oTx_n,
    P1A4);

    inout [7:0] ioFifoData;
    output P1A9;
    input P1A1;
    output P1A8;
    output oRx_n;
    output P1A7;
    output P1A3;
    input iTxE_n;
    input iRxF_n;
    input iClk;
    output P1A2;
    input BTN_N;
    input BTN1;
    output oTx_n;
    output P1A4;

    wire N__15651;
    wire N__15637;
    wire N__15636;
    wire N__15635;
    wire N__15628;
    wire N__15627;
    wire N__15626;
    wire N__15619;
    wire N__15618;
    wire N__15617;
    wire N__15610;
    wire N__15609;
    wire N__15608;
    wire N__15601;
    wire N__15600;
    wire N__15599;
    wire N__15592;
    wire N__15591;
    wire N__15590;
    wire N__15583;
    wire N__15582;
    wire N__15581;
    wire N__15574;
    wire N__15573;
    wire N__15572;
    wire N__15565;
    wire N__15564;
    wire N__15563;
    wire N__15556;
    wire N__15555;
    wire N__15554;
    wire N__15547;
    wire N__15546;
    wire N__15545;
    wire N__15538;
    wire N__15537;
    wire N__15536;
    wire N__15529;
    wire N__15528;
    wire N__15527;
    wire N__15520;
    wire N__15519;
    wire N__15518;
    wire N__15511;
    wire N__15510;
    wire N__15509;
    wire N__15502;
    wire N__15501;
    wire N__15500;
    wire N__15493;
    wire N__15492;
    wire N__15491;
    wire N__15484;
    wire N__15483;
    wire N__15482;
    wire N__15475;
    wire N__15474;
    wire N__15473;
    wire N__15466;
    wire N__15465;
    wire N__15464;
    wire N__15447;
    wire N__15444;
    wire N__15441;
    wire N__15438;
    wire N__15435;
    wire N__15432;
    wire N__15429;
    wire N__15426;
    wire N__15423;
    wire N__15422;
    wire N__15421;
    wire N__15418;
    wire N__15417;
    wire N__15414;
    wire N__15411;
    wire N__15410;
    wire N__15409;
    wire N__15408;
    wire N__15403;
    wire N__15396;
    wire N__15393;
    wire N__15392;
    wire N__15389;
    wire N__15388;
    wire N__15387;
    wire N__15384;
    wire N__15381;
    wire N__15376;
    wire N__15369;
    wire N__15360;
    wire N__15359;
    wire N__15358;
    wire N__15357;
    wire N__15356;
    wire N__15351;
    wire N__15344;
    wire N__15343;
    wire N__15342;
    wire N__15341;
    wire N__15340;
    wire N__15339;
    wire N__15336;
    wire N__15333;
    wire N__15328;
    wire N__15321;
    wire N__15312;
    wire N__15309;
    wire N__15306;
    wire N__15303;
    wire N__15302;
    wire N__15299;
    wire N__15296;
    wire N__15291;
    wire N__15290;
    wire N__15287;
    wire N__15286;
    wire N__15285;
    wire N__15284;
    wire N__15283;
    wire N__15282;
    wire N__15281;
    wire N__15280;
    wire N__15279;
    wire N__15278;
    wire N__15275;
    wire N__15266;
    wire N__15263;
    wire N__15260;
    wire N__15253;
    wire N__15250;
    wire N__15249;
    wire N__15248;
    wire N__15245;
    wire N__15242;
    wire N__15241;
    wire N__15240;
    wire N__15237;
    wire N__15236;
    wire N__15233;
    wire N__15232;
    wire N__15231;
    wire N__15230;
    wire N__15229;
    wire N__15226;
    wire N__15225;
    wire N__15224;
    wire N__15223;
    wire N__15220;
    wire N__15219;
    wire N__15218;
    wire N__15177;
    wire N__15174;
    wire N__15171;
    wire N__15168;
    wire N__15167;
    wire N__15166;
    wire N__15163;
    wire N__15160;
    wire N__15157;
    wire N__15154;
    wire N__15151;
    wire N__15148;
    wire N__15147;
    wire N__15146;
    wire N__15143;
    wire N__15140;
    wire N__15137;
    wire N__15134;
    wire N__15131;
    wire N__15120;
    wire N__15117;
    wire N__15114;
    wire N__15111;
    wire N__15110;
    wire N__15107;
    wire N__15106;
    wire N__15103;
    wire N__15100;
    wire N__15097;
    wire N__15094;
    wire N__15089;
    wire N__15086;
    wire N__15083;
    wire N__15082;
    wire N__15081;
    wire N__15076;
    wire N__15073;
    wire N__15070;
    wire N__15063;
    wire N__15060;
    wire N__15057;
    wire N__15054;
    wire N__15053;
    wire N__15052;
    wire N__15051;
    wire N__15050;
    wire N__15049;
    wire N__15048;
    wire N__15047;
    wire N__15046;
    wire N__15045;
    wire N__15044;
    wire N__15043;
    wire N__15042;
    wire N__15041;
    wire N__15040;
    wire N__15039;
    wire N__15038;
    wire N__15037;
    wire N__15036;
    wire N__15035;
    wire N__15034;
    wire N__15033;
    wire N__15032;
    wire N__15031;
    wire N__15030;
    wire N__15029;
    wire N__15028;
    wire N__15027;
    wire N__15026;
    wire N__15025;
    wire N__15024;
    wire N__15023;
    wire N__15022;
    wire N__15021;
    wire N__15020;
    wire N__15019;
    wire N__15018;
    wire N__15017;
    wire N__15016;
    wire N__15015;
    wire N__15014;
    wire N__15013;
    wire N__15012;
    wire N__15011;
    wire N__15010;
    wire N__15009;
    wire N__15008;
    wire N__15007;
    wire N__15006;
    wire N__15005;
    wire N__15004;
    wire N__15003;
    wire N__15002;
    wire N__15001;
    wire N__15000;
    wire N__14999;
    wire N__14998;
    wire N__14997;
    wire N__14996;
    wire N__14995;
    wire N__14994;
    wire N__14871;
    wire N__14868;
    wire N__14867;
    wire N__14866;
    wire N__14863;
    wire N__14860;
    wire N__14859;
    wire N__14856;
    wire N__14853;
    wire N__14850;
    wire N__14847;
    wire N__14844;
    wire N__14839;
    wire N__14836;
    wire N__14833;
    wire N__14826;
    wire N__14825;
    wire N__14824;
    wire N__14823;
    wire N__14820;
    wire N__14819;
    wire N__14818;
    wire N__14817;
    wire N__14816;
    wire N__14815;
    wire N__14814;
    wire N__14813;
    wire N__14812;
    wire N__14809;
    wire N__14806;
    wire N__14789;
    wire N__14786;
    wire N__14783;
    wire N__14780;
    wire N__14777;
    wire N__14774;
    wire N__14773;
    wire N__14770;
    wire N__14767;
    wire N__14764;
    wire N__14761;
    wire N__14758;
    wire N__14755;
    wire N__14750;
    wire N__14747;
    wire N__14744;
    wire N__14737;
    wire N__14730;
    wire N__14727;
    wire N__14724;
    wire N__14723;
    wire N__14720;
    wire N__14717;
    wire N__14714;
    wire N__14711;
    wire N__14710;
    wire N__14707;
    wire N__14704;
    wire N__14701;
    wire N__14694;
    wire N__14693;
    wire N__14692;
    wire N__14687;
    wire N__14684;
    wire N__14679;
    wire N__14676;
    wire N__14673;
    wire N__14670;
    wire N__14669;
    wire N__14666;
    wire N__14663;
    wire N__14658;
    wire N__14655;
    wire N__14652;
    wire N__14649;
    wire N__14648;
    wire N__14647;
    wire N__14644;
    wire N__14637;
    wire N__14636;
    wire N__14633;
    wire N__14630;
    wire N__14627;
    wire N__14624;
    wire N__14621;
    wire N__14618;
    wire N__14613;
    wire N__14610;
    wire N__14607;
    wire N__14604;
    wire N__14603;
    wire N__14600;
    wire N__14597;
    wire N__14592;
    wire N__14589;
    wire N__14588;
    wire N__14585;
    wire N__14582;
    wire N__14577;
    wire N__14576;
    wire N__14575;
    wire N__14574;
    wire N__14573;
    wire N__14572;
    wire N__14571;
    wire N__14568;
    wire N__14567;
    wire N__14566;
    wire N__14565;
    wire N__14564;
    wire N__14563;
    wire N__14562;
    wire N__14561;
    wire N__14558;
    wire N__14557;
    wire N__14556;
    wire N__14553;
    wire N__14552;
    wire N__14551;
    wire N__14550;
    wire N__14549;
    wire N__14548;
    wire N__14547;
    wire N__14546;
    wire N__14543;
    wire N__14540;
    wire N__14537;
    wire N__14530;
    wire N__14527;
    wire N__14522;
    wire N__14517;
    wire N__14514;
    wire N__14511;
    wire N__14508;
    wire N__14505;
    wire N__14502;
    wire N__14497;
    wire N__14492;
    wire N__14489;
    wire N__14486;
    wire N__14483;
    wire N__14480;
    wire N__14477;
    wire N__14474;
    wire N__14471;
    wire N__14468;
    wire N__14465;
    wire N__14462;
    wire N__14461;
    wire N__14460;
    wire N__14457;
    wire N__14456;
    wire N__14453;
    wire N__14452;
    wire N__14451;
    wire N__14450;
    wire N__14447;
    wire N__14444;
    wire N__14443;
    wire N__14440;
    wire N__14437;
    wire N__14436;
    wire N__14435;
    wire N__14432;
    wire N__14429;
    wire N__14428;
    wire N__14425;
    wire N__14422;
    wire N__14421;
    wire N__14364;
    wire N__14361;
    wire N__14358;
    wire N__14357;
    wire N__14356;
    wire N__14353;
    wire N__14348;
    wire N__14343;
    wire N__14340;
    wire N__14337;
    wire N__14336;
    wire N__14333;
    wire N__14330;
    wire N__14325;
    wire N__14324;
    wire N__14323;
    wire N__14322;
    wire N__14315;
    wire N__14312;
    wire N__14307;
    wire N__14304;
    wire N__14301;
    wire N__14298;
    wire N__14295;
    wire N__14292;
    wire N__14289;
    wire N__14286;
    wire N__14283;
    wire N__14280;
    wire N__14277;
    wire N__14274;
    wire N__14271;
    wire N__14268;
    wire N__14267;
    wire N__14266;
    wire N__14263;
    wire N__14260;
    wire N__14257;
    wire N__14254;
    wire N__14251;
    wire N__14248;
    wire N__14245;
    wire N__14240;
    wire N__14235;
    wire N__14232;
    wire N__14229;
    wire N__14226;
    wire N__14225;
    wire N__14222;
    wire N__14219;
    wire N__14216;
    wire N__14215;
    wire N__14212;
    wire N__14209;
    wire N__14206;
    wire N__14203;
    wire N__14198;
    wire N__14197;
    wire N__14194;
    wire N__14191;
    wire N__14188;
    wire N__14181;
    wire N__14178;
    wire N__14175;
    wire N__14174;
    wire N__14173;
    wire N__14172;
    wire N__14169;
    wire N__14162;
    wire N__14157;
    wire N__14156;
    wire N__14153;
    wire N__14150;
    wire N__14149;
    wire N__14146;
    wire N__14141;
    wire N__14136;
    wire N__14133;
    wire N__14130;
    wire N__14127;
    wire N__14126;
    wire N__14123;
    wire N__14120;
    wire N__14115;
    wire N__14114;
    wire N__14113;
    wire N__14110;
    wire N__14105;
    wire N__14100;
    wire N__14097;
    wire N__14094;
    wire N__14091;
    wire N__14088;
    wire N__14087;
    wire N__14086;
    wire N__14083;
    wire N__14080;
    wire N__14077;
    wire N__14074;
    wire N__14071;
    wire N__14068;
    wire N__14067;
    wire N__14066;
    wire N__14063;
    wire N__14060;
    wire N__14057;
    wire N__14054;
    wire N__14051;
    wire N__14040;
    wire N__14037;
    wire N__14034;
    wire N__14031;
    wire N__14028;
    wire N__14025;
    wire N__14022;
    wire N__14019;
    wire N__14016;
    wire N__14015;
    wire N__14012;
    wire N__14011;
    wire N__14008;
    wire N__14007;
    wire N__14006;
    wire N__14005;
    wire N__14002;
    wire N__13991;
    wire N__13986;
    wire N__13983;
    wire N__13980;
    wire N__13977;
    wire N__13976;
    wire N__13975;
    wire N__13972;
    wire N__13969;
    wire N__13968;
    wire N__13965;
    wire N__13958;
    wire N__13953;
    wire N__13950;
    wire N__13949;
    wire N__13948;
    wire N__13947;
    wire N__13944;
    wire N__13937;
    wire N__13932;
    wire N__13929;
    wire N__13928;
    wire N__13927;
    wire N__13926;
    wire N__13925;
    wire N__13924;
    wire N__13921;
    wire N__13910;
    wire N__13905;
    wire N__13902;
    wire N__13901;
    wire N__13898;
    wire N__13897;
    wire N__13896;
    wire N__13895;
    wire N__13894;
    wire N__13891;
    wire N__13888;
    wire N__13879;
    wire N__13872;
    wire N__13869;
    wire N__13866;
    wire N__13863;
    wire N__13860;
    wire N__13857;
    wire N__13854;
    wire N__13851;
    wire N__13848;
    wire N__13845;
    wire N__13842;
    wire N__13839;
    wire N__13836;
    wire N__13833;
    wire N__13830;
    wire N__13827;
    wire N__13824;
    wire N__13821;
    wire N__13818;
    wire N__13817;
    wire N__13816;
    wire N__13815;
    wire N__13814;
    wire N__13813;
    wire N__13812;
    wire N__13811;
    wire N__13810;
    wire N__13809;
    wire N__13808;
    wire N__13807;
    wire N__13802;
    wire N__13795;
    wire N__13792;
    wire N__13785;
    wire N__13778;
    wire N__13773;
    wire N__13764;
    wire N__13761;
    wire N__13758;
    wire N__13755;
    wire N__13752;
    wire N__13749;
    wire N__13746;
    wire N__13743;
    wire N__13740;
    wire N__13739;
    wire N__13738;
    wire N__13737;
    wire N__13736;
    wire N__13735;
    wire N__13734;
    wire N__13733;
    wire N__13732;
    wire N__13731;
    wire N__13730;
    wire N__13729;
    wire N__13726;
    wire N__13723;
    wire N__13722;
    wire N__13721;
    wire N__13720;
    wire N__13717;
    wire N__13716;
    wire N__13713;
    wire N__13710;
    wire N__13709;
    wire N__13708;
    wire N__13705;
    wire N__13704;
    wire N__13701;
    wire N__13700;
    wire N__13697;
    wire N__13684;
    wire N__13671;
    wire N__13668;
    wire N__13661;
    wire N__13654;
    wire N__13647;
    wire N__13638;
    wire N__13635;
    wire N__13632;
    wire N__13631;
    wire N__13630;
    wire N__13627;
    wire N__13624;
    wire N__13621;
    wire N__13616;
    wire N__13613;
    wire N__13612;
    wire N__13609;
    wire N__13606;
    wire N__13603;
    wire N__13596;
    wire N__13593;
    wire N__13590;
    wire N__13589;
    wire N__13588;
    wire N__13585;
    wire N__13582;
    wire N__13579;
    wire N__13574;
    wire N__13571;
    wire N__13570;
    wire N__13569;
    wire N__13566;
    wire N__13563;
    wire N__13560;
    wire N__13557;
    wire N__13548;
    wire N__13545;
    wire N__13542;
    wire N__13539;
    wire N__13536;
    wire N__13535;
    wire N__13534;
    wire N__13531;
    wire N__13528;
    wire N__13525;
    wire N__13522;
    wire N__13517;
    wire N__13516;
    wire N__13515;
    wire N__13512;
    wire N__13509;
    wire N__13506;
    wire N__13503;
    wire N__13494;
    wire N__13491;
    wire N__13488;
    wire N__13487;
    wire N__13484;
    wire N__13481;
    wire N__13480;
    wire N__13475;
    wire N__13472;
    wire N__13469;
    wire N__13468;
    wire N__13467;
    wire N__13464;
    wire N__13461;
    wire N__13458;
    wire N__13455;
    wire N__13446;
    wire N__13443;
    wire N__13440;
    wire N__13437;
    wire N__13434;
    wire N__13433;
    wire N__13430;
    wire N__13427;
    wire N__13426;
    wire N__13423;
    wire N__13420;
    wire N__13417;
    wire N__13416;
    wire N__13415;
    wire N__13412;
    wire N__13409;
    wire N__13406;
    wire N__13403;
    wire N__13400;
    wire N__13389;
    wire N__13386;
    wire N__13383;
    wire N__13380;
    wire N__13377;
    wire N__13374;
    wire N__13371;
    wire N__13368;
    wire N__13367;
    wire N__13366;
    wire N__13365;
    wire N__13362;
    wire N__13359;
    wire N__13356;
    wire N__13353;
    wire N__13344;
    wire N__13341;
    wire N__13338;
    wire N__13337;
    wire N__13336;
    wire N__13335;
    wire N__13334;
    wire N__13333;
    wire N__13332;
    wire N__13331;
    wire N__13314;
    wire N__13311;
    wire N__13308;
    wire N__13305;
    wire N__13302;
    wire N__13299;
    wire N__13296;
    wire N__13293;
    wire N__13292;
    wire N__13289;
    wire N__13286;
    wire N__13285;
    wire N__13282;
    wire N__13279;
    wire N__13276;
    wire N__13275;
    wire N__13268;
    wire N__13265;
    wire N__13260;
    wire N__13257;
    wire N__13254;
    wire N__13251;
    wire N__13248;
    wire N__13245;
    wire N__13242;
    wire N__13239;
    wire N__13236;
    wire N__13233;
    wire N__13230;
    wire N__13227;
    wire N__13224;
    wire N__13221;
    wire N__13218;
    wire N__13215;
    wire N__13212;
    wire N__13209;
    wire N__13206;
    wire N__13203;
    wire N__13200;
    wire N__13197;
    wire N__13194;
    wire N__13191;
    wire N__13188;
    wire N__13185;
    wire N__13182;
    wire N__13179;
    wire N__13176;
    wire N__13173;
    wire N__13170;
    wire N__13167;
    wire N__13164;
    wire N__13161;
    wire N__13158;
    wire N__13155;
    wire N__13152;
    wire N__13149;
    wire N__13146;
    wire N__13143;
    wire N__13140;
    wire N__13137;
    wire N__13134;
    wire N__13131;
    wire N__13128;
    wire N__13125;
    wire N__13122;
    wire N__13119;
    wire N__13116;
    wire N__13115;
    wire N__13112;
    wire N__13109;
    wire N__13108;
    wire N__13105;
    wire N__13104;
    wire N__13101;
    wire N__13098;
    wire N__13095;
    wire N__13092;
    wire N__13087;
    wire N__13082;
    wire N__13077;
    wire N__13074;
    wire N__13071;
    wire N__13068;
    wire N__13065;
    wire N__13062;
    wire N__13059;
    wire N__13058;
    wire N__13055;
    wire N__13052;
    wire N__13051;
    wire N__13050;
    wire N__13047;
    wire N__13044;
    wire N__13041;
    wire N__13038;
    wire N__13031;
    wire N__13028;
    wire N__13023;
    wire N__13020;
    wire N__13017;
    wire N__13014;
    wire N__13011;
    wire N__13008;
    wire N__13007;
    wire N__13004;
    wire N__13001;
    wire N__13000;
    wire N__12999;
    wire N__12996;
    wire N__12993;
    wire N__12990;
    wire N__12987;
    wire N__12984;
    wire N__12979;
    wire N__12976;
    wire N__12969;
    wire N__12966;
    wire N__12963;
    wire N__12960;
    wire N__12959;
    wire N__12958;
    wire N__12955;
    wire N__12952;
    wire N__12949;
    wire N__12948;
    wire N__12945;
    wire N__12942;
    wire N__12939;
    wire N__12936;
    wire N__12933;
    wire N__12930;
    wire N__12927;
    wire N__12924;
    wire N__12915;
    wire N__12912;
    wire N__12909;
    wire N__12906;
    wire N__12903;
    wire N__12902;
    wire N__12899;
    wire N__12896;
    wire N__12895;
    wire N__12894;
    wire N__12891;
    wire N__12888;
    wire N__12885;
    wire N__12882;
    wire N__12879;
    wire N__12874;
    wire N__12871;
    wire N__12868;
    wire N__12865;
    wire N__12862;
    wire N__12855;
    wire N__12852;
    wire N__12849;
    wire N__12846;
    wire N__12843;
    wire N__12840;
    wire N__12839;
    wire N__12838;
    wire N__12837;
    wire N__12834;
    wire N__12831;
    wire N__12828;
    wire N__12825;
    wire N__12816;
    wire N__12813;
    wire N__12810;
    wire N__12807;
    wire N__12804;
    wire N__12801;
    wire N__12798;
    wire N__12795;
    wire N__12792;
    wire N__12789;
    wire N__12786;
    wire N__12783;
    wire N__12780;
    wire N__12777;
    wire N__12774;
    wire N__12771;
    wire N__12768;
    wire N__12765;
    wire N__12762;
    wire N__12759;
    wire N__12756;
    wire N__12753;
    wire N__12750;
    wire N__12747;
    wire N__12744;
    wire N__12741;
    wire N__12738;
    wire N__12735;
    wire N__12732;
    wire N__12729;
    wire N__12726;
    wire N__12723;
    wire N__12720;
    wire N__12717;
    wire N__12714;
    wire N__12711;
    wire N__12708;
    wire N__12705;
    wire N__12702;
    wire N__12699;
    wire N__12696;
    wire N__12693;
    wire N__12690;
    wire N__12687;
    wire N__12684;
    wire N__12681;
    wire N__12678;
    wire N__12675;
    wire N__12672;
    wire N__12671;
    wire N__12668;
    wire N__12665;
    wire N__12660;
    wire N__12659;
    wire N__12656;
    wire N__12653;
    wire N__12648;
    wire N__12645;
    wire N__12642;
    wire N__12639;
    wire N__12636;
    wire N__12633;
    wire N__12630;
    wire N__12627;
    wire N__12624;
    wire N__12621;
    wire N__12618;
    wire N__12615;
    wire N__12612;
    wire N__12609;
    wire N__12608;
    wire N__12605;
    wire N__12604;
    wire N__12601;
    wire N__12596;
    wire N__12593;
    wire N__12592;
    wire N__12589;
    wire N__12586;
    wire N__12583;
    wire N__12580;
    wire N__12573;
    wire N__12572;
    wire N__12567;
    wire N__12566;
    wire N__12563;
    wire N__12560;
    wire N__12557;
    wire N__12554;
    wire N__12549;
    wire N__12546;
    wire N__12543;
    wire N__12540;
    wire N__12539;
    wire N__12536;
    wire N__12533;
    wire N__12528;
    wire N__12525;
    wire N__12522;
    wire N__12519;
    wire N__12516;
    wire N__12513;
    wire N__12512;
    wire N__12509;
    wire N__12506;
    wire N__12501;
    wire N__12498;
    wire N__12495;
    wire N__12492;
    wire N__12491;
    wire N__12488;
    wire N__12485;
    wire N__12482;
    wire N__12479;
    wire N__12474;
    wire N__12471;
    wire N__12468;
    wire N__12465;
    wire N__12462;
    wire N__12459;
    wire N__12456;
    wire N__12453;
    wire N__12450;
    wire N__12449;
    wire N__12446;
    wire N__12443;
    wire N__12440;
    wire N__12435;
    wire N__12434;
    wire N__12431;
    wire N__12428;
    wire N__12425;
    wire N__12422;
    wire N__12417;
    wire N__12416;
    wire N__12413;
    wire N__12410;
    wire N__12407;
    wire N__12402;
    wire N__12401;
    wire N__12400;
    wire N__12397;
    wire N__12396;
    wire N__12393;
    wire N__12390;
    wire N__12389;
    wire N__12388;
    wire N__12375;
    wire N__12374;
    wire N__12371;
    wire N__12370;
    wire N__12369;
    wire N__12366;
    wire N__12363;
    wire N__12356;
    wire N__12351;
    wire N__12350;
    wire N__12349;
    wire N__12348;
    wire N__12347;
    wire N__12346;
    wire N__12333;
    wire N__12330;
    wire N__12329;
    wire N__12328;
    wire N__12325;
    wire N__12320;
    wire N__12315;
    wire N__12314;
    wire N__12313;
    wire N__12312;
    wire N__12311;
    wire N__12308;
    wire N__12305;
    wire N__12302;
    wire N__12301;
    wire N__12296;
    wire N__12289;
    wire N__12286;
    wire N__12283;
    wire N__12276;
    wire N__12273;
    wire N__12272;
    wire N__12271;
    wire N__12268;
    wire N__12265;
    wire N__12264;
    wire N__12263;
    wire N__12260;
    wire N__12255;
    wire N__12250;
    wire N__12243;
    wire N__12242;
    wire N__12241;
    wire N__12240;
    wire N__12239;
    wire N__12238;
    wire N__12235;
    wire N__12232;
    wire N__12229;
    wire N__12226;
    wire N__12221;
    wire N__12214;
    wire N__12207;
    wire N__12204;
    wire N__12203;
    wire N__12200;
    wire N__12197;
    wire N__12194;
    wire N__12191;
    wire N__12186;
    wire N__12183;
    wire N__12180;
    wire N__12179;
    wire N__12174;
    wire N__12171;
    wire N__12170;
    wire N__12169;
    wire N__12168;
    wire N__12167;
    wire N__12166;
    wire N__12165;
    wire N__12164;
    wire N__12161;
    wire N__12158;
    wire N__12145;
    wire N__12138;
    wire N__12135;
    wire N__12132;
    wire N__12129;
    wire N__12126;
    wire N__12123;
    wire N__12120;
    wire N__12117;
    wire N__12114;
    wire N__12111;
    wire N__12108;
    wire N__12105;
    wire N__12102;
    wire N__12099;
    wire N__12096;
    wire N__12093;
    wire N__12090;
    wire N__12087;
    wire N__12084;
    wire N__12083;
    wire N__12080;
    wire N__12077;
    wire N__12074;
    wire N__12071;
    wire N__12068;
    wire N__12065;
    wire N__12060;
    wire N__12057;
    wire N__12054;
    wire N__12051;
    wire N__12048;
    wire N__12045;
    wire N__12042;
    wire N__12039;
    wire N__12036;
    wire N__12033;
    wire N__12030;
    wire N__12027;
    wire N__12026;
    wire N__12023;
    wire N__12020;
    wire N__12017;
    wire N__12012;
    wire N__12011;
    wire N__12008;
    wire N__12005;
    wire N__12002;
    wire N__11997;
    wire N__11994;
    wire N__11993;
    wire N__11990;
    wire N__11987;
    wire N__11984;
    wire N__11981;
    wire N__11978;
    wire N__11975;
    wire N__11972;
    wire N__11969;
    wire N__11964;
    wire N__11963;
    wire N__11960;
    wire N__11957;
    wire N__11954;
    wire N__11949;
    wire N__11948;
    wire N__11945;
    wire N__11942;
    wire N__11937;
    wire N__11936;
    wire N__11933;
    wire N__11930;
    wire N__11925;
    wire N__11922;
    wire N__11919;
    wire N__11916;
    wire N__11913;
    wire N__11910;
    wire N__11907;
    wire N__11904;
    wire N__11901;
    wire N__11898;
    wire N__11895;
    wire N__11892;
    wire N__11889;
    wire N__11886;
    wire N__11883;
    wire N__11880;
    wire N__11877;
    wire N__11874;
    wire N__11871;
    wire N__11868;
    wire N__11865;
    wire N__11862;
    wire N__11859;
    wire N__11856;
    wire N__11853;
    wire N__11852;
    wire N__11849;
    wire N__11848;
    wire N__11845;
    wire N__11842;
    wire N__11839;
    wire N__11838;
    wire N__11835;
    wire N__11834;
    wire N__11829;
    wire N__11826;
    wire N__11823;
    wire N__11820;
    wire N__11815;
    wire N__11812;
    wire N__11809;
    wire N__11806;
    wire N__11799;
    wire N__11796;
    wire N__11793;
    wire N__11790;
    wire N__11787;
    wire N__11784;
    wire N__11781;
    wire N__11778;
    wire N__11775;
    wire N__11772;
    wire N__11769;
    wire N__11766;
    wire N__11763;
    wire N__11760;
    wire N__11757;
    wire N__11754;
    wire N__11751;
    wire N__11748;
    wire N__11745;
    wire N__11744;
    wire N__11743;
    wire N__11742;
    wire N__11741;
    wire N__11740;
    wire N__11739;
    wire N__11732;
    wire N__11731;
    wire N__11730;
    wire N__11729;
    wire N__11728;
    wire N__11727;
    wire N__11726;
    wire N__11723;
    wire N__11716;
    wire N__11713;
    wire N__11708;
    wire N__11699;
    wire N__11688;
    wire N__11685;
    wire N__11682;
    wire N__11679;
    wire N__11678;
    wire N__11677;
    wire N__11676;
    wire N__11675;
    wire N__11674;
    wire N__11673;
    wire N__11670;
    wire N__11667;
    wire N__11666;
    wire N__11665;
    wire N__11664;
    wire N__11663;
    wire N__11662;
    wire N__11659;
    wire N__11658;
    wire N__11657;
    wire N__11656;
    wire N__11655;
    wire N__11654;
    wire N__11651;
    wire N__11638;
    wire N__11637;
    wire N__11636;
    wire N__11635;
    wire N__11632;
    wire N__11619;
    wire N__11610;
    wire N__11607;
    wire N__11598;
    wire N__11589;
    wire N__11586;
    wire N__11583;
    wire N__11580;
    wire N__11577;
    wire N__11574;
    wire N__11573;
    wire N__11572;
    wire N__11569;
    wire N__11568;
    wire N__11565;
    wire N__11564;
    wire N__11563;
    wire N__11562;
    wire N__11559;
    wire N__11552;
    wire N__11549;
    wire N__11548;
    wire N__11547;
    wire N__11546;
    wire N__11545;
    wire N__11544;
    wire N__11539;
    wire N__11536;
    wire N__11533;
    wire N__11530;
    wire N__11523;
    wire N__11520;
    wire N__11517;
    wire N__11510;
    wire N__11499;
    wire N__11498;
    wire N__11497;
    wire N__11494;
    wire N__11493;
    wire N__11492;
    wire N__11491;
    wire N__11490;
    wire N__11489;
    wire N__11488;
    wire N__11487;
    wire N__11484;
    wire N__11481;
    wire N__11480;
    wire N__11475;
    wire N__11468;
    wire N__11467;
    wire N__11462;
    wire N__11459;
    wire N__11456;
    wire N__11455;
    wire N__11452;
    wire N__11449;
    wire N__11444;
    wire N__11441;
    wire N__11438;
    wire N__11435;
    wire N__11432;
    wire N__11429;
    wire N__11426;
    wire N__11421;
    wire N__11418;
    wire N__11415;
    wire N__11400;
    wire N__11399;
    wire N__11398;
    wire N__11397;
    wire N__11394;
    wire N__11393;
    wire N__11392;
    wire N__11389;
    wire N__11384;
    wire N__11381;
    wire N__11380;
    wire N__11379;
    wire N__11378;
    wire N__11377;
    wire N__11374;
    wire N__11371;
    wire N__11368;
    wire N__11363;
    wire N__11356;
    wire N__11353;
    wire N__11350;
    wire N__11337;
    wire N__11336;
    wire N__11333;
    wire N__11332;
    wire N__11329;
    wire N__11326;
    wire N__11323;
    wire N__11322;
    wire N__11321;
    wire N__11318;
    wire N__11313;
    wire N__11308;
    wire N__11301;
    wire N__11298;
    wire N__11295;
    wire N__11292;
    wire N__11289;
    wire N__11286;
    wire N__11285;
    wire N__11282;
    wire N__11279;
    wire N__11276;
    wire N__11271;
    wire N__11268;
    wire N__11265;
    wire N__11264;
    wire N__11263;
    wire N__11262;
    wire N__11261;
    wire N__11258;
    wire N__11257;
    wire N__11256;
    wire N__11251;
    wire N__11246;
    wire N__11245;
    wire N__11244;
    wire N__11241;
    wire N__11238;
    wire N__11235;
    wire N__11230;
    wire N__11225;
    wire N__11224;
    wire N__11221;
    wire N__11220;
    wire N__11219;
    wire N__11218;
    wire N__11213;
    wire N__11208;
    wire N__11205;
    wire N__11202;
    wire N__11197;
    wire N__11194;
    wire N__11189;
    wire N__11186;
    wire N__11175;
    wire N__11174;
    wire N__11173;
    wire N__11170;
    wire N__11167;
    wire N__11164;
    wire N__11157;
    wire N__11156;
    wire N__11155;
    wire N__11154;
    wire N__11153;
    wire N__11150;
    wire N__11149;
    wire N__11146;
    wire N__11141;
    wire N__11140;
    wire N__11139;
    wire N__11136;
    wire N__11133;
    wire N__11128;
    wire N__11125;
    wire N__11120;
    wire N__11119;
    wire N__11118;
    wire N__11117;
    wire N__11116;
    wire N__11109;
    wire N__11104;
    wire N__11095;
    wire N__11092;
    wire N__11085;
    wire N__11082;
    wire N__11079;
    wire N__11076;
    wire N__11073;
    wire N__11070;
    wire N__11067;
    wire N__11064;
    wire N__11061;
    wire N__11058;
    wire N__11055;
    wire N__11052;
    wire N__11049;
    wire N__11048;
    wire N__11043;
    wire N__11040;
    wire N__11039;
    wire N__11036;
    wire N__11035;
    wire N__11032;
    wire N__11029;
    wire N__11026;
    wire N__11023;
    wire N__11016;
    wire N__11015;
    wire N__11014;
    wire N__11013;
    wire N__11012;
    wire N__11011;
    wire N__11010;
    wire N__11009;
    wire N__11006;
    wire N__11005;
    wire N__11004;
    wire N__11001;
    wire N__10998;
    wire N__10997;
    wire N__10996;
    wire N__10995;
    wire N__10994;
    wire N__10993;
    wire N__10990;
    wire N__10985;
    wire N__10976;
    wire N__10961;
    wire N__10960;
    wire N__10959;
    wire N__10956;
    wire N__10955;
    wire N__10954;
    wire N__10953;
    wire N__10952;
    wire N__10949;
    wire N__10946;
    wire N__10941;
    wire N__10928;
    wire N__10927;
    wire N__10926;
    wire N__10925;
    wire N__10922;
    wire N__10919;
    wire N__10916;
    wire N__10913;
    wire N__10910;
    wire N__10903;
    wire N__10890;
    wire N__10889;
    wire N__10886;
    wire N__10883;
    wire N__10880;
    wire N__10879;
    wire N__10878;
    wire N__10877;
    wire N__10876;
    wire N__10873;
    wire N__10870;
    wire N__10865;
    wire N__10860;
    wire N__10851;
    wire N__10848;
    wire N__10845;
    wire N__10842;
    wire N__10839;
    wire N__10836;
    wire N__10833;
    wire N__10830;
    wire N__10827;
    wire N__10824;
    wire N__10823;
    wire N__10822;
    wire N__10821;
    wire N__10818;
    wire N__10815;
    wire N__10814;
    wire N__10813;
    wire N__10812;
    wire N__10809;
    wire N__10806;
    wire N__10803;
    wire N__10800;
    wire N__10795;
    wire N__10792;
    wire N__10791;
    wire N__10788;
    wire N__10787;
    wire N__10784;
    wire N__10779;
    wire N__10776;
    wire N__10773;
    wire N__10770;
    wire N__10767;
    wire N__10764;
    wire N__10759;
    wire N__10752;
    wire N__10749;
    wire N__10746;
    wire N__10743;
    wire N__10740;
    wire N__10735;
    wire N__10730;
    wire N__10727;
    wire N__10724;
    wire N__10721;
    wire N__10718;
    wire N__10713;
    wire N__10710;
    wire N__10709;
    wire N__10708;
    wire N__10707;
    wire N__10706;
    wire N__10703;
    wire N__10702;
    wire N__10701;
    wire N__10700;
    wire N__10699;
    wire N__10696;
    wire N__10695;
    wire N__10694;
    wire N__10693;
    wire N__10692;
    wire N__10687;
    wire N__10686;
    wire N__10685;
    wire N__10684;
    wire N__10683;
    wire N__10682;
    wire N__10679;
    wire N__10678;
    wire N__10677;
    wire N__10676;
    wire N__10675;
    wire N__10672;
    wire N__10667;
    wire N__10664;
    wire N__10659;
    wire N__10656;
    wire N__10653;
    wire N__10648;
    wire N__10645;
    wire N__10642;
    wire N__10637;
    wire N__10632;
    wire N__10627;
    wire N__10622;
    wire N__10619;
    wire N__10608;
    wire N__10603;
    wire N__10600;
    wire N__10581;
    wire N__10578;
    wire N__10575;
    wire N__10572;
    wire N__10569;
    wire N__10568;
    wire N__10567;
    wire N__10566;
    wire N__10565;
    wire N__10564;
    wire N__10563;
    wire N__10562;
    wire N__10561;
    wire N__10560;
    wire N__10559;
    wire N__10558;
    wire N__10557;
    wire N__10556;
    wire N__10555;
    wire N__10552;
    wire N__10549;
    wire N__10548;
    wire N__10547;
    wire N__10544;
    wire N__10537;
    wire N__10536;
    wire N__10535;
    wire N__10532;
    wire N__10531;
    wire N__10528;
    wire N__10527;
    wire N__10526;
    wire N__10523;
    wire N__10520;
    wire N__10519;
    wire N__10518;
    wire N__10517;
    wire N__10514;
    wire N__10513;
    wire N__10510;
    wire N__10509;
    wire N__10506;
    wire N__10505;
    wire N__10504;
    wire N__10503;
    wire N__10502;
    wire N__10499;
    wire N__10494;
    wire N__10491;
    wire N__10488;
    wire N__10483;
    wire N__10482;
    wire N__10479;
    wire N__10474;
    wire N__10463;
    wire N__10456;
    wire N__10453;
    wire N__10450;
    wire N__10443;
    wire N__10430;
    wire N__10425;
    wire N__10424;
    wire N__10417;
    wire N__10414;
    wire N__10409;
    wire N__10406;
    wire N__10403;
    wire N__10400;
    wire N__10393;
    wire N__10390;
    wire N__10387;
    wire N__10384;
    wire N__10381;
    wire N__10376;
    wire N__10369;
    wire N__10360;
    wire N__10357;
    wire N__10354;
    wire N__10351;
    wire N__10348;
    wire N__10345;
    wire N__10338;
    wire N__10335;
    wire N__10332;
    wire N__10329;
    wire N__10326;
    wire N__10323;
    wire N__10320;
    wire N__10317;
    wire N__10314;
    wire N__10313;
    wire N__10310;
    wire N__10307;
    wire N__10302;
    wire N__10299;
    wire N__10296;
    wire N__10293;
    wire N__10292;
    wire N__10291;
    wire N__10290;
    wire N__10289;
    wire N__10286;
    wire N__10283;
    wire N__10278;
    wire N__10277;
    wire N__10276;
    wire N__10275;
    wire N__10274;
    wire N__10273;
    wire N__10272;
    wire N__10271;
    wire N__10268;
    wire N__10261;
    wire N__10258;
    wire N__10253;
    wire N__10246;
    wire N__10243;
    wire N__10230;
    wire N__10229;
    wire N__10228;
    wire N__10225;
    wire N__10222;
    wire N__10221;
    wire N__10220;
    wire N__10219;
    wire N__10218;
    wire N__10217;
    wire N__10216;
    wire N__10215;
    wire N__10214;
    wire N__10211;
    wire N__10206;
    wire N__10201;
    wire N__10198;
    wire N__10193;
    wire N__10190;
    wire N__10185;
    wire N__10170;
    wire N__10169;
    wire N__10168;
    wire N__10165;
    wire N__10164;
    wire N__10163;
    wire N__10160;
    wire N__10159;
    wire N__10158;
    wire N__10157;
    wire N__10154;
    wire N__10153;
    wire N__10152;
    wire N__10151;
    wire N__10148;
    wire N__10143;
    wire N__10142;
    wire N__10139;
    wire N__10136;
    wire N__10129;
    wire N__10122;
    wire N__10117;
    wire N__10114;
    wire N__10101;
    wire N__10100;
    wire N__10099;
    wire N__10098;
    wire N__10097;
    wire N__10094;
    wire N__10093;
    wire N__10090;
    wire N__10087;
    wire N__10082;
    wire N__10081;
    wire N__10080;
    wire N__10077;
    wire N__10072;
    wire N__10071;
    wire N__10066;
    wire N__10065;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10057;
    wire N__10052;
    wire N__10051;
    wire N__10050;
    wire N__10049;
    wire N__10046;
    wire N__10043;
    wire N__10038;
    wire N__10033;
    wire N__10030;
    wire N__10027;
    wire N__10022;
    wire N__10019;
    wire N__10002;
    wire N__10001;
    wire N__9998;
    wire N__9997;
    wire N__9996;
    wire N__9995;
    wire N__9992;
    wire N__9989;
    wire N__9986;
    wire N__9985;
    wire N__9984;
    wire N__9983;
    wire N__9982;
    wire N__9981;
    wire N__9978;
    wire N__9977;
    wire N__9974;
    wire N__9969;
    wire N__9966;
    wire N__9963;
    wire N__9958;
    wire N__9955;
    wire N__9948;
    wire N__9945;
    wire N__9940;
    wire N__9927;
    wire N__9926;
    wire N__9925;
    wire N__9922;
    wire N__9921;
    wire N__9920;
    wire N__9919;
    wire N__9914;
    wire N__9913;
    wire N__9910;
    wire N__9909;
    wire N__9908;
    wire N__9907;
    wire N__9904;
    wire N__9903;
    wire N__9900;
    wire N__9899;
    wire N__9896;
    wire N__9893;
    wire N__9890;
    wire N__9887;
    wire N__9884;
    wire N__9881;
    wire N__9878;
    wire N__9873;
    wire N__9868;
    wire N__9861;
    wire N__9846;
    wire N__9843;
    wire N__9840;
    wire N__9839;
    wire N__9838;
    wire N__9833;
    wire N__9830;
    wire N__9827;
    wire N__9822;
    wire N__9819;
    wire N__9816;
    wire N__9813;
    wire N__9810;
    wire N__9807;
    wire N__9804;
    wire N__9801;
    wire N__9798;
    wire N__9795;
    wire N__9792;
    wire N__9789;
    wire N__9786;
    wire N__9783;
    wire N__9780;
    wire N__9777;
    wire N__9774;
    wire N__9771;
    wire N__9768;
    wire N__9765;
    wire N__9764;
    wire N__9761;
    wire N__9758;
    wire N__9755;
    wire N__9754;
    wire N__9749;
    wire N__9746;
    wire N__9743;
    wire N__9740;
    wire N__9735;
    wire N__9732;
    wire N__9731;
    wire N__9730;
    wire N__9727;
    wire N__9724;
    wire N__9721;
    wire N__9714;
    wire N__9711;
    wire N__9708;
    wire N__9705;
    wire N__9704;
    wire N__9701;
    wire N__9698;
    wire N__9693;
    wire N__9690;
    wire N__9687;
    wire N__9684;
    wire N__9681;
    wire N__9678;
    wire N__9677;
    wire N__9676;
    wire N__9673;
    wire N__9670;
    wire N__9667;
    wire N__9660;
    wire N__9659;
    wire N__9654;
    wire N__9651;
    wire N__9648;
    wire N__9645;
    wire N__9642;
    wire N__9641;
    wire N__9640;
    wire N__9637;
    wire N__9634;
    wire N__9631;
    wire N__9624;
    wire N__9621;
    wire N__9618;
    wire N__9615;
    wire N__9612;
    wire N__9609;
    wire N__9606;
    wire N__9605;
    wire N__9602;
    wire N__9599;
    wire N__9594;
    wire N__9593;
    wire N__9592;
    wire N__9591;
    wire N__9590;
    wire N__9589;
    wire N__9588;
    wire N__9573;
    wire N__9570;
    wire N__9569;
    wire N__9566;
    wire N__9563;
    wire N__9560;
    wire N__9557;
    wire N__9556;
    wire N__9551;
    wire N__9548;
    wire N__9543;
    wire N__9540;
    wire N__9537;
    wire N__9534;
    wire N__9531;
    wire N__9528;
    wire N__9525;
    wire N__9522;
    wire N__9519;
    wire N__9516;
    wire N__9513;
    wire N__9512;
    wire N__9511;
    wire N__9508;
    wire N__9505;
    wire N__9502;
    wire N__9497;
    wire N__9496;
    wire N__9495;
    wire N__9492;
    wire N__9489;
    wire N__9484;
    wire N__9477;
    wire N__9476;
    wire N__9473;
    wire N__9470;
    wire N__9469;
    wire N__9464;
    wire N__9461;
    wire N__9458;
    wire N__9457;
    wire N__9456;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9442;
    wire N__9435;
    wire N__9434;
    wire N__9431;
    wire N__9430;
    wire N__9429;
    wire N__9426;
    wire N__9425;
    wire N__9422;
    wire N__9417;
    wire N__9416;
    wire N__9413;
    wire N__9412;
    wire N__9409;
    wire N__9408;
    wire N__9403;
    wire N__9400;
    wire N__9399;
    wire N__9398;
    wire N__9397;
    wire N__9394;
    wire N__9391;
    wire N__9388;
    wire N__9385;
    wire N__9382;
    wire N__9379;
    wire N__9374;
    wire N__9373;
    wire N__9372;
    wire N__9369;
    wire N__9366;
    wire N__9363;
    wire N__9360;
    wire N__9351;
    wire N__9346;
    wire N__9333;
    wire N__9332;
    wire N__9329;
    wire N__9326;
    wire N__9325;
    wire N__9320;
    wire N__9319;
    wire N__9318;
    wire N__9317;
    wire N__9314;
    wire N__9311;
    wire N__9304;
    wire N__9297;
    wire N__9294;
    wire N__9291;
    wire N__9290;
    wire N__9285;
    wire N__9282;
    wire N__9279;
    wire N__9276;
    wire N__9273;
    wire N__9270;
    wire N__9267;
    wire N__9264;
    wire N__9261;
    wire N__9258;
    wire N__9255;
    wire N__9252;
    wire N__9249;
    wire N__9246;
    wire N__9243;
    wire N__9240;
    wire N__9237;
    wire N__9234;
    wire N__9231;
    wire N__9228;
    wire N__9225;
    wire N__9222;
    wire N__9219;
    wire N__9216;
    wire N__9213;
    wire N__9210;
    wire N__9207;
    wire N__9204;
    wire N__9201;
    wire N__9198;
    wire N__9195;
    wire N__9194;
    wire N__9193;
    wire N__9192;
    wire N__9191;
    wire N__9190;
    wire N__9189;
    wire N__9188;
    wire N__9187;
    wire N__9186;
    wire N__9185;
    wire N__9184;
    wire N__9183;
    wire N__9182;
    wire N__9181;
    wire N__9180;
    wire N__9179;
    wire N__9178;
    wire N__9177;
    wire N__9174;
    wire N__9171;
    wire N__9168;
    wire N__9165;
    wire N__9162;
    wire N__9159;
    wire N__9156;
    wire N__9153;
    wire N__9150;
    wire N__9147;
    wire N__9144;
    wire N__9141;
    wire N__9138;
    wire N__9135;
    wire N__9132;
    wire N__9129;
    wire N__9128;
    wire N__9127;
    wire N__9126;
    wire N__9125;
    wire N__9124;
    wire N__9121;
    wire N__9116;
    wire N__9115;
    wire N__9114;
    wire N__9113;
    wire N__9110;
    wire N__9101;
    wire N__9094;
    wire N__9085;
    wire N__9076;
    wire N__9073;
    wire N__9070;
    wire N__9067;
    wire N__9064;
    wire N__9061;
    wire N__9060;
    wire N__9059;
    wire N__9058;
    wire N__9057;
    wire N__9056;
    wire N__9055;
    wire N__9054;
    wire N__9051;
    wire N__9048;
    wire N__9041;
    wire N__9034;
    wire N__9029;
    wire N__9024;
    wire N__9017;
    wire N__9014;
    wire N__9011;
    wire N__9008;
    wire N__9005;
    wire N__9002;
    wire N__8999;
    wire N__8996;
    wire N__8993;
    wire N__8990;
    wire N__8987;
    wire N__8978;
    wire N__8971;
    wire N__8962;
    wire N__8955;
    wire N__8948;
    wire N__8943;
    wire N__8940;
    wire N__8937;
    wire N__8934;
    wire N__8931;
    wire N__8928;
    wire N__8925;
    wire N__8922;
    wire N__8921;
    wire N__8916;
    wire N__8913;
    wire N__8910;
    wire N__8907;
    wire N__8906;
    wire N__8905;
    wire N__8902;
    wire N__8897;
    wire N__8894;
    wire N__8891;
    wire N__8888;
    wire N__8883;
    wire N__8880;
    wire N__8877;
    wire N__8874;
    wire N__8873;
    wire N__8870;
    wire N__8869;
    wire N__8868;
    wire N__8867;
    wire N__8866;
    wire N__8865;
    wire N__8864;
    wire N__8863;
    wire N__8860;
    wire N__8857;
    wire N__8854;
    wire N__8847;
    wire N__8840;
    wire N__8829;
    wire N__8826;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8816;
    wire N__8811;
    wire N__8808;
    wire N__8805;
    wire N__8802;
    wire N__8801;
    wire N__8800;
    wire N__8799;
    wire N__8798;
    wire N__8795;
    wire N__8792;
    wire N__8789;
    wire N__8788;
    wire N__8787;
    wire N__8786;
    wire N__8785;
    wire N__8784;
    wire N__8783;
    wire N__8780;
    wire N__8777;
    wire N__8770;
    wire N__8765;
    wire N__8762;
    wire N__8755;
    wire N__8742;
    wire N__8741;
    wire N__8740;
    wire N__8739;
    wire N__8732;
    wire N__8731;
    wire N__8730;
    wire N__8729;
    wire N__8726;
    wire N__8723;
    wire N__8714;
    wire N__8709;
    wire N__8708;
    wire N__8707;
    wire N__8704;
    wire N__8699;
    wire N__8694;
    wire N__8693;
    wire N__8692;
    wire N__8689;
    wire N__8688;
    wire N__8683;
    wire N__8680;
    wire N__8679;
    wire N__8678;
    wire N__8677;
    wire N__8676;
    wire N__8673;
    wire N__8668;
    wire N__8663;
    wire N__8656;
    wire N__8649;
    wire N__8648;
    wire N__8647;
    wire N__8640;
    wire N__8639;
    wire N__8638;
    wire N__8637;
    wire N__8634;
    wire N__8631;
    wire N__8626;
    wire N__8619;
    wire N__8616;
    wire N__8613;
    wire N__8610;
    wire N__8607;
    wire N__8604;
    wire N__8601;
    wire N__8598;
    wire N__8595;
    wire N__8592;
    wire N__8589;
    wire N__8586;
    wire N__8583;
    wire N__8580;
    wire N__8577;
    wire N__8574;
    wire N__8571;
    wire N__8568;
    wire N__8565;
    wire N__8562;
    wire N__8559;
    wire N__8556;
    wire N__8553;
    wire N__8550;
    wire N__8547;
    wire N__8544;
    wire N__8543;
    wire N__8540;
    wire N__8537;
    wire N__8536;
    wire N__8533;
    wire N__8530;
    wire N__8527;
    wire N__8524;
    wire N__8521;
    wire N__8514;
    wire N__8513;
    wire N__8510;
    wire N__8509;
    wire N__8506;
    wire N__8503;
    wire N__8500;
    wire N__8497;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8475;
    wire N__8472;
    wire N__8469;
    wire N__8466;
    wire N__8463;
    wire N__8462;
    wire N__8459;
    wire N__8458;
    wire N__8455;
    wire N__8452;
    wire N__8447;
    wire N__8442;
    wire N__8439;
    wire N__8436;
    wire N__8433;
    wire N__8430;
    wire N__8427;
    wire N__8424;
    wire N__8421;
    wire N__8418;
    wire N__8415;
    wire N__8412;
    wire N__8409;
    wire N__8406;
    wire N__8403;
    wire N__8400;
    wire N__8397;
    wire N__8394;
    wire N__8393;
    wire N__8392;
    wire N__8391;
    wire N__8390;
    wire N__8387;
    wire N__8386;
    wire N__8383;
    wire N__8382;
    wire N__8379;
    wire N__8376;
    wire N__8373;
    wire N__8370;
    wire N__8369;
    wire N__8366;
    wire N__8365;
    wire N__8364;
    wire N__8363;
    wire N__8362;
    wire N__8361;
    wire N__8358;
    wire N__8355;
    wire N__8352;
    wire N__8349;
    wire N__8344;
    wire N__8341;
    wire N__8334;
    wire N__8327;
    wire N__8310;
    wire N__8307;
    wire N__8304;
    wire N__8303;
    wire N__8302;
    wire N__8301;
    wire N__8300;
    wire N__8299;
    wire N__8298;
    wire N__8297;
    wire N__8294;
    wire N__8289;
    wire N__8286;
    wire N__8283;
    wire N__8280;
    wire N__8279;
    wire N__8278;
    wire N__8277;
    wire N__8274;
    wire N__8273;
    wire N__8272;
    wire N__8269;
    wire N__8268;
    wire N__8267;
    wire N__8266;
    wire N__8265;
    wire N__8264;
    wire N__8263;
    wire N__8262;
    wire N__8261;
    wire N__8260;
    wire N__8259;
    wire N__8256;
    wire N__8253;
    wire N__8252;
    wire N__8251;
    wire N__8250;
    wire N__8247;
    wire N__8244;
    wire N__8239;
    wire N__8236;
    wire N__8233;
    wire N__8228;
    wire N__8223;
    wire N__8218;
    wire N__8201;
    wire N__8196;
    wire N__8189;
    wire N__8182;
    wire N__8163;
    wire N__8160;
    wire N__8157;
    wire N__8156;
    wire N__8155;
    wire N__8152;
    wire N__8149;
    wire N__8146;
    wire N__8139;
    wire N__8136;
    wire N__8133;
    wire N__8130;
    wire N__8129;
    wire N__8128;
    wire N__8125;
    wire N__8120;
    wire N__8115;
    wire N__8112;
    wire N__8109;
    wire N__8106;
    wire N__8103;
    wire N__8102;
    wire N__8101;
    wire N__8098;
    wire N__8093;
    wire N__8088;
    wire N__8085;
    wire N__8082;
    wire N__8079;
    wire N__8076;
    wire N__8075;
    wire N__8074;
    wire N__8071;
    wire N__8066;
    wire N__8061;
    wire N__8058;
    wire N__8055;
    wire N__8052;
    wire N__8049;
    wire N__8048;
    wire N__8045;
    wire N__8042;
    wire N__8037;
    wire N__8034;
    wire N__8031;
    wire N__8028;
    wire N__8025;
    wire N__8022;
    wire N__8019;
    wire N__8016;
    wire N__8013;
    wire N__8010;
    wire N__8007;
    wire N__8004;
    wire N__8001;
    wire N__7998;
    wire N__7995;
    wire N__7992;
    wire N__7989;
    wire N__7986;
    wire N__7983;
    wire N__7980;
    wire N__7977;
    wire N__7974;
    wire N__7971;
    wire N__7970;
    wire N__7967;
    wire N__7964;
    wire N__7959;
    wire N__7958;
    wire N__7957;
    wire N__7950;
    wire N__7947;
    wire N__7944;
    wire N__7941;
    wire N__7938;
    wire N__7935;
    wire N__7932;
    wire N__7929;
    wire N__7926;
    wire N__7925;
    wire N__7924;
    wire N__7923;
    wire N__7918;
    wire N__7913;
    wire N__7908;
    wire N__7905;
    wire N__7902;
    wire N__7901;
    wire N__7900;
    wire N__7899;
    wire N__7898;
    wire N__7893;
    wire N__7886;
    wire N__7881;
    wire N__7880;
    wire N__7879;
    wire N__7878;
    wire N__7875;
    wire N__7872;
    wire N__7869;
    wire N__7868;
    wire N__7863;
    wire N__7856;
    wire N__7851;
    wire N__7848;
    wire N__7847;
    wire N__7846;
    wire N__7845;
    wire N__7840;
    wire N__7835;
    wire N__7830;
    wire N__7829;
    wire N__7828;
    wire N__7827;
    wire N__7826;
    wire N__7821;
    wire N__7814;
    wire N__7809;
    wire N__7806;
    wire N__7803;
    wire N__7800;
    wire N__7797;
    wire N__7794;
    wire N__7791;
    wire N__7790;
    wire N__7787;
    wire N__7784;
    wire N__7779;
    wire N__7778;
    wire N__7775;
    wire N__7772;
    wire N__7769;
    wire N__7768;
    wire N__7765;
    wire N__7762;
    wire N__7759;
    wire N__7758;
    wire N__7755;
    wire N__7752;
    wire N__7749;
    wire N__7746;
    wire N__7743;
    wire N__7734;
    wire N__7731;
    wire N__7728;
    wire N__7725;
    wire N__7722;
    wire N__7719;
    wire N__7716;
    wire N__7713;
    wire N__7710;
    wire N__7707;
    wire N__7704;
    wire N__7701;
    wire N__7698;
    wire N__7695;
    wire N__7692;
    wire N__7689;
    wire N__7686;
    wire N__7683;
    wire N__7680;
    wire N__7677;
    wire N__7674;
    wire N__7671;
    wire N__7668;
    wire N__7665;
    wire N__7664;
    wire N__7659;
    wire N__7656;
    wire N__7653;
    wire N__7650;
    wire N__7647;
    wire N__7644;
    wire N__7641;
    wire N__7638;
    wire N__7635;
    wire N__7632;
    wire N__7629;
    wire N__7626;
    wire N__7623;
    wire N__7620;
    wire N__7617;
    wire N__7614;
    wire N__7611;
    wire N__7608;
    wire N__7605;
    wire N__7602;
    wire N__7599;
    wire N__7596;
    wire N__7593;
    wire N__7590;
    wire N__7587;
    wire N__7584;
    wire N__7581;
    wire N__7578;
    wire N__7575;
    wire N__7572;
    wire N__7569;
    wire N__7566;
    wire N__7563;
    wire N__7560;
    wire N__7557;
    wire N__7554;
    wire N__7551;
    wire N__7548;
    wire N__7545;
    wire N__7542;
    wire N__7539;
    wire N__7538;
    wire N__7537;
    wire N__7534;
    wire N__7531;
    wire N__7528;
    wire N__7521;
    wire N__7518;
    wire N__7515;
    wire N__7512;
    wire N__7511;
    wire N__7510;
    wire N__7507;
    wire N__7504;
    wire N__7501;
    wire N__7494;
    wire N__7491;
    wire N__7488;
    wire N__7487;
    wire N__7484;
    wire N__7481;
    wire N__7476;
    wire N__7473;
    wire N__7470;
    wire N__7469;
    wire N__7466;
    wire N__7463;
    wire N__7458;
    wire N__7455;
    wire N__7452;
    wire N__7451;
    wire N__7450;
    wire N__7447;
    wire N__7444;
    wire N__7439;
    wire N__7434;
    wire N__7431;
    wire N__7428;
    wire N__7427;
    wire N__7426;
    wire N__7423;
    wire N__7420;
    wire N__7417;
    wire N__7414;
    wire N__7407;
    wire N__7404;
    wire N__7401;
    wire N__7398;
    wire N__7397;
    wire N__7394;
    wire N__7391;
    wire N__7386;
    wire N__7383;
    wire N__7380;
    wire N__7377;
    wire N__7374;
    wire N__7371;
    wire N__7368;
    wire N__7367;
    wire N__7366;
    wire N__7365;
    wire N__7364;
    wire N__7363;
    wire N__7358;
    wire N__7351;
    wire N__7348;
    wire N__7345;
    wire N__7342;
    wire N__7335;
    wire N__7332;
    wire N__7331;
    wire N__7328;
    wire N__7325;
    wire N__7322;
    wire N__7321;
    wire N__7320;
    wire N__7319;
    wire N__7318;
    wire N__7317;
    wire N__7314;
    wire N__7311;
    wire N__7308;
    wire N__7303;
    wire N__7298;
    wire N__7287;
    wire N__7286;
    wire N__7283;
    wire N__7280;
    wire N__7277;
    wire N__7274;
    wire N__7271;
    wire N__7266;
    wire N__7263;
    wire N__7260;
    wire N__7259;
    wire N__7258;
    wire N__7255;
    wire N__7252;
    wire N__7249;
    wire N__7242;
    wire N__7239;
    wire N__7236;
    wire N__7233;
    wire N__7232;
    wire N__7231;
    wire N__7228;
    wire N__7225;
    wire N__7222;
    wire N__7215;
    wire N__7212;
    wire N__7209;
    wire N__7208;
    wire N__7207;
    wire N__7204;
    wire N__7199;
    wire N__7194;
    wire N__7191;
    wire N__7188;
    wire N__7185;
    wire N__7184;
    wire N__7183;
    wire N__7180;
    wire N__7175;
    wire N__7170;
    wire N__7167;
    wire N__7164;
    wire N__7161;
    wire N__7160;
    wire N__7159;
    wire N__7156;
    wire N__7151;
    wire N__7146;
    wire N__7143;
    wire N__7142;
    wire N__7141;
    wire N__7138;
    wire N__7133;
    wire N__7128;
    wire N__7127;
    wire N__7126;
    wire N__7125;
    wire N__7124;
    wire N__7123;
    wire N__7122;
    wire N__7121;
    wire N__7120;
    wire N__7115;
    wire N__7110;
    wire N__7105;
    wire N__7098;
    wire N__7095;
    wire N__7088;
    wire N__7083;
    wire N__7082;
    wire N__7081;
    wire N__7080;
    wire N__7077;
    wire N__7076;
    wire N__7073;
    wire N__7072;
    wire N__7071;
    wire N__7070;
    wire N__7069;
    wire N__7066;
    wire N__7061;
    wire N__7058;
    wire N__7055;
    wire N__7048;
    wire N__7043;
    wire N__7032;
    wire N__7029;
    wire N__7028;
    wire N__7025;
    wire N__7022;
    wire N__7017;
    wire N__7014;
    wire N__7013;
    wire N__7012;
    wire N__7011;
    wire N__7010;
    wire N__7009;
    wire N__7008;
    wire N__7005;
    wire N__7002;
    wire N__7001;
    wire N__7000;
    wire N__6999;
    wire N__6998;
    wire N__6989;
    wire N__6986;
    wire N__6983;
    wire N__6980;
    wire N__6971;
    wire N__6960;
    wire N__6959;
    wire N__6958;
    wire N__6951;
    wire N__6948;
    wire N__6945;
    wire N__6942;
    wire N__6939;
    wire N__6938;
    wire N__6935;
    wire N__6934;
    wire N__6933;
    wire N__6928;
    wire N__6923;
    wire N__6918;
    wire N__6915;
    wire N__6912;
    wire N__6911;
    wire N__6910;
    wire N__6909;
    wire N__6908;
    wire N__6905;
    wire N__6900;
    wire N__6895;
    wire N__6888;
    wire N__6885;
    wire N__6882;
    wire N__6881;
    wire N__6880;
    wire N__6879;
    wire N__6878;
    wire N__6875;
    wire N__6870;
    wire N__6867;
    wire N__6864;
    wire N__6859;
    wire N__6852;
    wire N__6849;
    wire N__6846;
    wire N__6843;
    wire N__6842;
    wire N__6839;
    wire N__6838;
    wire N__6837;
    wire N__6836;
    wire N__6835;
    wire N__6832;
    wire N__6829;
    wire N__6824;
    wire N__6819;
    wire N__6810;
    wire N__6807;
    wire N__6806;
    wire N__6805;
    wire N__6802;
    wire N__6797;
    wire N__6792;
    wire N__6791;
    wire N__6790;
    wire N__6789;
    wire N__6788;
    wire N__6785;
    wire N__6784;
    wire N__6781;
    wire N__6780;
    wire N__6779;
    wire N__6778;
    wire N__6775;
    wire N__6772;
    wire N__6769;
    wire N__6766;
    wire N__6759;
    wire N__6750;
    wire N__6741;
    wire N__6740;
    wire N__6737;
    wire N__6734;
    wire N__6733;
    wire N__6732;
    wire N__6731;
    wire N__6730;
    wire N__6729;
    wire N__6728;
    wire N__6725;
    wire N__6722;
    wire N__6713;
    wire N__6708;
    wire N__6699;
    wire N__6696;
    wire N__6695;
    wire N__6694;
    wire N__6693;
    wire N__6688;
    wire N__6683;
    wire N__6678;
    wire N__6675;
    wire N__6672;
    wire N__6671;
    wire N__6670;
    wire N__6669;
    wire N__6666;
    wire N__6665;
    wire N__6662;
    wire N__6657;
    wire N__6654;
    wire N__6651;
    wire N__6648;
    wire N__6645;
    wire N__6636;
    wire N__6633;
    wire N__6630;
    wire N__6629;
    wire N__6626;
    wire N__6623;
    wire N__6618;
    wire N__6615;
    wire N__6612;
    wire N__6609;
    wire N__6606;
    wire N__6605;
    wire N__6602;
    wire N__6599;
    wire N__6594;
    wire N__6591;
    wire N__6588;
    wire N__6585;
    wire N__6584;
    wire N__6581;
    wire N__6580;
    wire N__6577;
    wire N__6574;
    wire N__6571;
    wire N__6564;
    wire N__6561;
    wire N__6558;
    wire N__6555;
    wire N__6554;
    wire N__6551;
    wire N__6548;
    wire N__6543;
    wire N__6540;
    wire N__6539;
    wire N__6536;
    wire N__6533;
    wire N__6530;
    wire N__6525;
    wire N__6522;
    wire N__6521;
    wire N__6518;
    wire N__6515;
    wire N__6510;
    wire N__6507;
    wire N__6504;
    wire N__6503;
    wire N__6500;
    wire N__6497;
    wire N__6494;
    wire N__6489;
    wire N__6486;
    wire N__6485;
    wire N__6484;
    wire N__6483;
    wire N__6480;
    wire N__6473;
    wire N__6468;
    wire N__6465;
    wire N__6464;
    wire N__6461;
    wire N__6460;
    wire N__6459;
    wire N__6458;
    wire N__6455;
    wire N__6452;
    wire N__6445;
    wire N__6438;
    wire N__6435;
    wire N__6432;
    wire N__6429;
    wire N__6428;
    wire N__6427;
    wire N__6426;
    wire N__6423;
    wire N__6422;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire N__6412;
    wire N__6409;
    wire N__6400;
    wire N__6393;
    wire N__6390;
    wire N__6387;
    wire N__6386;
    wire N__6383;
    wire N__6380;
    wire N__6375;
    wire N__6372;
    wire N__6371;
    wire N__6368;
    wire N__6365;
    wire N__6362;
    wire N__6357;
    wire N__6354;
    wire N__6353;
    wire N__6350;
    wire N__6347;
    wire N__6344;
    wire N__6339;
    wire N__6336;
    wire N__6335;
    wire N__6332;
    wire N__6329;
    wire N__6324;
    wire N__6321;
    wire N__6320;
    wire N__6317;
    wire N__6314;
    wire N__6309;
    wire N__6306;
    wire N__6305;
    wire N__6302;
    wire N__6299;
    wire N__6294;
    wire N__6291;
    wire N__6290;
    wire N__6287;
    wire N__6284;
    wire N__6279;
    wire N__6276;
    wire N__6275;
    wire N__6272;
    wire N__6269;
    wire N__6264;
    wire N__6261;
    wire N__6260;
    wire N__6257;
    wire N__6254;
    wire N__6249;
    wire N__6246;
    wire N__6245;
    wire N__6242;
    wire N__6239;
    wire N__6234;
    wire N__6231;
    wire N__6228;
    wire N__6225;
    wire N__6222;
    wire N__6219;
    wire N__6216;
    wire N__6213;
    wire N__6210;
    wire N__6207;
    wire N__6204;
    wire N__6201;
    wire N__6198;
    wire N__6195;
    wire N__6192;
    wire N__6189;
    wire N__6188;
    wire N__6187;
    wire N__6184;
    wire N__6179;
    wire N__6174;
    wire N__6173;
    wire N__6170;
    wire N__6167;
    wire N__6166;
    wire N__6159;
    wire N__6156;
    wire N__6153;
    wire N__6150;
    wire N__6147;
    wire N__6144;
    wire N__6141;
    wire N__6138;
    wire N__6135;
    wire N__6132;
    wire N__6129;
    wire N__6126;
    wire N__6123;
    wire N__6120;
    wire N__6117;
    wire N__6114;
    wire N__6111;
    wire N__6108;
    wire N__6105;
    wire N__6102;
    wire N__6099;
    wire N__6096;
    wire N__6093;
    wire N__6090;
    wire N__6087;
    wire N__6084;
    wire N__6081;
    wire N__6078;
    wire N__6075;
    wire N__6072;
    wire N__6069;
    wire N__6066;
    wire N__6063;
    wire N__6060;
    wire N__6057;
    wire N__6054;
    wire N__6051;
    wire N__6048;
    wire N__6045;
    wire N__6042;
    wire N__6039;
    wire N__6036;
    wire N__6033;
    wire N__6030;
    wire N__6027;
    wire N__6024;
    wire N__6021;
    wire N__6018;
    wire N__6015;
    wire N__6014;
    wire N__6009;
    wire N__6006;
    wire N__6003;
    wire N__6000;
    wire N__5997;
    wire N__5994;
    wire N__5991;
    wire N__5988;
    wire N__5985;
    wire N__5982;
    wire N__5979;
    wire N__5976;
    wire N__5973;
    wire N__5970;
    wire N__5967;
    wire N__5964;
    wire N__5961;
    wire N__5958;
    wire N__5955;
    wire N__5952;
    wire N__5949;
    wire N__5946;
    wire N__5943;
    wire N__5940;
    wire N__5937;
    wire N__5934;
    wire N__5931;
    wire N__5928;
    wire N__5925;
    wire N__5922;
    wire N__5919;
    wire N__5916;
    wire N__5913;
    wire N__5910;
    wire N__5907;
    wire N__5904;
    wire N__5901;
    wire N__5898;
    wire N__5895;
    wire N__5892;
    wire N__5889;
    wire N__5886;
    wire N__5883;
    wire N__5880;
    wire N__5877;
    wire N__5874;
    wire N__5871;
    wire N__5868;
    wire N__5865;
    wire N__5862;
    wire wRamRdData_1;
    wire wRamRdData_6;
    wire wRamRdData_2;
    wire wRamRdData_5;
    wire wRamRdData_4;
    wire BTN_N_c;
    wire wRamRdData_7;
    wire wRamRdData_0;
    wire VCCG0;
    wire wRamRdData_3;
    wire GNDG0;
    wire \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO ;
    wire \top_pll_inst.wPllLocked_iso_i ;
    wire \DUT.uart_inst0.N_6_0_cascade_ ;
    wire \DUT.uart_inst0.N_22_cascade_ ;
    wire \DUT.uart_inst0.N_22 ;
    wire \DUT.uart_inst0.g2_3_cascade_ ;
    wire \DUT.uart_inst0.g2 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_9 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_8 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_6_cascade_ ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_7 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_0_cascade_ ;
    wire \DUT.uart_inst0.N_152_cascade_ ;
    wire \DUT.uart_inst0.N_5 ;
    wire \DUT.uart_inst0.tx_countdown_7_m1_0_o2_2_2_cascade_ ;
    wire \DUT.uart_inst0.tx_out_6_iv_0_a3_0_1_cascade_ ;
    wire \DUT.uart_inst0.tx_out_6_iv_0_1_cascade_ ;
    wire \DUT.uart_inst0.N_119 ;
    wire \DUT.uart_inst0.tx_countdown_RNO_0Z0Z_4_cascade_ ;
    wire \DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0_cascade_ ;
    wire \DUT.uart_inst0.m25_e_3_cascade_ ;
    wire \DUT.uart_inst0.m3_0 ;
    wire bfn_13_7_0_;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_0 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_1 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_2 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_3 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_4 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_5 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_6 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_7 ;
    wire bfn_13_8_0_;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_8 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_9 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_10 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_11 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_12 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_13 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_14 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_15 ;
    wire bfn_13_9_0_;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_16 ;
    wire bfn_13_10_0_;
    wire \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0 ;
    wire \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1 ;
    wire \DUT.fifo_tx_inst.rFifoCount_RNISSQ21Z0Z_1 ;
    wire \DUT.fifo_tx_inst.N_108_cascade_ ;
    wire \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0 ;
    wire \DUT.fifo_tx_inst.N_108 ;
    wire rTxWriteZ0;
    wire \DUT.fifo_tx_inst.N_104_cascade_ ;
    wire \DUT.uart_inst0.rx_countdown_8_i_o2_1_2_cascade_ ;
    wire \DUT.uart_inst0.N_67 ;
    wire \DUT.uart_inst0.g0_0_0_a3_0_3_cascade_ ;
    wire \DUT.uart_inst0.N_159_0 ;
    wire \DUT.uart_inst0.N_4 ;
    wire bfn_14_2_0_;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_1 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_0 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_2 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_1 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_3 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_2 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_4 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_3 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_5 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_4 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_6 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_5 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_7 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_6 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_7 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_8 ;
    wire bfn_14_3_0_;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_9 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_8 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_10 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_9 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_11 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_10 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_12 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_11 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_12 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_13 ;
    wire \DUT.uart_inst0.tx_bits_remainingZ0Z_2 ;
    wire \DUT.uart_inst0.tx_bits_remainingZ0Z_1 ;
    wire \DUT.uart_inst0.m9_e_0_3 ;
    wire \DUT.uart_inst0.tx_bits_remainingZ0Z_0 ;
    wire \DUT.uart_inst0.m9_e_0_0 ;
    wire \DUT.uart_inst0.N_152 ;
    wire \DUT.uart_inst0.tx_state_0_sqmuxa_i_i_a3_c_cascade_ ;
    wire \DUT.uart_inst0.N_160_cascade_ ;
    wire \DUT.uart_inst0.tx_countdown_0_ac0_1 ;
    wire \DUT.uart_inst0.N_154 ;
    wire \DUT.uart_inst0.tx_bits_remainingZ0Z_3 ;
    wire \DUT.uart_inst0.N_72 ;
    wire \DUT.uart_inst0.N_99 ;
    wire \DUT.uart_inst0.tx_countdown_RNO_0Z0Z_1 ;
    wire \DUT.uart_inst0.N_88_i ;
    wire \DUT.uart_inst0.N_160 ;
    wire \DUT.uart_inst0.N_218 ;
    wire \DUT.uart_inst0.N_218_cascade_ ;
    wire \DUT.uart_inst0.N_109 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_1 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_0 ;
    wire \DUT.uart_inst0.N_120 ;
    wire \DUT.uart_inst0.tx_countdown_RNO_1Z0Z_3_cascade_ ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_0 ;
    wire \DUT.uart_inst0.N_164 ;
    wire \DUT.uart_inst0.N_164_cascade_ ;
    wire \DUT.uart_inst0.tx_countdown_RNO_0Z0Z_3 ;
    wire \DUT.uart_inst0.tx_state_ns_i_i_o2_a0_2_0 ;
    wire \DUT.uart_inst0.N_159 ;
    wire \DUT.uart_inst0.N_100 ;
    wire \DUT.uart_inst0.N_163 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_5 ;
    wire \DUT.uart_inst0.tx_countdown_0_c3 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_3 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_4 ;
    wire \DUT.uart_inst0.tx_countdown_30_5 ;
    wire \DUT.uart_inst0.tx_countdown_7_m1_0_a3_0_2 ;
    wire \DUT.uart_inst0.N_113 ;
    wire \DUT.uart_inst0.tx_countdown_7_sm0_0 ;
    wire \DUT.uart_inst0.N_84 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_17 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_13 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_14 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_15 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_10 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_9 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_11 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_7 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_5 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_5 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_6 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_6 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_8 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_12 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO ;
    wire \DUT.uart_inst0.m7_e_1_cascade_ ;
    wire \DUT.uart_inst0.m7_e_3_cascade_ ;
    wire \DUT.uart_inst0.m9_1_cascade_ ;
    wire \DUT.uart_inst0.N_11_mux ;
    wire \DUT.uart_inst0.N_66 ;
    wire \DUT.uart_inst0.m4_e_0 ;
    wire \DUT.uart_inst0.m4_e_3 ;
    wire \DUT.uart_inst0.N_21_0_cascade_ ;
    wire \DUT.uart_inst0.N_21_mux_0 ;
    wire \DUT.uart_inst0.m5_1 ;
    wire \DUT.uart_inst0.N_6 ;
    wire \DUT.uart_inst0.N_6_cascade_ ;
    wire \DUT.uart_inst0.N_18 ;
    wire \DUT.uart_inst0.N_18_mux_0 ;
    wire \DUT.uart_inst0.N_30 ;
    wire \DUT.uart_inst0.g1_i_a4_0_4 ;
    wire \DUT.uart_inst0.g1_i_a4_0_5_cascade_ ;
    wire \DUT.uart_inst0.g0_0_0_a3_0_4 ;
    wire \DUT.uart_inst0.g0_0_0_a3_4_cascade_ ;
    wire \DUT.uart_inst0.g0_0_0_a3_3 ;
    wire \DUT.fifo_tx_inst.un1_i11_i_cascade_ ;
    wire \DUT.fifo_rx_inst.N_57_cascade_ ;
    wire \DUT.fifo_rx_inst.un1_i11_i ;
    wire \DUT.uart_inst0.m13_2_cascade_ ;
    wire \DUT.uart_inst0.m13_3 ;
    wire \DUT.uart_inst0.P19_mux_cascade_ ;
    wire \DUT.uart_inst0.g0_0_1 ;
    wire N_1257_i;
    wire G_111_cascade_;
    wire \fifo_inst.ftdi_input_inst.SUMZ0Z_2_cascade_ ;
    wire G_110_cascade_;
    wire fifo_inst_ftdi_input_inst_oTxFull_0;
    wire G_108;
    wire \fifo_inst.ftdi_input_inst.SUMZ0Z_3 ;
    wire G_109;
    wire G_110;
    wire G_111;
    wire G_112;
    wire \fifo_inst.ftdi_input_inst.un2_oPacketAvail_iZ0 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_0 ;
    wire P1A7_c;
    wire \DUT.uart_inst0.N_116 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_1 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_2 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_3 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_4 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_5 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_7 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_6 ;
    wire \DUT.uart_inst0.N_22_i ;
    wire \DUT.uart_inst0.N_102 ;
    wire \DUT.uart_inst0.tx_state_0_sqmuxa_i_i_a3_0_1 ;
    wire \DUT.tx_state_1 ;
    wire \DUT.N_114_cascade_ ;
    wire \DUT.tx_state_0 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_16 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_9_cascade_ ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_1 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_dividerZ1Z_1 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_2 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_3 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_3 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_4 ;
    wire \DUT.uart_inst0.m6_3_cascade_ ;
    wire \top_pll_inst.m12_1_1_cascade_ ;
    wire \DUT.uart_inst0.G_30_1 ;
    wire P18_mux_cascade_;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_11 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_10 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_12 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_13 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_0_cascade_ ;
    wire bfn_15_9_0_;
    wire \DUT.uart_inst0.rx_countdown_3_cry_0_s1 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_1_s1 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_2_s1 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_3_s1 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_4_s1 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_0 ;
    wire \DUT.uart_inst0.N_20 ;
    wire \DUT.uart_inst0.N_21_cascade_ ;
    wire \DUT.uart_inst0.N_21_mux_cascade_ ;
    wire \DUT.uart_inst0.N_19_mux ;
    wire \DUT.uart_inst0.N_13_cascade_ ;
    wire \DUT.uart_inst0.N_13_0 ;
    wire \DUT.uart_inst0.rx_countdown_8_i_o2_2_0_2_cascade_ ;
    wire \DUT.fifo_tx_inst.un1_i11_i ;
    wire \DUT.uart_inst0.g0_0 ;
    wire \DUT.uart_inst0.N_49 ;
    wire \DUT.uart_inst0.m6_1 ;
    wire \DUT.uart_inst0.N_7 ;
    wire \DUT.uart_inst0.recv_state_srsts_1_5 ;
    wire \DUT.uart_inst0.rx_countdown_8_i_o2_2_2 ;
    wire \DUT.uart_inst0.recv_state_srsts_1_5_cascade_ ;
    wire \DUT.uart_inst0.recv_state_srsts_1_4 ;
    wire \DUT.uart_inst0.recv_stateZ0Z_1 ;
    wire \DUT.uart_inst0.N_43_cascade_ ;
    wire \DUT.uart_inst0.recv_state_RNIL139CZ0Z_1 ;
    wire \DUT.uart_inst0.m3_e_1_cascade_ ;
    wire DUT_uart_inst0_recv_state_2;
    wire \DUT.uart_inst0.rx_bits_remainingZ0Z_2 ;
    wire \DUT.uart_inst0.rx_bits_remainingZ0Z_3 ;
    wire \DUT.uart_inst0.rx_bits_remainingZ0Z_1 ;
    wire \DUT.uart_inst0.rx_bits_remainingZ0Z_0 ;
    wire \DUT.uart_inst0.recv_state_RNO_4Z0Z_2 ;
    wire \DUT.uart_inst0.N_19 ;
    wire \DUT.uart_inst0.G_8_i_a3_0_0 ;
    wire \DUT.uart_inst0.rx_countdown_8_i_o2_1_1_2 ;
    wire CONSTANT_ONE_NET;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_ ;
    wire \DUT.rFifoDatarx_7 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_7 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ;
    wire \DUT.rFifoDatarx_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1_cascade_ ;
    wire \DUT.rFifoDatarx_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_ ;
    wire \DUT.rFifoDatarx_4 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_4 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ;
    wire \DUT.rFifoDatarx_5 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_5 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_6 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_ ;
    wire \DUT.rFifoDatarx_6 ;
    wire \DUT.fifo_tx_inst.rFifoCountZ0Z_1 ;
    wire \DUT.fifo_tx_inst.rFifoCountZ0Z_0 ;
    wire \DUT.rTransmitZ0 ;
    wire \DUT.fifo_tx_inst.rFifoCountZ0Z_2 ;
    wire \DUT.fifo_tx_inst.rReadPtr11_cascade_ ;
    wire \DUT.fifo_tx_inst.un1_i11_2_i_cascade_ ;
    wire \DUT.fifo_tx_inst.rReadPtr11 ;
    wire \DUT.fifo_tx_inst.un1_i11_2_i ;
    wire \DUT.rFifoDataror_1 ;
    wire \DUT.rFifoDataror_1_cascade_ ;
    wire \DUT.rFifoDataror_0_0 ;
    wire \DUT.rFifoDataror_0 ;
    wire G_115;
    wire \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa ;
    wire \DUT.uart_inst0.m6_2 ;
    wire G_114;
    wire G_113;
    wire \fifo_inst.ftdi_input_inst.un1_rWrStateZ0Z_1_cascade_ ;
    wire G_118;
    wire G_118_cascade_;
    wire G_119;
    wire G_116;
    wire \fifo_inst.ftdi_input_inst.un1_rWrStateZ0Z_1 ;
    wire G_116_cascade_;
    wire G_117;
    wire \DUT.uart_inst0.g1_i_a4_1_5 ;
    wire \DUT.uart_inst0.g1_i_a4_1_3 ;
    wire \DUT.uart_inst0.N_78_cascade_ ;
    wire \DUT.uart_inst0.N_10_mux_cascade_ ;
    wire \DUT.uart_inst0.P6_mux ;
    wire \DUT.uart_inst0.G_19_0_a5_0_2_cascade_ ;
    wire \DUT.uart_inst0.G_19_0_1 ;
    wire \DUT.uart_inst0.G_19_0_a5_0_4_cascade_ ;
    wire \DUT.uart_inst0.rx_countdown_8_i_o2_2_0_2 ;
    wire \DUT.uart_inst0.G_8_i_a3_1 ;
    wire DUT_uart_inst0_rx_countdown_3_s1_4;
    wire DUT_uart_inst0_rx_countdown_3_s1_5;
    wire DUT_uart_inst0_rx_countdown_3_s1_3;
    wire \DUT.uart_inst0.rx_countdownZ0Z_3 ;
    wire DUT_uart_inst0_rx_countdown_3_s1_2;
    wire DUT_uart_inst0_rx_countdown_3_s1_1;
    wire \DUT.uart_inst0.G_19_0_a5_4 ;
    wire \DUT.uart_inst0.N_44 ;
    wire \DUT.fifo_rx_inst.N_77_mux ;
    wire \DUT.uart_inst0.g1_0 ;
    wire \DUT.uart_inst0.recv_stateZ0Z_0 ;
    wire \DUT.uart_inst0.recv_stateZ0Z_5 ;
    wire \DUT.uart_inst0.rx_countdown_8_i_a2_0_2 ;
    wire \DUT.uart_inst0.m10_e_3 ;
    wire \DUT.uart_inst0.m10_e_2 ;
    wire wPllLocked;
    wire \DUT.uart_inst0.N_20_mux_cascade_ ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_0 ;
    wire \DUT.uart_inst0.m7_3_cascade_ ;
    wire \DUT.uart_inst0.N_28_mux ;
    wire P1A1_c;
    wire \DUT.uart_inst0.m2_e_0 ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_5 ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_4 ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_1 ;
    wire \DUT.uart_inst0.recv_stateZ0Z_3 ;
    wire \DUT.uart_inst0.m6_e_2 ;
    wire \DUT.uart_inst0.m6_e_3_cascade_ ;
    wire \DUT.uart_inst0.N_15_mux ;
    wire \DUT.uart_inst0.N_18_mux_1 ;
    wire \DUT.uart_inst0.rx_countdownZ1Z_3 ;
    wire \DUT.uart_inst0.recv_stateZ0Z_4 ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_2 ;
    wire \DUT.uart_inst0.G_19_0_a5_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_4 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_5 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_6 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_7 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_ ;
    wire \DUT.rFifoDatarx_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_2 ;
    wire \DUT.fifo_tx_inst.rReadPtrZ0Z_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_3 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ;
    wire \DUT.fifo_tx_inst.rReadPtrZ0Z_1 ;
    wire \DUT.rFifoDatarx_3 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_3 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_3 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_4 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_5 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_6 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_7 ;
    wire \DUT.fifo_tx_inst.rFifoData_awe0 ;
    wire \DUT.fifo_tx_inst.rFifoDataro_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_awe1 ;
    wire \DUT.fifo_tx_inst.rFifoDataro_1 ;
    wire \DUT.fifo_tx_inst.rFifoDataro_2 ;
    wire \DUT.fifo_tx_inst.rFifoDataro_3 ;
    wire \DUT.fifo_rx_inst.N_57 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_6 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_6 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_7 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_7 ;
    wire \DUT.fifo_rx_inst.rFifoDataro_3 ;
    wire \DUT.fifo_rx_inst.rFifoDataror_1_0_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_3 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_3 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_4 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_4 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_5 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoDataro_0 ;
    wire \DUT.fifo_rx_inst.rFifoDataro_1 ;
    wire \DUT.fifo_rx_inst.rFifoDataro_2 ;
    wire \DUT.fifo_rx_inst.rWritePtrZ0Z_0 ;
    wire \DUT.fifo_rx_inst.rWritePtrZ0Z_1 ;
    wire \DUT.fifo_tx_inst.rWritePtrZ0Z_0 ;
    wire \DUT.fifo_tx_inst.rWritePtrZ0Z_1 ;
    wire \DUT.fifo_tx_inst.N_104 ;
    wire \DUT.fifo_tx_inst.rFifoData_awe2 ;
    wire \DUT.fifo_rx_inst.rWritePtr16_cascade_ ;
    wire \DUT.fifo_rx_inst.rWritePtr16 ;
    wire \DUT.wRcvd ;
    wire \DUT.fifo_rx_inst.N_46 ;
    wire N_69_mux;
    wire N_69_mux_cascade_;
    wire N_1258_i;
    wire P1A4_c_i;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_3 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_4 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_5 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_6 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_7 ;
    wire \DUT.fifo_tx_inst.rFifoData_awe3 ;
    wire ioFifoData_in_3;
    wire ioFifoData_in_1;
    wire ioFifoData_in_5;
    wire ioFifoData_in_2;
    wire ioFifoData_in_0;
    wire ioFifoData_in_6;
    wire ioFifoData_in_4;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_3 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_4 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_5 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_6 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_7 ;
    wire \DUT.fifo_rx_inst.rFifoData_awe2 ;
    wire \DUT.fifo_rx_inst.rFifoDatarx_6 ;
    wire wRxFifoData_6;
    wire rTxByteZ0Z_6;
    wire wRxFifoData_5;
    wire \DUT.fifo_rx_inst.rFifoDatarx_5 ;
    wire rTxByteZ0Z_5;
    wire wRxFifoData_0;
    wire rTxByteZ0Z_0;
    wire \DUT.fifo_rx_inst.rFifoDatarx_7 ;
    wire rTxByteZ0Z_7;
    wire wRxFifoData_1;
    wire rTxByteZ0Z_1;
    wire wRxFifoData_2;
    wire rTxByteZ0Z_2;
    wire \DUT.fifo_rx_inst.rFifoDatarx_3 ;
    wire wRxFifoData_3;
    wire rTxByteZ0Z_3;
    wire \DUT.fifo_rx_inst.rFifoDataror_0 ;
    wire wRxFifoData_4;
    wire \DUT.fifo_rx_inst.rFifoDatarx_4 ;
    wire rTxByteZ0Z_4;
    wire rTxByte_1_sqmuxa_i_0;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoDatarx_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_1 ;
    wire \DUT.fifo_rx_inst.rFifoDatarx_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_1 ;
    wire \DUT.fifo_rx_inst.rReadPtrZ0Z_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_2 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_2 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2_cascade_ ;
    wire \DUT.fifo_rx_inst.rReadPtrZ0Z_1 ;
    wire \DUT.fifo_rx_inst.rFifoDatarx_2 ;
    wire \DUT.wRxByte_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_0 ;
    wire \DUT.wRxByte_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_2 ;
    wire \DUT.wRxByte_3 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_3 ;
    wire \DUT.wRxByte_4 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_4 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_5 ;
    wire \DUT.wRxByte_6 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_6 ;
    wire \DUT.wRxByte_7 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_7 ;
    wire \DUT.fifo_rx_inst.rFifoData_awe1 ;
    wire \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0 ;
    wire \DUT.fifo_rx_inst.rFifoCountZ0Z_0 ;
    wire bfn_18_12_0_;
    wire \DUT.fifo_rx_inst.rFifoCount_RNIPTFQ1Z0Z_1 ;
    wire \DUT.fifo_rx_inst.rFifoCountZ0Z_1 ;
    wire \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0 ;
    wire \DUT.fifo_rx_inst.N_4_0 ;
    wire rRxReadZ0;
    wire \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1 ;
    wire \DUT.fifo_rx_inst.rFifoCountZ0Z_2 ;
    wire N_1261_i;
    wire oTx_n_rep4_ess;
    wire oTx_n_rep1_ess;
    wire oTx_n_rep0_ess;
    wire \fifo_inst.ftdi_output_inst.N_77_0_cascade_ ;
    wire P1A4_c;
    wire \fifo_inst.ftdi_output_inst.oPacketRead_1_sqmuxa_1_cascade_ ;
    wire \fifo_inst.wRamRdAddr_0 ;
    wire \fifo_inst.wRamRdAddr_1 ;
    wire \fifo_inst.ftdi_output_inst.oPacketRead_1_sqmuxa_1 ;
    wire \fifo_inst.wRamRdAddr_2 ;
    wire \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_3 ;
    wire P1A2_c;
    wire P1A3_c;
    wire \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1 ;
    wire iTxE_n_c;
    wire iRxF_n_c;
    wire G_120;
    wire wPllLocked_g;
    wire \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2 ;
    wire \fifo_inst.ftdi_output_inst.N_87_cascade_ ;
    wire \fifo_inst.ftdi_output_inst.N_77_0 ;
    wire \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0 ;
    wire ioFifoData_in_7;
    wire wRxFifoData_7;
    wire \fifo_inst.ftdi_output_inst.rFifoState_0_1 ;
    wire N_1260_i;
    wire N_1259_i;
    wire oTx_n_rep3_ess;
    wire \fifo_inst.ftdi_output_inst.rWrDelayZ0 ;
    wire \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4 ;
    wire oTx_n_rep2_ess;
    wire \fifo_inst.ftdi_output_inst.N_88_i_0 ;
    wire wPllLocked_iso_i_g;
    wire \DUT.wRxByte_2 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_2 ;
    wire \DUT.wRxByte_5 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_5 ;
    wire clk_48mhz;
    wire \DUT.fifo_rx_inst.rFifoData_awe0 ;
    wire _gnd_net_;

    defparam \fifo_inst.ftdi_input_inst.ram512x8_inst_physical .WRITE_MODE=1;
    defparam \fifo_inst.ftdi_input_inst.ram512x8_inst_physical .READ_MODE=1;
    SB_RAM40_4K \fifo_inst.ftdi_input_inst.ram512x8_inst_physical  (
            .RDATA({dangling_wire_0,wRamRdData_7,dangling_wire_1,wRamRdData_6,dangling_wire_2,wRamRdData_5,dangling_wire_3,wRamRdData_4,dangling_wire_4,wRamRdData_3,dangling_wire_5,wRamRdData_2,dangling_wire_6,wRamRdData_1,dangling_wire_7,wRamRdData_0}),
            .RADDR({dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,N__14130,N__14157,N__14178}),
            .WADDR({dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,N__9711,N__9648,N__9684}),
            .MASK({dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39}),
            .WDATA({dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55}),
            .RCLKE(),
            .RCLK(GNDG0),
            .RE(N__9179),
            .WCLKE(),
            .WCLK(N__15047),
            .WE(N__9569));
    defparam \top_pll_inst.top_pll_inst_pll .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \top_pll_inst.top_pll_inst_pll .TEST_MODE=1'b0;
    defparam \top_pll_inst.top_pll_inst_pll .SHIFTREG_DIV_MODE=2'b00;
    defparam \top_pll_inst.top_pll_inst_pll .PLLOUT_SELECT="GENCLK";
    defparam \top_pll_inst.top_pll_inst_pll .FILTER_RANGE=3'b001;
    defparam \top_pll_inst.top_pll_inst_pll .FEEDBACK_PATH="SIMPLE";
    defparam \top_pll_inst.top_pll_inst_pll .FDA_RELATIVE=4'b0000;
    defparam \top_pll_inst.top_pll_inst_pll .FDA_FEEDBACK=4'b0000;
    defparam \top_pll_inst.top_pll_inst_pll .ENABLE_ICEGATE=1'b0;
    defparam \top_pll_inst.top_pll_inst_pll .DIVR=4'b0000;
    defparam \top_pll_inst.top_pll_inst_pll .DIVQ=3'b100;
    defparam \top_pll_inst.top_pll_inst_pll .DIVF=7'b0111111;
    defparam \top_pll_inst.top_pll_inst_pll .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    PLL40 \top_pll_inst.top_pll_inst_pll  (
            .PLLOUTGLOBAL(clk_48mhz),
            .SDI(GNDG0),
            .BYPASS(GNDG0),
            .RESETB(N__5949),
            .PLLOUTCORE(),
            .LOCK(\PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO ),
            .SDO(),
            .SCLK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .EXTFEEDBACK(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLIN(N__15651));
    IO_PAD \top_pll_inst.top_pll_inst_iopad  (
            .OE(VCCG0),
            .DIN(),
            .DOUT(N__15651),
            .PACKAGEPIN(iClk));
    IO_PAD P1A8_obuft_iopad (
            .OE(N__15637),
            .DIN(N__15636),
            .DOUT(N__15635),
            .PACKAGEPIN(P1A8));
    defparam P1A8_obuft_preio.NEG_TRIGGER=1'b0;
    defparam P1A8_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO P1A8_obuft_preio (
            .PADOEN(N__15637),
            .PADOUT(N__15636),
            .PADIN(N__15635),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_3_iopad (
            .OE(N__15628),
            .DIN(N__15627),
            .DOUT(N__15626),
            .PACKAGEPIN(ioFifoData[3]));
    defparam ioFifoData_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_3_preio (
            .PADOEN(N__15628),
            .PADOUT(N__15627),
            .PADIN(N__15626),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__15447),
            .DIN0(ioFifoData_in_3),
            .DOUT0(N__5988),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A4_obuf_iopad (
            .OE(N__15619),
            .DIN(N__15618),
            .DOUT(N__15617),
            .PACKAGEPIN(P1A4));
    defparam P1A4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO P1A4_obuf_preio (
            .PADOEN(N__15619),
            .PADOUT(N__15618),
            .PADIN(N__15617),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14232),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD oRx_n_obuf_iopad (
            .OE(N__15610),
            .DIN(N__15609),
            .DOUT(N__15608),
            .PACKAGEPIN(oRx_n));
    defparam oRx_n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam oRx_n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO oRx_n_obuf_preio (
            .PADOEN(N__15610),
            .PADOUT(N__15609),
            .PADIN(N__15608),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14723),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A2_obuf_iopad (
            .OE(N__15601),
            .DIN(N__15600),
            .DOUT(N__15599),
            .PACKAGEPIN(P1A2));
    defparam P1A2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO P1A2_obuf_preio (
            .PADOEN(N__15601),
            .PADOUT(N__15600),
            .PADIN(N__15599),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14825),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_0_iopad (
            .OE(N__15592),
            .DIN(N__15591),
            .DOUT(N__15590),
            .PACKAGEPIN(ioFifoData[0]));
    defparam ioFifoData_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_0_preio (
            .PADOEN(N__15592),
            .PADOUT(N__15591),
            .PADIN(N__15590),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7704),
            .DIN0(ioFifoData_in_0),
            .DOUT0(N__6006),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD iRxF_n_ibuf_iopad (
            .OE(N__15583),
            .DIN(N__15582),
            .DOUT(N__15581),
            .PACKAGEPIN(iRxF_n));
    defparam iRxF_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam iRxF_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO iRxF_n_ibuf_preio (
            .PADOEN(N__15583),
            .PADOUT(N__15582),
            .PADIN(N__15581),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(iRxF_n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A3_obuf_iopad (
            .OE(N__15574),
            .DIN(N__15573),
            .DOUT(N__15572),
            .PACKAGEPIN(P1A3));
    defparam P1A3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO P1A3_obuf_preio (
            .PADOEN(N__15574),
            .PADOUT(N__15573),
            .PADIN(N__15572),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14730),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A7_obuf_iopad (
            .OE(N__15565),
            .DIN(N__15564),
            .DOUT(N__15563),
            .PACKAGEPIN(P1A7));
    defparam P1A7_obuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A7_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO P1A7_obuf_preio (
            .PADOEN(N__15565),
            .PADOUT(N__15564),
            .PADIN(N__15563),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7779),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_7_iopad (
            .OE(N__15556),
            .DIN(N__15555),
            .DOUT(N__15554),
            .PACKAGEPIN(ioFifoData[7]));
    defparam ioFifoData_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_7_preio (
            .PADOEN(N__15556),
            .PADOUT(N__15555),
            .PADIN(N__15554),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__12513),
            .DIN0(ioFifoData_in_7),
            .DOUT0(N__5934),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BTN_N_ibuf_iopad (
            .OE(N__15547),
            .DIN(N__15546),
            .DOUT(N__15545),
            .PACKAGEPIN(BTN_N));
    defparam BTN_N_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam BTN_N_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO BTN_N_ibuf_preio (
            .PADOEN(N__15547),
            .PADOUT(N__15546),
            .PADIN(N__15545),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(BTN_N_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_4_iopad (
            .OE(N__15538),
            .DIN(N__15537),
            .DOUT(N__15536),
            .PACKAGEPIN(ioFifoData[4]));
    defparam ioFifoData_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_4_preio (
            .PADOEN(N__15538),
            .PADOUT(N__15537),
            .PADIN(N__15536),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__13872),
            .DIN0(ioFifoData_in_4),
            .DOUT0(N__5961),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_1_iopad (
            .OE(N__15529),
            .DIN(N__15528),
            .DOUT(N__15527),
            .PACKAGEPIN(ioFifoData[1]));
    defparam ioFifoData_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_1_preio (
            .PADOEN(N__15529),
            .PADOUT(N__15528),
            .PADIN(N__15527),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__12525),
            .DIN0(ioFifoData_in_1),
            .DOUT0(N__5919),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_5_iopad (
            .OE(N__15520),
            .DIN(N__15519),
            .DOUT(N__15518),
            .PACKAGEPIN(ioFifoData[5]));
    defparam ioFifoData_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_5_preio (
            .PADOEN(N__15520),
            .PADOUT(N__15519),
            .PADIN(N__15518),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__12491),
            .DIN0(ioFifoData_in_5),
            .DOUT0(N__5871),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD oTx_n_obuf_iopad (
            .OE(N__15511),
            .DIN(N__15510),
            .DOUT(N__15509),
            .PACKAGEPIN(oTx_n));
    defparam oTx_n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam oTx_n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO oTx_n_obuf_preio (
            .PADOEN(N__15511),
            .PADOUT(N__15510),
            .PADIN(N__15509),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14225),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD iTxE_n_ibuf_iopad (
            .OE(N__15502),
            .DIN(N__15501),
            .DOUT(N__15500),
            .PACKAGEPIN(iTxE_n));
    defparam iTxE_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam iTxE_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO iTxE_n_ibuf_preio (
            .PADOEN(N__15502),
            .PADOUT(N__15501),
            .PADIN(N__15500),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(iTxE_n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A1_ibuf_iopad (
            .OE(N__15493),
            .DIN(N__15492),
            .DOUT(N__15491),
            .PACKAGEPIN(P1A1));
    defparam P1A1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO P1A1_ibuf_preio (
            .PADOEN(N__15493),
            .PADOUT(N__15492),
            .PADIN(N__15491),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(P1A1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_2_iopad (
            .OE(N__15484),
            .DIN(N__15483),
            .DOUT(N__15482),
            .PACKAGEPIN(ioFifoData[2]));
    defparam ioFifoData_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_2_preio (
            .PADOEN(N__15484),
            .PADOUT(N__15483),
            .PADIN(N__15482),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__15441),
            .DIN0(ioFifoData_in_2),
            .DOUT0(N__5886),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A9_obuft_iopad (
            .OE(N__15475),
            .DIN(N__15474),
            .DOUT(N__15473),
            .PACKAGEPIN(P1A9));
    defparam P1A9_obuft_preio.NEG_TRIGGER=1'b0;
    defparam P1A9_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO P1A9_obuft_preio (
            .PADOEN(N__15475),
            .PADOUT(N__15474),
            .PADIN(N__15473),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_6_iopad (
            .OE(N__15466),
            .DIN(N__15465),
            .DOUT(N__15464),
            .PACKAGEPIN(ioFifoData[6]));
    defparam ioFifoData_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_6_preio (
            .PADOEN(N__15466),
            .PADOUT(N__15465),
            .PADIN(N__15464),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__12512),
            .DIN0(ioFifoData_in_6),
            .DOUT0(N__5901),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IoInMux I__3682 (
            .O(N__15447),
            .I(N__15444));
    LocalMux I__3681 (
            .O(N__15444),
            .I(N_1260_i));
    IoInMux I__3680 (
            .O(N__15441),
            .I(N__15438));
    LocalMux I__3679 (
            .O(N__15438),
            .I(N__15435));
    Odrv4 I__3678 (
            .O(N__15435),
            .I(N_1259_i));
    InMux I__3677 (
            .O(N__15432),
            .I(N__15429));
    LocalMux I__3676 (
            .O(N__15429),
            .I(N__15426));
    Odrv12 I__3675 (
            .O(N__15426),
            .I(oTx_n_rep3_ess));
    CascadeMux I__3674 (
            .O(N__15423),
            .I(N__15418));
    CascadeMux I__3673 (
            .O(N__15422),
            .I(N__15414));
    CascadeMux I__3672 (
            .O(N__15421),
            .I(N__15411));
    InMux I__3671 (
            .O(N__15418),
            .I(N__15403));
    InMux I__3670 (
            .O(N__15417),
            .I(N__15403));
    InMux I__3669 (
            .O(N__15414),
            .I(N__15396));
    InMux I__3668 (
            .O(N__15411),
            .I(N__15396));
    InMux I__3667 (
            .O(N__15410),
            .I(N__15396));
    CascadeMux I__3666 (
            .O(N__15409),
            .I(N__15393));
    CascadeMux I__3665 (
            .O(N__15408),
            .I(N__15389));
    LocalMux I__3664 (
            .O(N__15403),
            .I(N__15384));
    LocalMux I__3663 (
            .O(N__15396),
            .I(N__15381));
    InMux I__3662 (
            .O(N__15393),
            .I(N__15376));
    InMux I__3661 (
            .O(N__15392),
            .I(N__15376));
    InMux I__3660 (
            .O(N__15389),
            .I(N__15369));
    InMux I__3659 (
            .O(N__15388),
            .I(N__15369));
    InMux I__3658 (
            .O(N__15387),
            .I(N__15369));
    Odrv4 I__3657 (
            .O(N__15384),
            .I(\fifo_inst.ftdi_output_inst.rWrDelayZ0 ));
    Odrv4 I__3656 (
            .O(N__15381),
            .I(\fifo_inst.ftdi_output_inst.rWrDelayZ0 ));
    LocalMux I__3655 (
            .O(N__15376),
            .I(\fifo_inst.ftdi_output_inst.rWrDelayZ0 ));
    LocalMux I__3654 (
            .O(N__15369),
            .I(\fifo_inst.ftdi_output_inst.rWrDelayZ0 ));
    InMux I__3653 (
            .O(N__15360),
            .I(N__15351));
    InMux I__3652 (
            .O(N__15359),
            .I(N__15351));
    InMux I__3651 (
            .O(N__15358),
            .I(N__15344));
    InMux I__3650 (
            .O(N__15357),
            .I(N__15344));
    InMux I__3649 (
            .O(N__15356),
            .I(N__15344));
    LocalMux I__3648 (
            .O(N__15351),
            .I(N__15336));
    LocalMux I__3647 (
            .O(N__15344),
            .I(N__15333));
    InMux I__3646 (
            .O(N__15343),
            .I(N__15328));
    InMux I__3645 (
            .O(N__15342),
            .I(N__15328));
    InMux I__3644 (
            .O(N__15341),
            .I(N__15321));
    InMux I__3643 (
            .O(N__15340),
            .I(N__15321));
    InMux I__3642 (
            .O(N__15339),
            .I(N__15321));
    Odrv4 I__3641 (
            .O(N__15336),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4 ));
    Odrv4 I__3640 (
            .O(N__15333),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4 ));
    LocalMux I__3639 (
            .O(N__15328),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4 ));
    LocalMux I__3638 (
            .O(N__15321),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4 ));
    InMux I__3637 (
            .O(N__15312),
            .I(N__15309));
    LocalMux I__3636 (
            .O(N__15309),
            .I(N__15306));
    Odrv4 I__3635 (
            .O(N__15306),
            .I(oTx_n_rep2_ess));
    CEMux I__3634 (
            .O(N__15303),
            .I(N__15299));
    CEMux I__3633 (
            .O(N__15302),
            .I(N__15296));
    LocalMux I__3632 (
            .O(N__15299),
            .I(\fifo_inst.ftdi_output_inst.N_88_i_0 ));
    LocalMux I__3631 (
            .O(N__15296),
            .I(\fifo_inst.ftdi_output_inst.N_88_i_0 ));
    CascadeMux I__3630 (
            .O(N__15291),
            .I(N__15287));
    InMux I__3629 (
            .O(N__15290),
            .I(N__15275));
    InMux I__3628 (
            .O(N__15287),
            .I(N__15266));
    InMux I__3627 (
            .O(N__15286),
            .I(N__15266));
    InMux I__3626 (
            .O(N__15285),
            .I(N__15266));
    InMux I__3625 (
            .O(N__15284),
            .I(N__15266));
    InMux I__3624 (
            .O(N__15283),
            .I(N__15263));
    InMux I__3623 (
            .O(N__15282),
            .I(N__15260));
    InMux I__3622 (
            .O(N__15281),
            .I(N__15253));
    InMux I__3621 (
            .O(N__15280),
            .I(N__15253));
    InMux I__3620 (
            .O(N__15279),
            .I(N__15253));
    InMux I__3619 (
            .O(N__15278),
            .I(N__15250));
    LocalMux I__3618 (
            .O(N__15275),
            .I(N__15245));
    LocalMux I__3617 (
            .O(N__15266),
            .I(N__15242));
    LocalMux I__3616 (
            .O(N__15263),
            .I(N__15237));
    LocalMux I__3615 (
            .O(N__15260),
            .I(N__15233));
    LocalMux I__3614 (
            .O(N__15253),
            .I(N__15226));
    LocalMux I__3613 (
            .O(N__15250),
            .I(N__15220));
    SRMux I__3612 (
            .O(N__15249),
            .I(N__15177));
    SRMux I__3611 (
            .O(N__15248),
            .I(N__15177));
    Glb2LocalMux I__3610 (
            .O(N__15245),
            .I(N__15177));
    Glb2LocalMux I__3609 (
            .O(N__15242),
            .I(N__15177));
    SRMux I__3608 (
            .O(N__15241),
            .I(N__15177));
    SRMux I__3607 (
            .O(N__15240),
            .I(N__15177));
    Glb2LocalMux I__3606 (
            .O(N__15237),
            .I(N__15177));
    SRMux I__3605 (
            .O(N__15236),
            .I(N__15177));
    Glb2LocalMux I__3604 (
            .O(N__15233),
            .I(N__15177));
    SRMux I__3603 (
            .O(N__15232),
            .I(N__15177));
    SRMux I__3602 (
            .O(N__15231),
            .I(N__15177));
    SRMux I__3601 (
            .O(N__15230),
            .I(N__15177));
    SRMux I__3600 (
            .O(N__15229),
            .I(N__15177));
    Glb2LocalMux I__3599 (
            .O(N__15226),
            .I(N__15177));
    SRMux I__3598 (
            .O(N__15225),
            .I(N__15177));
    SRMux I__3597 (
            .O(N__15224),
            .I(N__15177));
    SRMux I__3596 (
            .O(N__15223),
            .I(N__15177));
    Glb2LocalMux I__3595 (
            .O(N__15220),
            .I(N__15177));
    SRMux I__3594 (
            .O(N__15219),
            .I(N__15177));
    SRMux I__3593 (
            .O(N__15218),
            .I(N__15177));
    GlobalMux I__3592 (
            .O(N__15177),
            .I(N__15174));
    gio2CtrlBuf I__3591 (
            .O(N__15174),
            .I(wPllLocked_iso_i_g));
    InMux I__3590 (
            .O(N__15171),
            .I(N__15168));
    LocalMux I__3589 (
            .O(N__15168),
            .I(N__15163));
    InMux I__3588 (
            .O(N__15167),
            .I(N__15160));
    InMux I__3587 (
            .O(N__15166),
            .I(N__15157));
    Span4Mux_h I__3586 (
            .O(N__15163),
            .I(N__15154));
    LocalMux I__3585 (
            .O(N__15160),
            .I(N__15151));
    LocalMux I__3584 (
            .O(N__15157),
            .I(N__15148));
    Span4Mux_h I__3583 (
            .O(N__15154),
            .I(N__15143));
    Span4Mux_v I__3582 (
            .O(N__15151),
            .I(N__15140));
    Span4Mux_h I__3581 (
            .O(N__15148),
            .I(N__15137));
    InMux I__3580 (
            .O(N__15147),
            .I(N__15134));
    InMux I__3579 (
            .O(N__15146),
            .I(N__15131));
    Odrv4 I__3578 (
            .O(N__15143),
            .I(\DUT.wRxByte_2 ));
    Odrv4 I__3577 (
            .O(N__15140),
            .I(\DUT.wRxByte_2 ));
    Odrv4 I__3576 (
            .O(N__15137),
            .I(\DUT.wRxByte_2 ));
    LocalMux I__3575 (
            .O(N__15134),
            .I(\DUT.wRxByte_2 ));
    LocalMux I__3574 (
            .O(N__15131),
            .I(\DUT.wRxByte_2 ));
    InMux I__3573 (
            .O(N__15120),
            .I(N__15117));
    LocalMux I__3572 (
            .O(N__15117),
            .I(N__15114));
    Odrv12 I__3571 (
            .O(N__15114),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_2 ));
    InMux I__3570 (
            .O(N__15111),
            .I(N__15107));
    InMux I__3569 (
            .O(N__15110),
            .I(N__15103));
    LocalMux I__3568 (
            .O(N__15107),
            .I(N__15100));
    InMux I__3567 (
            .O(N__15106),
            .I(N__15097));
    LocalMux I__3566 (
            .O(N__15103),
            .I(N__15094));
    Span4Mux_v I__3565 (
            .O(N__15100),
            .I(N__15089));
    LocalMux I__3564 (
            .O(N__15097),
            .I(N__15089));
    Span4Mux_v I__3563 (
            .O(N__15094),
            .I(N__15086));
    Sp12to4 I__3562 (
            .O(N__15089),
            .I(N__15083));
    Sp12to4 I__3561 (
            .O(N__15086),
            .I(N__15076));
    Span12Mux_s6_v I__3560 (
            .O(N__15083),
            .I(N__15076));
    InMux I__3559 (
            .O(N__15082),
            .I(N__15073));
    InMux I__3558 (
            .O(N__15081),
            .I(N__15070));
    Odrv12 I__3557 (
            .O(N__15076),
            .I(\DUT.wRxByte_5 ));
    LocalMux I__3556 (
            .O(N__15073),
            .I(\DUT.wRxByte_5 ));
    LocalMux I__3555 (
            .O(N__15070),
            .I(\DUT.wRxByte_5 ));
    InMux I__3554 (
            .O(N__15063),
            .I(N__15060));
    LocalMux I__3553 (
            .O(N__15060),
            .I(N__15057));
    Odrv12 I__3552 (
            .O(N__15057),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_5 ));
    ClkMux I__3551 (
            .O(N__15054),
            .I(N__14871));
    ClkMux I__3550 (
            .O(N__15053),
            .I(N__14871));
    ClkMux I__3549 (
            .O(N__15052),
            .I(N__14871));
    ClkMux I__3548 (
            .O(N__15051),
            .I(N__14871));
    ClkMux I__3547 (
            .O(N__15050),
            .I(N__14871));
    ClkMux I__3546 (
            .O(N__15049),
            .I(N__14871));
    ClkMux I__3545 (
            .O(N__15048),
            .I(N__14871));
    ClkMux I__3544 (
            .O(N__15047),
            .I(N__14871));
    ClkMux I__3543 (
            .O(N__15046),
            .I(N__14871));
    ClkMux I__3542 (
            .O(N__15045),
            .I(N__14871));
    ClkMux I__3541 (
            .O(N__15044),
            .I(N__14871));
    ClkMux I__3540 (
            .O(N__15043),
            .I(N__14871));
    ClkMux I__3539 (
            .O(N__15042),
            .I(N__14871));
    ClkMux I__3538 (
            .O(N__15041),
            .I(N__14871));
    ClkMux I__3537 (
            .O(N__15040),
            .I(N__14871));
    ClkMux I__3536 (
            .O(N__15039),
            .I(N__14871));
    ClkMux I__3535 (
            .O(N__15038),
            .I(N__14871));
    ClkMux I__3534 (
            .O(N__15037),
            .I(N__14871));
    ClkMux I__3533 (
            .O(N__15036),
            .I(N__14871));
    ClkMux I__3532 (
            .O(N__15035),
            .I(N__14871));
    ClkMux I__3531 (
            .O(N__15034),
            .I(N__14871));
    ClkMux I__3530 (
            .O(N__15033),
            .I(N__14871));
    ClkMux I__3529 (
            .O(N__15032),
            .I(N__14871));
    ClkMux I__3528 (
            .O(N__15031),
            .I(N__14871));
    ClkMux I__3527 (
            .O(N__15030),
            .I(N__14871));
    ClkMux I__3526 (
            .O(N__15029),
            .I(N__14871));
    ClkMux I__3525 (
            .O(N__15028),
            .I(N__14871));
    ClkMux I__3524 (
            .O(N__15027),
            .I(N__14871));
    ClkMux I__3523 (
            .O(N__15026),
            .I(N__14871));
    ClkMux I__3522 (
            .O(N__15025),
            .I(N__14871));
    ClkMux I__3521 (
            .O(N__15024),
            .I(N__14871));
    ClkMux I__3520 (
            .O(N__15023),
            .I(N__14871));
    ClkMux I__3519 (
            .O(N__15022),
            .I(N__14871));
    ClkMux I__3518 (
            .O(N__15021),
            .I(N__14871));
    ClkMux I__3517 (
            .O(N__15020),
            .I(N__14871));
    ClkMux I__3516 (
            .O(N__15019),
            .I(N__14871));
    ClkMux I__3515 (
            .O(N__15018),
            .I(N__14871));
    ClkMux I__3514 (
            .O(N__15017),
            .I(N__14871));
    ClkMux I__3513 (
            .O(N__15016),
            .I(N__14871));
    ClkMux I__3512 (
            .O(N__15015),
            .I(N__14871));
    ClkMux I__3511 (
            .O(N__15014),
            .I(N__14871));
    ClkMux I__3510 (
            .O(N__15013),
            .I(N__14871));
    ClkMux I__3509 (
            .O(N__15012),
            .I(N__14871));
    ClkMux I__3508 (
            .O(N__15011),
            .I(N__14871));
    ClkMux I__3507 (
            .O(N__15010),
            .I(N__14871));
    ClkMux I__3506 (
            .O(N__15009),
            .I(N__14871));
    ClkMux I__3505 (
            .O(N__15008),
            .I(N__14871));
    ClkMux I__3504 (
            .O(N__15007),
            .I(N__14871));
    ClkMux I__3503 (
            .O(N__15006),
            .I(N__14871));
    ClkMux I__3502 (
            .O(N__15005),
            .I(N__14871));
    ClkMux I__3501 (
            .O(N__15004),
            .I(N__14871));
    ClkMux I__3500 (
            .O(N__15003),
            .I(N__14871));
    ClkMux I__3499 (
            .O(N__15002),
            .I(N__14871));
    ClkMux I__3498 (
            .O(N__15001),
            .I(N__14871));
    ClkMux I__3497 (
            .O(N__15000),
            .I(N__14871));
    ClkMux I__3496 (
            .O(N__14999),
            .I(N__14871));
    ClkMux I__3495 (
            .O(N__14998),
            .I(N__14871));
    ClkMux I__3494 (
            .O(N__14997),
            .I(N__14871));
    ClkMux I__3493 (
            .O(N__14996),
            .I(N__14871));
    ClkMux I__3492 (
            .O(N__14995),
            .I(N__14871));
    ClkMux I__3491 (
            .O(N__14994),
            .I(N__14871));
    GlobalMux I__3490 (
            .O(N__14871),
            .I(clk_48mhz));
    CEMux I__3489 (
            .O(N__14868),
            .I(N__14863));
    CEMux I__3488 (
            .O(N__14867),
            .I(N__14860));
    CEMux I__3487 (
            .O(N__14866),
            .I(N__14856));
    LocalMux I__3486 (
            .O(N__14863),
            .I(N__14853));
    LocalMux I__3485 (
            .O(N__14860),
            .I(N__14850));
    CEMux I__3484 (
            .O(N__14859),
            .I(N__14847));
    LocalMux I__3483 (
            .O(N__14856),
            .I(N__14844));
    Span4Mux_h I__3482 (
            .O(N__14853),
            .I(N__14839));
    Span4Mux_h I__3481 (
            .O(N__14850),
            .I(N__14839));
    LocalMux I__3480 (
            .O(N__14847),
            .I(N__14836));
    Span4Mux_v I__3479 (
            .O(N__14844),
            .I(N__14833));
    Odrv4 I__3478 (
            .O(N__14839),
            .I(\DUT.fifo_rx_inst.rFifoData_awe0 ));
    Odrv4 I__3477 (
            .O(N__14836),
            .I(\DUT.fifo_rx_inst.rFifoData_awe0 ));
    Odrv4 I__3476 (
            .O(N__14833),
            .I(\DUT.fifo_rx_inst.rFifoData_awe0 ));
    CascadeMux I__3475 (
            .O(N__14826),
            .I(N__14820));
    IoInMux I__3474 (
            .O(N__14825),
            .I(N__14809));
    InMux I__3473 (
            .O(N__14824),
            .I(N__14806));
    InMux I__3472 (
            .O(N__14823),
            .I(N__14789));
    InMux I__3471 (
            .O(N__14820),
            .I(N__14789));
    InMux I__3470 (
            .O(N__14819),
            .I(N__14789));
    InMux I__3469 (
            .O(N__14818),
            .I(N__14789));
    InMux I__3468 (
            .O(N__14817),
            .I(N__14789));
    InMux I__3467 (
            .O(N__14816),
            .I(N__14789));
    InMux I__3466 (
            .O(N__14815),
            .I(N__14789));
    InMux I__3465 (
            .O(N__14814),
            .I(N__14789));
    InMux I__3464 (
            .O(N__14813),
            .I(N__14786));
    InMux I__3463 (
            .O(N__14812),
            .I(N__14783));
    LocalMux I__3462 (
            .O(N__14809),
            .I(N__14780));
    LocalMux I__3461 (
            .O(N__14806),
            .I(N__14777));
    LocalMux I__3460 (
            .O(N__14789),
            .I(N__14774));
    LocalMux I__3459 (
            .O(N__14786),
            .I(N__14770));
    LocalMux I__3458 (
            .O(N__14783),
            .I(N__14767));
    Span12Mux_s1_v I__3457 (
            .O(N__14780),
            .I(N__14764));
    Span4Mux_h I__3456 (
            .O(N__14777),
            .I(N__14761));
    Span4Mux_v I__3455 (
            .O(N__14774),
            .I(N__14758));
    InMux I__3454 (
            .O(N__14773),
            .I(N__14755));
    Span4Mux_h I__3453 (
            .O(N__14770),
            .I(N__14750));
    Span4Mux_h I__3452 (
            .O(N__14767),
            .I(N__14750));
    Span12Mux_h I__3451 (
            .O(N__14764),
            .I(N__14747));
    Span4Mux_h I__3450 (
            .O(N__14761),
            .I(N__14744));
    Span4Mux_h I__3449 (
            .O(N__14758),
            .I(N__14737));
    LocalMux I__3448 (
            .O(N__14755),
            .I(N__14737));
    Span4Mux_v I__3447 (
            .O(N__14750),
            .I(N__14737));
    Odrv12 I__3446 (
            .O(N__14747),
            .I(P1A2_c));
    Odrv4 I__3445 (
            .O(N__14744),
            .I(P1A2_c));
    Odrv4 I__3444 (
            .O(N__14737),
            .I(P1A2_c));
    IoInMux I__3443 (
            .O(N__14730),
            .I(N__14727));
    LocalMux I__3442 (
            .O(N__14727),
            .I(N__14724));
    IoSpan4Mux I__3441 (
            .O(N__14724),
            .I(N__14720));
    IoInMux I__3440 (
            .O(N__14723),
            .I(N__14717));
    Sp12to4 I__3439 (
            .O(N__14720),
            .I(N__14714));
    LocalMux I__3438 (
            .O(N__14717),
            .I(N__14711));
    Span12Mux_s7_v I__3437 (
            .O(N__14714),
            .I(N__14707));
    Span12Mux_s7_v I__3436 (
            .O(N__14711),
            .I(N__14704));
    InMux I__3435 (
            .O(N__14710),
            .I(N__14701));
    Odrv12 I__3434 (
            .O(N__14707),
            .I(P1A3_c));
    Odrv12 I__3433 (
            .O(N__14704),
            .I(P1A3_c));
    LocalMux I__3432 (
            .O(N__14701),
            .I(P1A3_c));
    InMux I__3431 (
            .O(N__14694),
            .I(N__14687));
    InMux I__3430 (
            .O(N__14693),
            .I(N__14687));
    InMux I__3429 (
            .O(N__14692),
            .I(N__14684));
    LocalMux I__3428 (
            .O(N__14687),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1 ));
    LocalMux I__3427 (
            .O(N__14684),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1 ));
    CascadeMux I__3426 (
            .O(N__14679),
            .I(N__14676));
    InMux I__3425 (
            .O(N__14676),
            .I(N__14673));
    LocalMux I__3424 (
            .O(N__14673),
            .I(N__14670));
    Span4Mux_v I__3423 (
            .O(N__14670),
            .I(N__14666));
    InMux I__3422 (
            .O(N__14669),
            .I(N__14663));
    Sp12to4 I__3421 (
            .O(N__14666),
            .I(N__14658));
    LocalMux I__3420 (
            .O(N__14663),
            .I(N__14658));
    Span12Mux_s7_h I__3419 (
            .O(N__14658),
            .I(N__14655));
    Span12Mux_v I__3418 (
            .O(N__14655),
            .I(N__14652));
    Odrv12 I__3417 (
            .O(N__14652),
            .I(iTxE_n_c));
    CascadeMux I__3416 (
            .O(N__14649),
            .I(N__14644));
    InMux I__3415 (
            .O(N__14648),
            .I(N__14637));
    InMux I__3414 (
            .O(N__14647),
            .I(N__14637));
    InMux I__3413 (
            .O(N__14644),
            .I(N__14637));
    LocalMux I__3412 (
            .O(N__14637),
            .I(N__14633));
    InMux I__3411 (
            .O(N__14636),
            .I(N__14630));
    Span4Mux_v I__3410 (
            .O(N__14633),
            .I(N__14627));
    LocalMux I__3409 (
            .O(N__14630),
            .I(N__14624));
    Sp12to4 I__3408 (
            .O(N__14627),
            .I(N__14621));
    Span4Mux_h I__3407 (
            .O(N__14624),
            .I(N__14618));
    Span12Mux_s7_h I__3406 (
            .O(N__14621),
            .I(N__14613));
    Sp12to4 I__3405 (
            .O(N__14618),
            .I(N__14613));
    Span12Mux_v I__3404 (
            .O(N__14613),
            .I(N__14610));
    Odrv12 I__3403 (
            .O(N__14610),
            .I(iRxF_n_c));
    CascadeMux I__3402 (
            .O(N__14607),
            .I(N__14604));
    InMux I__3401 (
            .O(N__14604),
            .I(N__14600));
    InMux I__3400 (
            .O(N__14603),
            .I(N__14597));
    LocalMux I__3399 (
            .O(N__14600),
            .I(N__14592));
    LocalMux I__3398 (
            .O(N__14597),
            .I(N__14592));
    Span4Mux_v I__3397 (
            .O(N__14592),
            .I(N__14589));
    Span4Mux_h I__3396 (
            .O(N__14589),
            .I(N__14585));
    InMux I__3395 (
            .O(N__14588),
            .I(N__14582));
    Odrv4 I__3394 (
            .O(N__14585),
            .I(G_120));
    LocalMux I__3393 (
            .O(N__14582),
            .I(G_120));
    CascadeMux I__3392 (
            .O(N__14577),
            .I(N__14568));
    CascadeMux I__3391 (
            .O(N__14576),
            .I(N__14558));
    CascadeMux I__3390 (
            .O(N__14575),
            .I(N__14553));
    InMux I__3389 (
            .O(N__14574),
            .I(N__14543));
    InMux I__3388 (
            .O(N__14573),
            .I(N__14540));
    InMux I__3387 (
            .O(N__14572),
            .I(N__14537));
    InMux I__3386 (
            .O(N__14571),
            .I(N__14530));
    InMux I__3385 (
            .O(N__14568),
            .I(N__14530));
    InMux I__3384 (
            .O(N__14567),
            .I(N__14530));
    InMux I__3383 (
            .O(N__14566),
            .I(N__14527));
    InMux I__3382 (
            .O(N__14565),
            .I(N__14522));
    InMux I__3381 (
            .O(N__14564),
            .I(N__14522));
    InMux I__3380 (
            .O(N__14563),
            .I(N__14517));
    InMux I__3379 (
            .O(N__14562),
            .I(N__14517));
    InMux I__3378 (
            .O(N__14561),
            .I(N__14514));
    InMux I__3377 (
            .O(N__14558),
            .I(N__14511));
    InMux I__3376 (
            .O(N__14557),
            .I(N__14508));
    InMux I__3375 (
            .O(N__14556),
            .I(N__14505));
    InMux I__3374 (
            .O(N__14553),
            .I(N__14502));
    InMux I__3373 (
            .O(N__14552),
            .I(N__14497));
    InMux I__3372 (
            .O(N__14551),
            .I(N__14497));
    InMux I__3371 (
            .O(N__14550),
            .I(N__14492));
    InMux I__3370 (
            .O(N__14549),
            .I(N__14492));
    InMux I__3369 (
            .O(N__14548),
            .I(N__14489));
    InMux I__3368 (
            .O(N__14547),
            .I(N__14486));
    InMux I__3367 (
            .O(N__14546),
            .I(N__14483));
    LocalMux I__3366 (
            .O(N__14543),
            .I(N__14480));
    LocalMux I__3365 (
            .O(N__14540),
            .I(N__14477));
    LocalMux I__3364 (
            .O(N__14537),
            .I(N__14474));
    LocalMux I__3363 (
            .O(N__14530),
            .I(N__14471));
    LocalMux I__3362 (
            .O(N__14527),
            .I(N__14468));
    LocalMux I__3361 (
            .O(N__14522),
            .I(N__14465));
    LocalMux I__3360 (
            .O(N__14517),
            .I(N__14462));
    LocalMux I__3359 (
            .O(N__14514),
            .I(N__14457));
    LocalMux I__3358 (
            .O(N__14511),
            .I(N__14453));
    LocalMux I__3357 (
            .O(N__14508),
            .I(N__14447));
    LocalMux I__3356 (
            .O(N__14505),
            .I(N__14444));
    LocalMux I__3355 (
            .O(N__14502),
            .I(N__14440));
    LocalMux I__3354 (
            .O(N__14497),
            .I(N__14437));
    LocalMux I__3353 (
            .O(N__14492),
            .I(N__14432));
    LocalMux I__3352 (
            .O(N__14489),
            .I(N__14429));
    LocalMux I__3351 (
            .O(N__14486),
            .I(N__14425));
    LocalMux I__3350 (
            .O(N__14483),
            .I(N__14422));
    Glb2LocalMux I__3349 (
            .O(N__14480),
            .I(N__14364));
    Glb2LocalMux I__3348 (
            .O(N__14477),
            .I(N__14364));
    Glb2LocalMux I__3347 (
            .O(N__14474),
            .I(N__14364));
    Glb2LocalMux I__3346 (
            .O(N__14471),
            .I(N__14364));
    Glb2LocalMux I__3345 (
            .O(N__14468),
            .I(N__14364));
    Glb2LocalMux I__3344 (
            .O(N__14465),
            .I(N__14364));
    Glb2LocalMux I__3343 (
            .O(N__14462),
            .I(N__14364));
    CEMux I__3342 (
            .O(N__14461),
            .I(N__14364));
    CEMux I__3341 (
            .O(N__14460),
            .I(N__14364));
    Glb2LocalMux I__3340 (
            .O(N__14457),
            .I(N__14364));
    CEMux I__3339 (
            .O(N__14456),
            .I(N__14364));
    Glb2LocalMux I__3338 (
            .O(N__14453),
            .I(N__14364));
    CEMux I__3337 (
            .O(N__14452),
            .I(N__14364));
    CEMux I__3336 (
            .O(N__14451),
            .I(N__14364));
    CEMux I__3335 (
            .O(N__14450),
            .I(N__14364));
    Glb2LocalMux I__3334 (
            .O(N__14447),
            .I(N__14364));
    Glb2LocalMux I__3333 (
            .O(N__14444),
            .I(N__14364));
    CEMux I__3332 (
            .O(N__14443),
            .I(N__14364));
    Glb2LocalMux I__3331 (
            .O(N__14440),
            .I(N__14364));
    Glb2LocalMux I__3330 (
            .O(N__14437),
            .I(N__14364));
    CEMux I__3329 (
            .O(N__14436),
            .I(N__14364));
    CEMux I__3328 (
            .O(N__14435),
            .I(N__14364));
    Glb2LocalMux I__3327 (
            .O(N__14432),
            .I(N__14364));
    Glb2LocalMux I__3326 (
            .O(N__14429),
            .I(N__14364));
    CEMux I__3325 (
            .O(N__14428),
            .I(N__14364));
    Glb2LocalMux I__3324 (
            .O(N__14425),
            .I(N__14364));
    Glb2LocalMux I__3323 (
            .O(N__14422),
            .I(N__14364));
    CEMux I__3322 (
            .O(N__14421),
            .I(N__14364));
    GlobalMux I__3321 (
            .O(N__14364),
            .I(N__14361));
    gio2CtrlBuf I__3320 (
            .O(N__14361),
            .I(wPllLocked_g));
    InMux I__3319 (
            .O(N__14358),
            .I(N__14353));
    InMux I__3318 (
            .O(N__14357),
            .I(N__14348));
    InMux I__3317 (
            .O(N__14356),
            .I(N__14348));
    LocalMux I__3316 (
            .O(N__14353),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2 ));
    LocalMux I__3315 (
            .O(N__14348),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2 ));
    CascadeMux I__3314 (
            .O(N__14343),
            .I(\fifo_inst.ftdi_output_inst.N_87_cascade_ ));
    InMux I__3313 (
            .O(N__14340),
            .I(N__14337));
    LocalMux I__3312 (
            .O(N__14337),
            .I(N__14333));
    InMux I__3311 (
            .O(N__14336),
            .I(N__14330));
    Odrv4 I__3310 (
            .O(N__14333),
            .I(\fifo_inst.ftdi_output_inst.N_77_0 ));
    LocalMux I__3309 (
            .O(N__14330),
            .I(\fifo_inst.ftdi_output_inst.N_77_0 ));
    InMux I__3308 (
            .O(N__14325),
            .I(N__14315));
    InMux I__3307 (
            .O(N__14324),
            .I(N__14315));
    InMux I__3306 (
            .O(N__14323),
            .I(N__14315));
    InMux I__3305 (
            .O(N__14322),
            .I(N__14312));
    LocalMux I__3304 (
            .O(N__14315),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0 ));
    LocalMux I__3303 (
            .O(N__14312),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0 ));
    InMux I__3302 (
            .O(N__14307),
            .I(N__14304));
    LocalMux I__3301 (
            .O(N__14304),
            .I(N__14301));
    Span4Mux_v I__3300 (
            .O(N__14301),
            .I(N__14298));
    Sp12to4 I__3299 (
            .O(N__14298),
            .I(N__14295));
    Span12Mux_s6_h I__3298 (
            .O(N__14295),
            .I(N__14292));
    Span12Mux_v I__3297 (
            .O(N__14292),
            .I(N__14289));
    Odrv12 I__3296 (
            .O(N__14289),
            .I(ioFifoData_in_7));
    CascadeMux I__3295 (
            .O(N__14286),
            .I(N__14283));
    InMux I__3294 (
            .O(N__14283),
            .I(N__14280));
    LocalMux I__3293 (
            .O(N__14280),
            .I(N__14277));
    Span4Mux_v I__3292 (
            .O(N__14277),
            .I(N__14274));
    Span4Mux_h I__3291 (
            .O(N__14274),
            .I(N__14271));
    Odrv4 I__3290 (
            .O(N__14271),
            .I(wRxFifoData_7));
    CEMux I__3289 (
            .O(N__14268),
            .I(N__14263));
    CEMux I__3288 (
            .O(N__14267),
            .I(N__14260));
    CEMux I__3287 (
            .O(N__14266),
            .I(N__14257));
    LocalMux I__3286 (
            .O(N__14263),
            .I(N__14254));
    LocalMux I__3285 (
            .O(N__14260),
            .I(N__14251));
    LocalMux I__3284 (
            .O(N__14257),
            .I(N__14248));
    Span4Mux_h I__3283 (
            .O(N__14254),
            .I(N__14245));
    Span4Mux_h I__3282 (
            .O(N__14251),
            .I(N__14240));
    Span4Mux_h I__3281 (
            .O(N__14248),
            .I(N__14240));
    Odrv4 I__3280 (
            .O(N__14245),
            .I(\fifo_inst.ftdi_output_inst.rFifoState_0_1 ));
    Odrv4 I__3279 (
            .O(N__14240),
            .I(\fifo_inst.ftdi_output_inst.rFifoState_0_1 ));
    CascadeMux I__3278 (
            .O(N__14235),
            .I(\fifo_inst.ftdi_output_inst.N_77_0_cascade_ ));
    IoInMux I__3277 (
            .O(N__14232),
            .I(N__14229));
    LocalMux I__3276 (
            .O(N__14229),
            .I(N__14226));
    IoSpan4Mux I__3275 (
            .O(N__14226),
            .I(N__14222));
    IoInMux I__3274 (
            .O(N__14225),
            .I(N__14219));
    Span4Mux_s2_v I__3273 (
            .O(N__14222),
            .I(N__14216));
    LocalMux I__3272 (
            .O(N__14219),
            .I(N__14212));
    Span4Mux_h I__3271 (
            .O(N__14216),
            .I(N__14209));
    InMux I__3270 (
            .O(N__14215),
            .I(N__14206));
    Span12Mux_s11_v I__3269 (
            .O(N__14212),
            .I(N__14203));
    Span4Mux_h I__3268 (
            .O(N__14209),
            .I(N__14198));
    LocalMux I__3267 (
            .O(N__14206),
            .I(N__14198));
    Span12Mux_v I__3266 (
            .O(N__14203),
            .I(N__14194));
    Span4Mux_h I__3265 (
            .O(N__14198),
            .I(N__14191));
    InMux I__3264 (
            .O(N__14197),
            .I(N__14188));
    Odrv12 I__3263 (
            .O(N__14194),
            .I(P1A4_c));
    Odrv4 I__3262 (
            .O(N__14191),
            .I(P1A4_c));
    LocalMux I__3261 (
            .O(N__14188),
            .I(P1A4_c));
    CascadeMux I__3260 (
            .O(N__14181),
            .I(\fifo_inst.ftdi_output_inst.oPacketRead_1_sqmuxa_1_cascade_ ));
    CascadeMux I__3259 (
            .O(N__14178),
            .I(N__14175));
    InMux I__3258 (
            .O(N__14175),
            .I(N__14169));
    InMux I__3257 (
            .O(N__14174),
            .I(N__14162));
    InMux I__3256 (
            .O(N__14173),
            .I(N__14162));
    InMux I__3255 (
            .O(N__14172),
            .I(N__14162));
    LocalMux I__3254 (
            .O(N__14169),
            .I(\fifo_inst.wRamRdAddr_0 ));
    LocalMux I__3253 (
            .O(N__14162),
            .I(\fifo_inst.wRamRdAddr_0 ));
    CascadeMux I__3252 (
            .O(N__14157),
            .I(N__14153));
    CascadeMux I__3251 (
            .O(N__14156),
            .I(N__14150));
    InMux I__3250 (
            .O(N__14153),
            .I(N__14146));
    InMux I__3249 (
            .O(N__14150),
            .I(N__14141));
    InMux I__3248 (
            .O(N__14149),
            .I(N__14141));
    LocalMux I__3247 (
            .O(N__14146),
            .I(\fifo_inst.wRamRdAddr_1 ));
    LocalMux I__3246 (
            .O(N__14141),
            .I(\fifo_inst.wRamRdAddr_1 ));
    InMux I__3245 (
            .O(N__14136),
            .I(N__14133));
    LocalMux I__3244 (
            .O(N__14133),
            .I(\fifo_inst.ftdi_output_inst.oPacketRead_1_sqmuxa_1 ));
    CascadeMux I__3243 (
            .O(N__14130),
            .I(N__14127));
    InMux I__3242 (
            .O(N__14127),
            .I(N__14123));
    InMux I__3241 (
            .O(N__14126),
            .I(N__14120));
    LocalMux I__3240 (
            .O(N__14123),
            .I(\fifo_inst.wRamRdAddr_2 ));
    LocalMux I__3239 (
            .O(N__14120),
            .I(\fifo_inst.wRamRdAddr_2 ));
    InMux I__3238 (
            .O(N__14115),
            .I(N__14110));
    InMux I__3237 (
            .O(N__14114),
            .I(N__14105));
    InMux I__3236 (
            .O(N__14113),
            .I(N__14105));
    LocalMux I__3235 (
            .O(N__14110),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_3 ));
    LocalMux I__3234 (
            .O(N__14105),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_3 ));
    CascadeMux I__3233 (
            .O(N__14100),
            .I(N__14097));
    InMux I__3232 (
            .O(N__14097),
            .I(N__14094));
    LocalMux I__3231 (
            .O(N__14094),
            .I(N__14091));
    Odrv4 I__3230 (
            .O(N__14091),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_6 ));
    InMux I__3229 (
            .O(N__14088),
            .I(N__14083));
    InMux I__3228 (
            .O(N__14087),
            .I(N__14080));
    InMux I__3227 (
            .O(N__14086),
            .I(N__14077));
    LocalMux I__3226 (
            .O(N__14083),
            .I(N__14074));
    LocalMux I__3225 (
            .O(N__14080),
            .I(N__14071));
    LocalMux I__3224 (
            .O(N__14077),
            .I(N__14068));
    Span4Mux_v I__3223 (
            .O(N__14074),
            .I(N__14063));
    Span4Mux_h I__3222 (
            .O(N__14071),
            .I(N__14060));
    Span4Mux_h I__3221 (
            .O(N__14068),
            .I(N__14057));
    InMux I__3220 (
            .O(N__14067),
            .I(N__14054));
    InMux I__3219 (
            .O(N__14066),
            .I(N__14051));
    Odrv4 I__3218 (
            .O(N__14063),
            .I(\DUT.wRxByte_7 ));
    Odrv4 I__3217 (
            .O(N__14060),
            .I(\DUT.wRxByte_7 ));
    Odrv4 I__3216 (
            .O(N__14057),
            .I(\DUT.wRxByte_7 ));
    LocalMux I__3215 (
            .O(N__14054),
            .I(\DUT.wRxByte_7 ));
    LocalMux I__3214 (
            .O(N__14051),
            .I(\DUT.wRxByte_7 ));
    InMux I__3213 (
            .O(N__14040),
            .I(N__14037));
    LocalMux I__3212 (
            .O(N__14037),
            .I(N__14034));
    Span4Mux_h I__3211 (
            .O(N__14034),
            .I(N__14031));
    Odrv4 I__3210 (
            .O(N__14031),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_7 ));
    CEMux I__3209 (
            .O(N__14028),
            .I(N__14025));
    LocalMux I__3208 (
            .O(N__14025),
            .I(\DUT.fifo_rx_inst.rFifoData_awe1 ));
    InMux I__3207 (
            .O(N__14022),
            .I(N__14019));
    LocalMux I__3206 (
            .O(N__14019),
            .I(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0 ));
    CascadeMux I__3205 (
            .O(N__14016),
            .I(N__14012));
    CascadeMux I__3204 (
            .O(N__14015),
            .I(N__14008));
    InMux I__3203 (
            .O(N__14012),
            .I(N__14002));
    InMux I__3202 (
            .O(N__14011),
            .I(N__13991));
    InMux I__3201 (
            .O(N__14008),
            .I(N__13991));
    InMux I__3200 (
            .O(N__14007),
            .I(N__13991));
    InMux I__3199 (
            .O(N__14006),
            .I(N__13991));
    InMux I__3198 (
            .O(N__14005),
            .I(N__13991));
    LocalMux I__3197 (
            .O(N__14002),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_0 ));
    LocalMux I__3196 (
            .O(N__13991),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_0 ));
    CascadeMux I__3195 (
            .O(N__13986),
            .I(N__13983));
    InMux I__3194 (
            .O(N__13983),
            .I(N__13980));
    LocalMux I__3193 (
            .O(N__13980),
            .I(\DUT.fifo_rx_inst.rFifoCount_RNIPTFQ1Z0Z_1 ));
    CascadeMux I__3192 (
            .O(N__13977),
            .I(N__13972));
    CascadeMux I__3191 (
            .O(N__13976),
            .I(N__13969));
    InMux I__3190 (
            .O(N__13975),
            .I(N__13965));
    InMux I__3189 (
            .O(N__13972),
            .I(N__13958));
    InMux I__3188 (
            .O(N__13969),
            .I(N__13958));
    InMux I__3187 (
            .O(N__13968),
            .I(N__13958));
    LocalMux I__3186 (
            .O(N__13965),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_1 ));
    LocalMux I__3185 (
            .O(N__13958),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_1 ));
    InMux I__3184 (
            .O(N__13953),
            .I(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0 ));
    InMux I__3183 (
            .O(N__13950),
            .I(N__13944));
    InMux I__3182 (
            .O(N__13949),
            .I(N__13937));
    InMux I__3181 (
            .O(N__13948),
            .I(N__13937));
    InMux I__3180 (
            .O(N__13947),
            .I(N__13937));
    LocalMux I__3179 (
            .O(N__13944),
            .I(\DUT.fifo_rx_inst.N_4_0 ));
    LocalMux I__3178 (
            .O(N__13937),
            .I(\DUT.fifo_rx_inst.N_4_0 ));
    CascadeMux I__3177 (
            .O(N__13932),
            .I(N__13929));
    InMux I__3176 (
            .O(N__13929),
            .I(N__13921));
    InMux I__3175 (
            .O(N__13928),
            .I(N__13910));
    InMux I__3174 (
            .O(N__13927),
            .I(N__13910));
    InMux I__3173 (
            .O(N__13926),
            .I(N__13910));
    InMux I__3172 (
            .O(N__13925),
            .I(N__13910));
    InMux I__3171 (
            .O(N__13924),
            .I(N__13910));
    LocalMux I__3170 (
            .O(N__13921),
            .I(rRxReadZ0));
    LocalMux I__3169 (
            .O(N__13910),
            .I(rRxReadZ0));
    InMux I__3168 (
            .O(N__13905),
            .I(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1 ));
    InMux I__3167 (
            .O(N__13902),
            .I(N__13898));
    InMux I__3166 (
            .O(N__13901),
            .I(N__13891));
    LocalMux I__3165 (
            .O(N__13898),
            .I(N__13888));
    InMux I__3164 (
            .O(N__13897),
            .I(N__13879));
    InMux I__3163 (
            .O(N__13896),
            .I(N__13879));
    InMux I__3162 (
            .O(N__13895),
            .I(N__13879));
    InMux I__3161 (
            .O(N__13894),
            .I(N__13879));
    LocalMux I__3160 (
            .O(N__13891),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ));
    Odrv12 I__3159 (
            .O(N__13888),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ));
    LocalMux I__3158 (
            .O(N__13879),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ));
    IoInMux I__3157 (
            .O(N__13872),
            .I(N__13869));
    LocalMux I__3156 (
            .O(N__13869),
            .I(N__13866));
    Span4Mux_s2_v I__3155 (
            .O(N__13866),
            .I(N__13863));
    Odrv4 I__3154 (
            .O(N__13863),
            .I(N_1261_i));
    InMux I__3153 (
            .O(N__13860),
            .I(N__13857));
    LocalMux I__3152 (
            .O(N__13857),
            .I(N__13854));
    Odrv4 I__3151 (
            .O(N__13854),
            .I(oTx_n_rep4_ess));
    InMux I__3150 (
            .O(N__13851),
            .I(N__13848));
    LocalMux I__3149 (
            .O(N__13848),
            .I(N__13845));
    Span4Mux_s1_v I__3148 (
            .O(N__13845),
            .I(N__13842));
    Span4Mux_v I__3147 (
            .O(N__13842),
            .I(N__13839));
    Odrv4 I__3146 (
            .O(N__13839),
            .I(oTx_n_rep1_ess));
    InMux I__3145 (
            .O(N__13836),
            .I(N__13833));
    LocalMux I__3144 (
            .O(N__13833),
            .I(N__13830));
    Span4Mux_h I__3143 (
            .O(N__13830),
            .I(N__13827));
    Span4Mux_v I__3142 (
            .O(N__13827),
            .I(N__13824));
    Odrv4 I__3141 (
            .O(N__13824),
            .I(oTx_n_rep0_ess));
    CascadeMux I__3140 (
            .O(N__13821),
            .I(N__13818));
    InMux I__3139 (
            .O(N__13818),
            .I(N__13802));
    InMux I__3138 (
            .O(N__13817),
            .I(N__13802));
    InMux I__3137 (
            .O(N__13816),
            .I(N__13795));
    InMux I__3136 (
            .O(N__13815),
            .I(N__13795));
    InMux I__3135 (
            .O(N__13814),
            .I(N__13795));
    InMux I__3134 (
            .O(N__13813),
            .I(N__13792));
    InMux I__3133 (
            .O(N__13812),
            .I(N__13785));
    InMux I__3132 (
            .O(N__13811),
            .I(N__13785));
    InMux I__3131 (
            .O(N__13810),
            .I(N__13785));
    InMux I__3130 (
            .O(N__13809),
            .I(N__13778));
    InMux I__3129 (
            .O(N__13808),
            .I(N__13778));
    InMux I__3128 (
            .O(N__13807),
            .I(N__13778));
    LocalMux I__3127 (
            .O(N__13802),
            .I(N__13773));
    LocalMux I__3126 (
            .O(N__13795),
            .I(N__13773));
    LocalMux I__3125 (
            .O(N__13792),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__3124 (
            .O(N__13785),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__3123 (
            .O(N__13778),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    Odrv4 I__3122 (
            .O(N__13773),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    InMux I__3121 (
            .O(N__13764),
            .I(N__13761));
    LocalMux I__3120 (
            .O(N__13761),
            .I(N__13758));
    Span4Mux_v I__3119 (
            .O(N__13758),
            .I(N__13755));
    Odrv4 I__3118 (
            .O(N__13755),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_2 ));
    InMux I__3117 (
            .O(N__13752),
            .I(N__13749));
    LocalMux I__3116 (
            .O(N__13749),
            .I(N__13746));
    Odrv4 I__3115 (
            .O(N__13746),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_2 ));
    CascadeMux I__3114 (
            .O(N__13743),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2_cascade_ ));
    CascadeMux I__3113 (
            .O(N__13740),
            .I(N__13726));
    CascadeMux I__3112 (
            .O(N__13739),
            .I(N__13723));
    CascadeMux I__3111 (
            .O(N__13738),
            .I(N__13717));
    CascadeMux I__3110 (
            .O(N__13737),
            .I(N__13713));
    InMux I__3109 (
            .O(N__13736),
            .I(N__13710));
    CascadeMux I__3108 (
            .O(N__13735),
            .I(N__13705));
    CascadeMux I__3107 (
            .O(N__13734),
            .I(N__13701));
    InMux I__3106 (
            .O(N__13733),
            .I(N__13697));
    InMux I__3105 (
            .O(N__13732),
            .I(N__13684));
    InMux I__3104 (
            .O(N__13731),
            .I(N__13684));
    InMux I__3103 (
            .O(N__13730),
            .I(N__13684));
    InMux I__3102 (
            .O(N__13729),
            .I(N__13684));
    InMux I__3101 (
            .O(N__13726),
            .I(N__13684));
    InMux I__3100 (
            .O(N__13723),
            .I(N__13684));
    InMux I__3099 (
            .O(N__13722),
            .I(N__13671));
    InMux I__3098 (
            .O(N__13721),
            .I(N__13671));
    InMux I__3097 (
            .O(N__13720),
            .I(N__13671));
    InMux I__3096 (
            .O(N__13717),
            .I(N__13671));
    InMux I__3095 (
            .O(N__13716),
            .I(N__13671));
    InMux I__3094 (
            .O(N__13713),
            .I(N__13671));
    LocalMux I__3093 (
            .O(N__13710),
            .I(N__13668));
    InMux I__3092 (
            .O(N__13709),
            .I(N__13661));
    InMux I__3091 (
            .O(N__13708),
            .I(N__13661));
    InMux I__3090 (
            .O(N__13705),
            .I(N__13661));
    InMux I__3089 (
            .O(N__13704),
            .I(N__13654));
    InMux I__3088 (
            .O(N__13701),
            .I(N__13654));
    InMux I__3087 (
            .O(N__13700),
            .I(N__13654));
    LocalMux I__3086 (
            .O(N__13697),
            .I(N__13647));
    LocalMux I__3085 (
            .O(N__13684),
            .I(N__13647));
    LocalMux I__3084 (
            .O(N__13671),
            .I(N__13647));
    Odrv4 I__3083 (
            .O(N__13668),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__3082 (
            .O(N__13661),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__3081 (
            .O(N__13654),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    Odrv4 I__3080 (
            .O(N__13647),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    InMux I__3079 (
            .O(N__13638),
            .I(N__13635));
    LocalMux I__3078 (
            .O(N__13635),
            .I(\DUT.fifo_rx_inst.rFifoDatarx_2 ));
    InMux I__3077 (
            .O(N__13632),
            .I(N__13627));
    InMux I__3076 (
            .O(N__13631),
            .I(N__13624));
    InMux I__3075 (
            .O(N__13630),
            .I(N__13621));
    LocalMux I__3074 (
            .O(N__13627),
            .I(N__13616));
    LocalMux I__3073 (
            .O(N__13624),
            .I(N__13616));
    LocalMux I__3072 (
            .O(N__13621),
            .I(N__13613));
    Span4Mux_v I__3071 (
            .O(N__13616),
            .I(N__13609));
    Span4Mux_h I__3070 (
            .O(N__13613),
            .I(N__13606));
    InMux I__3069 (
            .O(N__13612),
            .I(N__13603));
    Odrv4 I__3068 (
            .O(N__13609),
            .I(\DUT.wRxByte_0 ));
    Odrv4 I__3067 (
            .O(N__13606),
            .I(\DUT.wRxByte_0 ));
    LocalMux I__3066 (
            .O(N__13603),
            .I(\DUT.wRxByte_0 ));
    InMux I__3065 (
            .O(N__13596),
            .I(N__13593));
    LocalMux I__3064 (
            .O(N__13593),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_0 ));
    InMux I__3063 (
            .O(N__13590),
            .I(N__13585));
    InMux I__3062 (
            .O(N__13589),
            .I(N__13582));
    InMux I__3061 (
            .O(N__13588),
            .I(N__13579));
    LocalMux I__3060 (
            .O(N__13585),
            .I(N__13574));
    LocalMux I__3059 (
            .O(N__13582),
            .I(N__13574));
    LocalMux I__3058 (
            .O(N__13579),
            .I(N__13571));
    Span4Mux_v I__3057 (
            .O(N__13574),
            .I(N__13566));
    Span4Mux_h I__3056 (
            .O(N__13571),
            .I(N__13563));
    InMux I__3055 (
            .O(N__13570),
            .I(N__13560));
    InMux I__3054 (
            .O(N__13569),
            .I(N__13557));
    Odrv4 I__3053 (
            .O(N__13566),
            .I(\DUT.wRxByte_1 ));
    Odrv4 I__3052 (
            .O(N__13563),
            .I(\DUT.wRxByte_1 ));
    LocalMux I__3051 (
            .O(N__13560),
            .I(\DUT.wRxByte_1 ));
    LocalMux I__3050 (
            .O(N__13557),
            .I(\DUT.wRxByte_1 ));
    InMux I__3049 (
            .O(N__13548),
            .I(N__13545));
    LocalMux I__3048 (
            .O(N__13545),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_1 ));
    InMux I__3047 (
            .O(N__13542),
            .I(N__13539));
    LocalMux I__3046 (
            .O(N__13539),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_2 ));
    InMux I__3045 (
            .O(N__13536),
            .I(N__13531));
    InMux I__3044 (
            .O(N__13535),
            .I(N__13528));
    InMux I__3043 (
            .O(N__13534),
            .I(N__13525));
    LocalMux I__3042 (
            .O(N__13531),
            .I(N__13522));
    LocalMux I__3041 (
            .O(N__13528),
            .I(N__13517));
    LocalMux I__3040 (
            .O(N__13525),
            .I(N__13517));
    Span4Mux_h I__3039 (
            .O(N__13522),
            .I(N__13512));
    Span4Mux_v I__3038 (
            .O(N__13517),
            .I(N__13509));
    InMux I__3037 (
            .O(N__13516),
            .I(N__13506));
    InMux I__3036 (
            .O(N__13515),
            .I(N__13503));
    Odrv4 I__3035 (
            .O(N__13512),
            .I(\DUT.wRxByte_3 ));
    Odrv4 I__3034 (
            .O(N__13509),
            .I(\DUT.wRxByte_3 ));
    LocalMux I__3033 (
            .O(N__13506),
            .I(\DUT.wRxByte_3 ));
    LocalMux I__3032 (
            .O(N__13503),
            .I(\DUT.wRxByte_3 ));
    InMux I__3031 (
            .O(N__13494),
            .I(N__13491));
    LocalMux I__3030 (
            .O(N__13491),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_3 ));
    InMux I__3029 (
            .O(N__13488),
            .I(N__13484));
    InMux I__3028 (
            .O(N__13487),
            .I(N__13481));
    LocalMux I__3027 (
            .O(N__13484),
            .I(N__13475));
    LocalMux I__3026 (
            .O(N__13481),
            .I(N__13475));
    InMux I__3025 (
            .O(N__13480),
            .I(N__13472));
    Span4Mux_v I__3024 (
            .O(N__13475),
            .I(N__13469));
    LocalMux I__3023 (
            .O(N__13472),
            .I(N__13464));
    Sp12to4 I__3022 (
            .O(N__13469),
            .I(N__13461));
    InMux I__3021 (
            .O(N__13468),
            .I(N__13458));
    InMux I__3020 (
            .O(N__13467),
            .I(N__13455));
    Odrv4 I__3019 (
            .O(N__13464),
            .I(\DUT.wRxByte_4 ));
    Odrv12 I__3018 (
            .O(N__13461),
            .I(\DUT.wRxByte_4 ));
    LocalMux I__3017 (
            .O(N__13458),
            .I(\DUT.wRxByte_4 ));
    LocalMux I__3016 (
            .O(N__13455),
            .I(\DUT.wRxByte_4 ));
    InMux I__3015 (
            .O(N__13446),
            .I(N__13443));
    LocalMux I__3014 (
            .O(N__13443),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_4 ));
    InMux I__3013 (
            .O(N__13440),
            .I(N__13437));
    LocalMux I__3012 (
            .O(N__13437),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_5 ));
    InMux I__3011 (
            .O(N__13434),
            .I(N__13430));
    InMux I__3010 (
            .O(N__13433),
            .I(N__13427));
    LocalMux I__3009 (
            .O(N__13430),
            .I(N__13423));
    LocalMux I__3008 (
            .O(N__13427),
            .I(N__13420));
    InMux I__3007 (
            .O(N__13426),
            .I(N__13417));
    Span4Mux_v I__3006 (
            .O(N__13423),
            .I(N__13412));
    Span4Mux_h I__3005 (
            .O(N__13420),
            .I(N__13409));
    LocalMux I__3004 (
            .O(N__13417),
            .I(N__13406));
    InMux I__3003 (
            .O(N__13416),
            .I(N__13403));
    InMux I__3002 (
            .O(N__13415),
            .I(N__13400));
    Odrv4 I__3001 (
            .O(N__13412),
            .I(\DUT.wRxByte_6 ));
    Odrv4 I__3000 (
            .O(N__13409),
            .I(\DUT.wRxByte_6 ));
    Odrv4 I__2999 (
            .O(N__13406),
            .I(\DUT.wRxByte_6 ));
    LocalMux I__2998 (
            .O(N__13403),
            .I(\DUT.wRxByte_6 ));
    LocalMux I__2997 (
            .O(N__13400),
            .I(\DUT.wRxByte_6 ));
    InMux I__2996 (
            .O(N__13389),
            .I(N__13386));
    LocalMux I__2995 (
            .O(N__13386),
            .I(\DUT.fifo_rx_inst.rFifoDatarx_3 ));
    CascadeMux I__2994 (
            .O(N__13383),
            .I(N__13380));
    InMux I__2993 (
            .O(N__13380),
            .I(N__13377));
    LocalMux I__2992 (
            .O(N__13377),
            .I(N__13374));
    Odrv4 I__2991 (
            .O(N__13374),
            .I(wRxFifoData_3));
    InMux I__2990 (
            .O(N__13371),
            .I(N__13368));
    LocalMux I__2989 (
            .O(N__13368),
            .I(N__13362));
    InMux I__2988 (
            .O(N__13367),
            .I(N__13359));
    InMux I__2987 (
            .O(N__13366),
            .I(N__13356));
    InMux I__2986 (
            .O(N__13365),
            .I(N__13353));
    Span4Mux_h I__2985 (
            .O(N__13362),
            .I(N__13344));
    LocalMux I__2984 (
            .O(N__13359),
            .I(N__13344));
    LocalMux I__2983 (
            .O(N__13356),
            .I(N__13344));
    LocalMux I__2982 (
            .O(N__13353),
            .I(N__13344));
    Span4Mux_v I__2981 (
            .O(N__13344),
            .I(N__13341));
    Odrv4 I__2980 (
            .O(N__13341),
            .I(rTxByteZ0Z_3));
    InMux I__2979 (
            .O(N__13338),
            .I(N__13314));
    InMux I__2978 (
            .O(N__13337),
            .I(N__13314));
    InMux I__2977 (
            .O(N__13336),
            .I(N__13314));
    InMux I__2976 (
            .O(N__13335),
            .I(N__13314));
    InMux I__2975 (
            .O(N__13334),
            .I(N__13314));
    InMux I__2974 (
            .O(N__13333),
            .I(N__13314));
    InMux I__2973 (
            .O(N__13332),
            .I(N__13314));
    InMux I__2972 (
            .O(N__13331),
            .I(N__13314));
    LocalMux I__2971 (
            .O(N__13314),
            .I(\DUT.fifo_rx_inst.rFifoDataror_0 ));
    CascadeMux I__2970 (
            .O(N__13311),
            .I(N__13308));
    InMux I__2969 (
            .O(N__13308),
            .I(N__13305));
    LocalMux I__2968 (
            .O(N__13305),
            .I(N__13302));
    Odrv12 I__2967 (
            .O(N__13302),
            .I(wRxFifoData_4));
    InMux I__2966 (
            .O(N__13299),
            .I(N__13296));
    LocalMux I__2965 (
            .O(N__13296),
            .I(\DUT.fifo_rx_inst.rFifoDatarx_4 ));
    InMux I__2964 (
            .O(N__13293),
            .I(N__13289));
    InMux I__2963 (
            .O(N__13292),
            .I(N__13286));
    LocalMux I__2962 (
            .O(N__13289),
            .I(N__13282));
    LocalMux I__2961 (
            .O(N__13286),
            .I(N__13279));
    InMux I__2960 (
            .O(N__13285),
            .I(N__13276));
    Span4Mux_v I__2959 (
            .O(N__13282),
            .I(N__13268));
    Span4Mux_h I__2958 (
            .O(N__13279),
            .I(N__13268));
    LocalMux I__2957 (
            .O(N__13276),
            .I(N__13268));
    InMux I__2956 (
            .O(N__13275),
            .I(N__13265));
    Sp12to4 I__2955 (
            .O(N__13268),
            .I(N__13260));
    LocalMux I__2954 (
            .O(N__13265),
            .I(N__13260));
    Odrv12 I__2953 (
            .O(N__13260),
            .I(rTxByteZ0Z_4));
    CEMux I__2952 (
            .O(N__13257),
            .I(N__13254));
    LocalMux I__2951 (
            .O(N__13254),
            .I(N__13251));
    Span4Mux_v I__2950 (
            .O(N__13251),
            .I(N__13248));
    Odrv4 I__2949 (
            .O(N__13248),
            .I(rTxByte_1_sqmuxa_i_0));
    InMux I__2948 (
            .O(N__13245),
            .I(N__13242));
    LocalMux I__2947 (
            .O(N__13242),
            .I(N__13239));
    Odrv4 I__2946 (
            .O(N__13239),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_0 ));
    InMux I__2945 (
            .O(N__13236),
            .I(N__13233));
    LocalMux I__2944 (
            .O(N__13233),
            .I(N__13230));
    Span4Mux_h I__2943 (
            .O(N__13230),
            .I(N__13227));
    Odrv4 I__2942 (
            .O(N__13227),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_0 ));
    CascadeMux I__2941 (
            .O(N__13224),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ));
    InMux I__2940 (
            .O(N__13221),
            .I(N__13218));
    LocalMux I__2939 (
            .O(N__13218),
            .I(\DUT.fifo_rx_inst.rFifoDatarx_0 ));
    InMux I__2938 (
            .O(N__13215),
            .I(N__13212));
    LocalMux I__2937 (
            .O(N__13212),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_0 ));
    InMux I__2936 (
            .O(N__13209),
            .I(N__13206));
    LocalMux I__2935 (
            .O(N__13206),
            .I(N__13203));
    Span4Mux_h I__2934 (
            .O(N__13203),
            .I(N__13200));
    Odrv4 I__2933 (
            .O(N__13200),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_1 ));
    CascadeMux I__2932 (
            .O(N__13197),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1_cascade_ ));
    InMux I__2931 (
            .O(N__13194),
            .I(N__13191));
    LocalMux I__2930 (
            .O(N__13191),
            .I(N__13188));
    Odrv4 I__2929 (
            .O(N__13188),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_1 ));
    InMux I__2928 (
            .O(N__13185),
            .I(N__13182));
    LocalMux I__2927 (
            .O(N__13182),
            .I(\DUT.fifo_rx_inst.rFifoDatarx_1 ));
    CascadeMux I__2926 (
            .O(N__13179),
            .I(N__13176));
    InMux I__2925 (
            .O(N__13176),
            .I(N__13173));
    LocalMux I__2924 (
            .O(N__13173),
            .I(N__13170));
    Odrv4 I__2923 (
            .O(N__13170),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_1 ));
    InMux I__2922 (
            .O(N__13167),
            .I(N__13164));
    LocalMux I__2921 (
            .O(N__13164),
            .I(N__13161));
    Span4Mux_h I__2920 (
            .O(N__13161),
            .I(N__13158));
    Odrv4 I__2919 (
            .O(N__13158),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_5 ));
    InMux I__2918 (
            .O(N__13155),
            .I(N__13152));
    LocalMux I__2917 (
            .O(N__13152),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_6 ));
    InMux I__2916 (
            .O(N__13149),
            .I(N__13146));
    LocalMux I__2915 (
            .O(N__13146),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_7 ));
    CEMux I__2914 (
            .O(N__13143),
            .I(N__13140));
    LocalMux I__2913 (
            .O(N__13140),
            .I(N__13137));
    Span4Mux_v I__2912 (
            .O(N__13137),
            .I(N__13134));
    Odrv4 I__2911 (
            .O(N__13134),
            .I(\DUT.fifo_rx_inst.rFifoData_awe2 ));
    InMux I__2910 (
            .O(N__13131),
            .I(N__13128));
    LocalMux I__2909 (
            .O(N__13128),
            .I(\DUT.fifo_rx_inst.rFifoDatarx_6 ));
    InMux I__2908 (
            .O(N__13125),
            .I(N__13122));
    LocalMux I__2907 (
            .O(N__13122),
            .I(N__13119));
    Odrv12 I__2906 (
            .O(N__13119),
            .I(wRxFifoData_6));
    InMux I__2905 (
            .O(N__13116),
            .I(N__13112));
    InMux I__2904 (
            .O(N__13115),
            .I(N__13109));
    LocalMux I__2903 (
            .O(N__13112),
            .I(N__13105));
    LocalMux I__2902 (
            .O(N__13109),
            .I(N__13101));
    InMux I__2901 (
            .O(N__13108),
            .I(N__13098));
    Span4Mux_h I__2900 (
            .O(N__13105),
            .I(N__13095));
    InMux I__2899 (
            .O(N__13104),
            .I(N__13092));
    Span4Mux_v I__2898 (
            .O(N__13101),
            .I(N__13087));
    LocalMux I__2897 (
            .O(N__13098),
            .I(N__13087));
    Sp12to4 I__2896 (
            .O(N__13095),
            .I(N__13082));
    LocalMux I__2895 (
            .O(N__13092),
            .I(N__13082));
    Odrv4 I__2894 (
            .O(N__13087),
            .I(rTxByteZ0Z_6));
    Odrv12 I__2893 (
            .O(N__13082),
            .I(rTxByteZ0Z_6));
    CascadeMux I__2892 (
            .O(N__13077),
            .I(N__13074));
    InMux I__2891 (
            .O(N__13074),
            .I(N__13071));
    LocalMux I__2890 (
            .O(N__13071),
            .I(N__13068));
    Odrv4 I__2889 (
            .O(N__13068),
            .I(wRxFifoData_5));
    InMux I__2888 (
            .O(N__13065),
            .I(N__13062));
    LocalMux I__2887 (
            .O(N__13062),
            .I(\DUT.fifo_rx_inst.rFifoDatarx_5 ));
    InMux I__2886 (
            .O(N__13059),
            .I(N__13055));
    InMux I__2885 (
            .O(N__13058),
            .I(N__13052));
    LocalMux I__2884 (
            .O(N__13055),
            .I(N__13047));
    LocalMux I__2883 (
            .O(N__13052),
            .I(N__13044));
    InMux I__2882 (
            .O(N__13051),
            .I(N__13041));
    InMux I__2881 (
            .O(N__13050),
            .I(N__13038));
    Span4Mux_v I__2880 (
            .O(N__13047),
            .I(N__13031));
    Span4Mux_h I__2879 (
            .O(N__13044),
            .I(N__13031));
    LocalMux I__2878 (
            .O(N__13041),
            .I(N__13031));
    LocalMux I__2877 (
            .O(N__13038),
            .I(N__13028));
    Odrv4 I__2876 (
            .O(N__13031),
            .I(rTxByteZ0Z_5));
    Odrv12 I__2875 (
            .O(N__13028),
            .I(rTxByteZ0Z_5));
    CascadeMux I__2874 (
            .O(N__13023),
            .I(N__13020));
    InMux I__2873 (
            .O(N__13020),
            .I(N__13017));
    LocalMux I__2872 (
            .O(N__13017),
            .I(N__13014));
    Odrv4 I__2871 (
            .O(N__13014),
            .I(wRxFifoData_0));
    InMux I__2870 (
            .O(N__13011),
            .I(N__13008));
    LocalMux I__2869 (
            .O(N__13008),
            .I(N__13004));
    InMux I__2868 (
            .O(N__13007),
            .I(N__13001));
    Span4Mux_h I__2867 (
            .O(N__13004),
            .I(N__12996));
    LocalMux I__2866 (
            .O(N__13001),
            .I(N__12993));
    InMux I__2865 (
            .O(N__13000),
            .I(N__12990));
    InMux I__2864 (
            .O(N__12999),
            .I(N__12987));
    Span4Mux_v I__2863 (
            .O(N__12996),
            .I(N__12984));
    Span4Mux_v I__2862 (
            .O(N__12993),
            .I(N__12979));
    LocalMux I__2861 (
            .O(N__12990),
            .I(N__12979));
    LocalMux I__2860 (
            .O(N__12987),
            .I(N__12976));
    Odrv4 I__2859 (
            .O(N__12984),
            .I(rTxByteZ0Z_0));
    Odrv4 I__2858 (
            .O(N__12979),
            .I(rTxByteZ0Z_0));
    Odrv12 I__2857 (
            .O(N__12976),
            .I(rTxByteZ0Z_0));
    InMux I__2856 (
            .O(N__12969),
            .I(N__12966));
    LocalMux I__2855 (
            .O(N__12966),
            .I(\DUT.fifo_rx_inst.rFifoDatarx_7 ));
    InMux I__2854 (
            .O(N__12963),
            .I(N__12960));
    LocalMux I__2853 (
            .O(N__12960),
            .I(N__12955));
    InMux I__2852 (
            .O(N__12959),
            .I(N__12952));
    InMux I__2851 (
            .O(N__12958),
            .I(N__12949));
    Span4Mux_h I__2850 (
            .O(N__12955),
            .I(N__12945));
    LocalMux I__2849 (
            .O(N__12952),
            .I(N__12942));
    LocalMux I__2848 (
            .O(N__12949),
            .I(N__12939));
    InMux I__2847 (
            .O(N__12948),
            .I(N__12936));
    Span4Mux_v I__2846 (
            .O(N__12945),
            .I(N__12933));
    Span4Mux_v I__2845 (
            .O(N__12942),
            .I(N__12930));
    Span4Mux_h I__2844 (
            .O(N__12939),
            .I(N__12927));
    LocalMux I__2843 (
            .O(N__12936),
            .I(N__12924));
    Odrv4 I__2842 (
            .O(N__12933),
            .I(rTxByteZ0Z_7));
    Odrv4 I__2841 (
            .O(N__12930),
            .I(rTxByteZ0Z_7));
    Odrv4 I__2840 (
            .O(N__12927),
            .I(rTxByteZ0Z_7));
    Odrv12 I__2839 (
            .O(N__12924),
            .I(rTxByteZ0Z_7));
    CascadeMux I__2838 (
            .O(N__12915),
            .I(N__12912));
    InMux I__2837 (
            .O(N__12912),
            .I(N__12909));
    LocalMux I__2836 (
            .O(N__12909),
            .I(N__12906));
    Odrv4 I__2835 (
            .O(N__12906),
            .I(wRxFifoData_1));
    InMux I__2834 (
            .O(N__12903),
            .I(N__12899));
    InMux I__2833 (
            .O(N__12902),
            .I(N__12896));
    LocalMux I__2832 (
            .O(N__12899),
            .I(N__12891));
    LocalMux I__2831 (
            .O(N__12896),
            .I(N__12888));
    InMux I__2830 (
            .O(N__12895),
            .I(N__12885));
    InMux I__2829 (
            .O(N__12894),
            .I(N__12882));
    Span4Mux_h I__2828 (
            .O(N__12891),
            .I(N__12879));
    Span4Mux_h I__2827 (
            .O(N__12888),
            .I(N__12874));
    LocalMux I__2826 (
            .O(N__12885),
            .I(N__12874));
    LocalMux I__2825 (
            .O(N__12882),
            .I(N__12871));
    Span4Mux_v I__2824 (
            .O(N__12879),
            .I(N__12868));
    Span4Mux_v I__2823 (
            .O(N__12874),
            .I(N__12865));
    Span4Mux_h I__2822 (
            .O(N__12871),
            .I(N__12862));
    Odrv4 I__2821 (
            .O(N__12868),
            .I(rTxByteZ0Z_1));
    Odrv4 I__2820 (
            .O(N__12865),
            .I(rTxByteZ0Z_1));
    Odrv4 I__2819 (
            .O(N__12862),
            .I(rTxByteZ0Z_1));
    CascadeMux I__2818 (
            .O(N__12855),
            .I(N__12852));
    InMux I__2817 (
            .O(N__12852),
            .I(N__12849));
    LocalMux I__2816 (
            .O(N__12849),
            .I(N__12846));
    Odrv4 I__2815 (
            .O(N__12846),
            .I(wRxFifoData_2));
    InMux I__2814 (
            .O(N__12843),
            .I(N__12840));
    LocalMux I__2813 (
            .O(N__12840),
            .I(N__12834));
    InMux I__2812 (
            .O(N__12839),
            .I(N__12831));
    InMux I__2811 (
            .O(N__12838),
            .I(N__12828));
    InMux I__2810 (
            .O(N__12837),
            .I(N__12825));
    Span4Mux_h I__2809 (
            .O(N__12834),
            .I(N__12816));
    LocalMux I__2808 (
            .O(N__12831),
            .I(N__12816));
    LocalMux I__2807 (
            .O(N__12828),
            .I(N__12816));
    LocalMux I__2806 (
            .O(N__12825),
            .I(N__12816));
    Span4Mux_v I__2805 (
            .O(N__12816),
            .I(N__12813));
    Odrv4 I__2804 (
            .O(N__12813),
            .I(rTxByteZ0Z_2));
    InMux I__2803 (
            .O(N__12810),
            .I(N__12807));
    LocalMux I__2802 (
            .O(N__12807),
            .I(N__12804));
    Span12Mux_h I__2801 (
            .O(N__12804),
            .I(N__12801));
    Odrv12 I__2800 (
            .O(N__12801),
            .I(ioFifoData_in_2));
    InMux I__2799 (
            .O(N__12798),
            .I(N__12795));
    LocalMux I__2798 (
            .O(N__12795),
            .I(N__12792));
    Span12Mux_h I__2797 (
            .O(N__12792),
            .I(N__12789));
    Odrv12 I__2796 (
            .O(N__12789),
            .I(ioFifoData_in_0));
    InMux I__2795 (
            .O(N__12786),
            .I(N__12783));
    LocalMux I__2794 (
            .O(N__12783),
            .I(N__12780));
    Sp12to4 I__2793 (
            .O(N__12780),
            .I(N__12777));
    Span12Mux_v I__2792 (
            .O(N__12777),
            .I(N__12774));
    Odrv12 I__2791 (
            .O(N__12774),
            .I(ioFifoData_in_6));
    InMux I__2790 (
            .O(N__12771),
            .I(N__12768));
    LocalMux I__2789 (
            .O(N__12768),
            .I(N__12765));
    Span4Mux_v I__2788 (
            .O(N__12765),
            .I(N__12762));
    Odrv4 I__2787 (
            .O(N__12762),
            .I(ioFifoData_in_4));
    InMux I__2786 (
            .O(N__12759),
            .I(N__12756));
    LocalMux I__2785 (
            .O(N__12756),
            .I(N__12753));
    Span4Mux_v I__2784 (
            .O(N__12753),
            .I(N__12750));
    Odrv4 I__2783 (
            .O(N__12750),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_3 ));
    InMux I__2782 (
            .O(N__12747),
            .I(N__12744));
    LocalMux I__2781 (
            .O(N__12744),
            .I(N__12741));
    Odrv4 I__2780 (
            .O(N__12741),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_4 ));
    InMux I__2779 (
            .O(N__12738),
            .I(N__12735));
    LocalMux I__2778 (
            .O(N__12735),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_2 ));
    InMux I__2777 (
            .O(N__12732),
            .I(N__12729));
    LocalMux I__2776 (
            .O(N__12729),
            .I(N__12726));
    Odrv4 I__2775 (
            .O(N__12726),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_3 ));
    InMux I__2774 (
            .O(N__12723),
            .I(N__12720));
    LocalMux I__2773 (
            .O(N__12720),
            .I(N__12717));
    Span4Mux_h I__2772 (
            .O(N__12717),
            .I(N__12714));
    Odrv4 I__2771 (
            .O(N__12714),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_4 ));
    InMux I__2770 (
            .O(N__12711),
            .I(N__12708));
    LocalMux I__2769 (
            .O(N__12708),
            .I(N__12705));
    Span4Mux_h I__2768 (
            .O(N__12705),
            .I(N__12702));
    Odrv4 I__2767 (
            .O(N__12702),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_5 ));
    InMux I__2766 (
            .O(N__12699),
            .I(N__12696));
    LocalMux I__2765 (
            .O(N__12696),
            .I(N__12693));
    Odrv12 I__2764 (
            .O(N__12693),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_6 ));
    InMux I__2763 (
            .O(N__12690),
            .I(N__12687));
    LocalMux I__2762 (
            .O(N__12687),
            .I(N__12684));
    Span4Mux_h I__2761 (
            .O(N__12684),
            .I(N__12681));
    Odrv4 I__2760 (
            .O(N__12681),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_7 ));
    CEMux I__2759 (
            .O(N__12678),
            .I(N__12675));
    LocalMux I__2758 (
            .O(N__12675),
            .I(N__12672));
    Span4Mux_v I__2757 (
            .O(N__12672),
            .I(N__12668));
    InMux I__2756 (
            .O(N__12671),
            .I(N__12665));
    Span4Mux_h I__2755 (
            .O(N__12668),
            .I(N__12660));
    LocalMux I__2754 (
            .O(N__12665),
            .I(N__12660));
    Span4Mux_h I__2753 (
            .O(N__12660),
            .I(N__12656));
    InMux I__2752 (
            .O(N__12659),
            .I(N__12653));
    Odrv4 I__2751 (
            .O(N__12656),
            .I(\DUT.fifo_tx_inst.rFifoData_awe3 ));
    LocalMux I__2750 (
            .O(N__12653),
            .I(\DUT.fifo_tx_inst.rFifoData_awe3 ));
    InMux I__2749 (
            .O(N__12648),
            .I(N__12645));
    LocalMux I__2748 (
            .O(N__12645),
            .I(N__12642));
    Span4Mux_h I__2747 (
            .O(N__12642),
            .I(N__12639));
    Span4Mux_v I__2746 (
            .O(N__12639),
            .I(N__12636));
    Odrv4 I__2745 (
            .O(N__12636),
            .I(ioFifoData_in_3));
    InMux I__2744 (
            .O(N__12633),
            .I(N__12630));
    LocalMux I__2743 (
            .O(N__12630),
            .I(N__12627));
    Span4Mux_h I__2742 (
            .O(N__12627),
            .I(N__12624));
    Span4Mux_v I__2741 (
            .O(N__12624),
            .I(N__12621));
    Odrv4 I__2740 (
            .O(N__12621),
            .I(ioFifoData_in_1));
    InMux I__2739 (
            .O(N__12618),
            .I(N__12615));
    LocalMux I__2738 (
            .O(N__12615),
            .I(N__12612));
    Odrv12 I__2737 (
            .O(N__12612),
            .I(ioFifoData_in_5));
    CascadeMux I__2736 (
            .O(N__12609),
            .I(N__12605));
    InMux I__2735 (
            .O(N__12608),
            .I(N__12601));
    InMux I__2734 (
            .O(N__12605),
            .I(N__12596));
    InMux I__2733 (
            .O(N__12604),
            .I(N__12596));
    LocalMux I__2732 (
            .O(N__12601),
            .I(N__12593));
    LocalMux I__2731 (
            .O(N__12596),
            .I(N__12589));
    Span4Mux_v I__2730 (
            .O(N__12593),
            .I(N__12586));
    InMux I__2729 (
            .O(N__12592),
            .I(N__12583));
    Span4Mux_h I__2728 (
            .O(N__12589),
            .I(N__12580));
    Odrv4 I__2727 (
            .O(N__12586),
            .I(\DUT.wRcvd ));
    LocalMux I__2726 (
            .O(N__12583),
            .I(\DUT.wRcvd ));
    Odrv4 I__2725 (
            .O(N__12580),
            .I(\DUT.wRcvd ));
    InMux I__2724 (
            .O(N__12573),
            .I(N__12567));
    InMux I__2723 (
            .O(N__12572),
            .I(N__12567));
    LocalMux I__2722 (
            .O(N__12567),
            .I(N__12563));
    CascadeMux I__2721 (
            .O(N__12566),
            .I(N__12560));
    Span4Mux_h I__2720 (
            .O(N__12563),
            .I(N__12557));
    InMux I__2719 (
            .O(N__12560),
            .I(N__12554));
    Odrv4 I__2718 (
            .O(N__12557),
            .I(\DUT.fifo_rx_inst.N_46 ));
    LocalMux I__2717 (
            .O(N__12554),
            .I(\DUT.fifo_rx_inst.N_46 ));
    InMux I__2716 (
            .O(N__12549),
            .I(N__12546));
    LocalMux I__2715 (
            .O(N__12546),
            .I(N__12543));
    Span4Mux_h I__2714 (
            .O(N__12543),
            .I(N__12540));
    Span4Mux_h I__2713 (
            .O(N__12540),
            .I(N__12536));
    InMux I__2712 (
            .O(N__12539),
            .I(N__12533));
    Odrv4 I__2711 (
            .O(N__12536),
            .I(N_69_mux));
    LocalMux I__2710 (
            .O(N__12533),
            .I(N_69_mux));
    CascadeMux I__2709 (
            .O(N__12528),
            .I(N_69_mux_cascade_));
    IoInMux I__2708 (
            .O(N__12525),
            .I(N__12522));
    LocalMux I__2707 (
            .O(N__12522),
            .I(N__12519));
    IoSpan4Mux I__2706 (
            .O(N__12519),
            .I(N__12516));
    Odrv4 I__2705 (
            .O(N__12516),
            .I(N_1258_i));
    IoInMux I__2704 (
            .O(N__12513),
            .I(N__12509));
    IoInMux I__2703 (
            .O(N__12512),
            .I(N__12506));
    LocalMux I__2702 (
            .O(N__12509),
            .I(N__12501));
    LocalMux I__2701 (
            .O(N__12506),
            .I(N__12501));
    Span4Mux_s1_v I__2700 (
            .O(N__12501),
            .I(N__12498));
    Sp12to4 I__2699 (
            .O(N__12498),
            .I(N__12495));
    Span12Mux_s7_h I__2698 (
            .O(N__12495),
            .I(N__12492));
    Span12Mux_v I__2697 (
            .O(N__12492),
            .I(N__12488));
    IoInMux I__2696 (
            .O(N__12491),
            .I(N__12485));
    Span12Mux_v I__2695 (
            .O(N__12488),
            .I(N__12482));
    LocalMux I__2694 (
            .O(N__12485),
            .I(N__12479));
    Odrv12 I__2693 (
            .O(N__12482),
            .I(P1A4_c_i));
    Odrv4 I__2692 (
            .O(N__12479),
            .I(P1A4_c_i));
    InMux I__2691 (
            .O(N__12474),
            .I(N__12471));
    LocalMux I__2690 (
            .O(N__12471),
            .I(N__12468));
    Span4Mux_v I__2689 (
            .O(N__12468),
            .I(N__12465));
    Odrv4 I__2688 (
            .O(N__12465),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_0 ));
    InMux I__2687 (
            .O(N__12462),
            .I(N__12459));
    LocalMux I__2686 (
            .O(N__12459),
            .I(N__12456));
    Span4Mux_v I__2685 (
            .O(N__12456),
            .I(N__12453));
    Odrv4 I__2684 (
            .O(N__12453),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_1 ));
    InMux I__2683 (
            .O(N__12450),
            .I(N__12446));
    InMux I__2682 (
            .O(N__12449),
            .I(N__12443));
    LocalMux I__2681 (
            .O(N__12446),
            .I(N__12440));
    LocalMux I__2680 (
            .O(N__12443),
            .I(\DUT.fifo_rx_inst.rFifoDataro_0 ));
    Odrv4 I__2679 (
            .O(N__12440),
            .I(\DUT.fifo_rx_inst.rFifoDataro_0 ));
    CascadeMux I__2678 (
            .O(N__12435),
            .I(N__12431));
    InMux I__2677 (
            .O(N__12434),
            .I(N__12428));
    InMux I__2676 (
            .O(N__12431),
            .I(N__12425));
    LocalMux I__2675 (
            .O(N__12428),
            .I(N__12422));
    LocalMux I__2674 (
            .O(N__12425),
            .I(\DUT.fifo_rx_inst.rFifoDataro_1 ));
    Odrv4 I__2673 (
            .O(N__12422),
            .I(\DUT.fifo_rx_inst.rFifoDataro_1 ));
    InMux I__2672 (
            .O(N__12417),
            .I(N__12413));
    InMux I__2671 (
            .O(N__12416),
            .I(N__12410));
    LocalMux I__2670 (
            .O(N__12413),
            .I(N__12407));
    LocalMux I__2669 (
            .O(N__12410),
            .I(\DUT.fifo_rx_inst.rFifoDataro_2 ));
    Odrv4 I__2668 (
            .O(N__12407),
            .I(\DUT.fifo_rx_inst.rFifoDataro_2 ));
    CascadeMux I__2667 (
            .O(N__12402),
            .I(N__12397));
    CascadeMux I__2666 (
            .O(N__12401),
            .I(N__12393));
    CascadeMux I__2665 (
            .O(N__12400),
            .I(N__12390));
    InMux I__2664 (
            .O(N__12397),
            .I(N__12375));
    InMux I__2663 (
            .O(N__12396),
            .I(N__12375));
    InMux I__2662 (
            .O(N__12393),
            .I(N__12375));
    InMux I__2661 (
            .O(N__12390),
            .I(N__12375));
    InMux I__2660 (
            .O(N__12389),
            .I(N__12375));
    InMux I__2659 (
            .O(N__12388),
            .I(N__12375));
    LocalMux I__2658 (
            .O(N__12375),
            .I(N__12371));
    CascadeMux I__2657 (
            .O(N__12374),
            .I(N__12366));
    Span4Mux_v I__2656 (
            .O(N__12371),
            .I(N__12363));
    InMux I__2655 (
            .O(N__12370),
            .I(N__12356));
    InMux I__2654 (
            .O(N__12369),
            .I(N__12356));
    InMux I__2653 (
            .O(N__12366),
            .I(N__12356));
    Odrv4 I__2652 (
            .O(N__12363),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_0 ));
    LocalMux I__2651 (
            .O(N__12356),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_0 ));
    InMux I__2650 (
            .O(N__12351),
            .I(N__12333));
    InMux I__2649 (
            .O(N__12350),
            .I(N__12333));
    InMux I__2648 (
            .O(N__12349),
            .I(N__12333));
    InMux I__2647 (
            .O(N__12348),
            .I(N__12333));
    InMux I__2646 (
            .O(N__12347),
            .I(N__12333));
    InMux I__2645 (
            .O(N__12346),
            .I(N__12333));
    LocalMux I__2644 (
            .O(N__12333),
            .I(N__12330));
    Span4Mux_v I__2643 (
            .O(N__12330),
            .I(N__12325));
    InMux I__2642 (
            .O(N__12329),
            .I(N__12320));
    InMux I__2641 (
            .O(N__12328),
            .I(N__12320));
    Odrv4 I__2640 (
            .O(N__12325),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_1 ));
    LocalMux I__2639 (
            .O(N__12320),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_1 ));
    InMux I__2638 (
            .O(N__12315),
            .I(N__12308));
    InMux I__2637 (
            .O(N__12314),
            .I(N__12305));
    InMux I__2636 (
            .O(N__12313),
            .I(N__12302));
    InMux I__2635 (
            .O(N__12312),
            .I(N__12296));
    InMux I__2634 (
            .O(N__12311),
            .I(N__12296));
    LocalMux I__2633 (
            .O(N__12308),
            .I(N__12289));
    LocalMux I__2632 (
            .O(N__12305),
            .I(N__12289));
    LocalMux I__2631 (
            .O(N__12302),
            .I(N__12289));
    InMux I__2630 (
            .O(N__12301),
            .I(N__12286));
    LocalMux I__2629 (
            .O(N__12296),
            .I(N__12283));
    Odrv4 I__2628 (
            .O(N__12289),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_0 ));
    LocalMux I__2627 (
            .O(N__12286),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_0 ));
    Odrv4 I__2626 (
            .O(N__12283),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_0 ));
    InMux I__2625 (
            .O(N__12276),
            .I(N__12273));
    LocalMux I__2624 (
            .O(N__12273),
            .I(N__12268));
    InMux I__2623 (
            .O(N__12272),
            .I(N__12265));
    InMux I__2622 (
            .O(N__12271),
            .I(N__12260));
    Span4Mux_h I__2621 (
            .O(N__12268),
            .I(N__12255));
    LocalMux I__2620 (
            .O(N__12265),
            .I(N__12255));
    InMux I__2619 (
            .O(N__12264),
            .I(N__12250));
    InMux I__2618 (
            .O(N__12263),
            .I(N__12250));
    LocalMux I__2617 (
            .O(N__12260),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_1 ));
    Odrv4 I__2616 (
            .O(N__12255),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_1 ));
    LocalMux I__2615 (
            .O(N__12250),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_1 ));
    InMux I__2614 (
            .O(N__12243),
            .I(N__12235));
    InMux I__2613 (
            .O(N__12242),
            .I(N__12232));
    InMux I__2612 (
            .O(N__12241),
            .I(N__12229));
    InMux I__2611 (
            .O(N__12240),
            .I(N__12226));
    InMux I__2610 (
            .O(N__12239),
            .I(N__12221));
    InMux I__2609 (
            .O(N__12238),
            .I(N__12221));
    LocalMux I__2608 (
            .O(N__12235),
            .I(N__12214));
    LocalMux I__2607 (
            .O(N__12232),
            .I(N__12214));
    LocalMux I__2606 (
            .O(N__12229),
            .I(N__12214));
    LocalMux I__2605 (
            .O(N__12226),
            .I(\DUT.fifo_tx_inst.N_104 ));
    LocalMux I__2604 (
            .O(N__12221),
            .I(\DUT.fifo_tx_inst.N_104 ));
    Odrv12 I__2603 (
            .O(N__12214),
            .I(\DUT.fifo_tx_inst.N_104 ));
    CEMux I__2602 (
            .O(N__12207),
            .I(N__12204));
    LocalMux I__2601 (
            .O(N__12204),
            .I(N__12200));
    InMux I__2600 (
            .O(N__12203),
            .I(N__12197));
    Span4Mux_v I__2599 (
            .O(N__12200),
            .I(N__12194));
    LocalMux I__2598 (
            .O(N__12197),
            .I(N__12191));
    Odrv4 I__2597 (
            .O(N__12194),
            .I(\DUT.fifo_tx_inst.rFifoData_awe2 ));
    Odrv12 I__2596 (
            .O(N__12191),
            .I(\DUT.fifo_tx_inst.rFifoData_awe2 ));
    CascadeMux I__2595 (
            .O(N__12186),
            .I(\DUT.fifo_rx_inst.rWritePtr16_cascade_ ));
    CascadeMux I__2594 (
            .O(N__12183),
            .I(N__12180));
    InMux I__2593 (
            .O(N__12180),
            .I(N__12174));
    InMux I__2592 (
            .O(N__12179),
            .I(N__12174));
    LocalMux I__2591 (
            .O(N__12174),
            .I(N__12171));
    Span4Mux_h I__2590 (
            .O(N__12171),
            .I(N__12161));
    InMux I__2589 (
            .O(N__12170),
            .I(N__12158));
    InMux I__2588 (
            .O(N__12169),
            .I(N__12145));
    InMux I__2587 (
            .O(N__12168),
            .I(N__12145));
    InMux I__2586 (
            .O(N__12167),
            .I(N__12145));
    InMux I__2585 (
            .O(N__12166),
            .I(N__12145));
    InMux I__2584 (
            .O(N__12165),
            .I(N__12145));
    InMux I__2583 (
            .O(N__12164),
            .I(N__12145));
    Odrv4 I__2582 (
            .O(N__12161),
            .I(\DUT.fifo_rx_inst.rWritePtr16 ));
    LocalMux I__2581 (
            .O(N__12158),
            .I(\DUT.fifo_rx_inst.rWritePtr16 ));
    LocalMux I__2580 (
            .O(N__12145),
            .I(\DUT.fifo_rx_inst.rWritePtr16 ));
    CascadeMux I__2579 (
            .O(N__12138),
            .I(\DUT.fifo_rx_inst.rFifoDataror_1_0_cascade_ ));
    InMux I__2578 (
            .O(N__12135),
            .I(N__12132));
    LocalMux I__2577 (
            .O(N__12132),
            .I(N__12129));
    Odrv4 I__2576 (
            .O(N__12129),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_3 ));
    CascadeMux I__2575 (
            .O(N__12126),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ));
    InMux I__2574 (
            .O(N__12123),
            .I(N__12120));
    LocalMux I__2573 (
            .O(N__12120),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_3 ));
    InMux I__2572 (
            .O(N__12117),
            .I(N__12114));
    LocalMux I__2571 (
            .O(N__12114),
            .I(N__12111));
    Odrv4 I__2570 (
            .O(N__12111),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_4 ));
    CascadeMux I__2569 (
            .O(N__12108),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4_cascade_ ));
    CascadeMux I__2568 (
            .O(N__12105),
            .I(N__12102));
    InMux I__2567 (
            .O(N__12102),
            .I(N__12099));
    LocalMux I__2566 (
            .O(N__12099),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_4 ));
    InMux I__2565 (
            .O(N__12096),
            .I(N__12093));
    LocalMux I__2564 (
            .O(N__12093),
            .I(N__12090));
    Odrv12 I__2563 (
            .O(N__12090),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_5 ));
    CascadeMux I__2562 (
            .O(N__12087),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ));
    CEMux I__2561 (
            .O(N__12084),
            .I(N__12080));
    InMux I__2560 (
            .O(N__12083),
            .I(N__12077));
    LocalMux I__2559 (
            .O(N__12080),
            .I(N__12074));
    LocalMux I__2558 (
            .O(N__12077),
            .I(N__12071));
    Span4Mux_v I__2557 (
            .O(N__12074),
            .I(N__12068));
    Span4Mux_h I__2556 (
            .O(N__12071),
            .I(N__12065));
    Span4Mux_h I__2555 (
            .O(N__12068),
            .I(N__12060));
    Span4Mux_v I__2554 (
            .O(N__12065),
            .I(N__12060));
    Odrv4 I__2553 (
            .O(N__12060),
            .I(\DUT.fifo_rx_inst.N_57 ));
    InMux I__2552 (
            .O(N__12057),
            .I(N__12054));
    LocalMux I__2551 (
            .O(N__12054),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_6 ));
    CascadeMux I__2550 (
            .O(N__12051),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6_cascade_ ));
    InMux I__2549 (
            .O(N__12048),
            .I(N__12045));
    LocalMux I__2548 (
            .O(N__12045),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_6 ));
    InMux I__2547 (
            .O(N__12042),
            .I(N__12039));
    LocalMux I__2546 (
            .O(N__12039),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_7 ));
    CascadeMux I__2545 (
            .O(N__12036),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7_cascade_ ));
    InMux I__2544 (
            .O(N__12033),
            .I(N__12030));
    LocalMux I__2543 (
            .O(N__12030),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_7 ));
    InMux I__2542 (
            .O(N__12027),
            .I(N__12023));
    InMux I__2541 (
            .O(N__12026),
            .I(N__12020));
    LocalMux I__2540 (
            .O(N__12023),
            .I(N__12017));
    LocalMux I__2539 (
            .O(N__12020),
            .I(\DUT.fifo_rx_inst.rFifoDataro_3 ));
    Odrv4 I__2538 (
            .O(N__12017),
            .I(\DUT.fifo_rx_inst.rFifoDataro_3 ));
    InMux I__2537 (
            .O(N__12012),
            .I(N__12008));
    InMux I__2536 (
            .O(N__12011),
            .I(N__12005));
    LocalMux I__2535 (
            .O(N__12008),
            .I(N__12002));
    LocalMux I__2534 (
            .O(N__12005),
            .I(\DUT.fifo_tx_inst.rFifoDataro_0 ));
    Odrv4 I__2533 (
            .O(N__12002),
            .I(\DUT.fifo_tx_inst.rFifoDataro_0 ));
    CEMux I__2532 (
            .O(N__11997),
            .I(N__11994));
    LocalMux I__2531 (
            .O(N__11994),
            .I(N__11990));
    InMux I__2530 (
            .O(N__11993),
            .I(N__11987));
    Span4Mux_v I__2529 (
            .O(N__11990),
            .I(N__11984));
    LocalMux I__2528 (
            .O(N__11987),
            .I(N__11981));
    Span4Mux_v I__2527 (
            .O(N__11984),
            .I(N__11978));
    Span4Mux_h I__2526 (
            .O(N__11981),
            .I(N__11975));
    Span4Mux_h I__2525 (
            .O(N__11978),
            .I(N__11972));
    Span4Mux_v I__2524 (
            .O(N__11975),
            .I(N__11969));
    Odrv4 I__2523 (
            .O(N__11972),
            .I(\DUT.fifo_tx_inst.rFifoData_awe1 ));
    Odrv4 I__2522 (
            .O(N__11969),
            .I(\DUT.fifo_tx_inst.rFifoData_awe1 ));
    CascadeMux I__2521 (
            .O(N__11964),
            .I(N__11960));
    InMux I__2520 (
            .O(N__11963),
            .I(N__11957));
    InMux I__2519 (
            .O(N__11960),
            .I(N__11954));
    LocalMux I__2518 (
            .O(N__11957),
            .I(\DUT.fifo_tx_inst.rFifoDataro_1 ));
    LocalMux I__2517 (
            .O(N__11954),
            .I(\DUT.fifo_tx_inst.rFifoDataro_1 ));
    InMux I__2516 (
            .O(N__11949),
            .I(N__11945));
    InMux I__2515 (
            .O(N__11948),
            .I(N__11942));
    LocalMux I__2514 (
            .O(N__11945),
            .I(\DUT.fifo_tx_inst.rFifoDataro_2 ));
    LocalMux I__2513 (
            .O(N__11942),
            .I(\DUT.fifo_tx_inst.rFifoDataro_2 ));
    InMux I__2512 (
            .O(N__11937),
            .I(N__11933));
    InMux I__2511 (
            .O(N__11936),
            .I(N__11930));
    LocalMux I__2510 (
            .O(N__11933),
            .I(\DUT.fifo_tx_inst.rFifoDataro_3 ));
    LocalMux I__2509 (
            .O(N__11930),
            .I(\DUT.fifo_tx_inst.rFifoDataro_3 ));
    InMux I__2508 (
            .O(N__11925),
            .I(N__11922));
    LocalMux I__2507 (
            .O(N__11922),
            .I(N__11919));
    Span4Mux_h I__2506 (
            .O(N__11919),
            .I(N__11916));
    Odrv4 I__2505 (
            .O(N__11916),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_0 ));
    InMux I__2504 (
            .O(N__11913),
            .I(N__11910));
    LocalMux I__2503 (
            .O(N__11910),
            .I(N__11907));
    Span4Mux_h I__2502 (
            .O(N__11907),
            .I(N__11904));
    Odrv4 I__2501 (
            .O(N__11904),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_1 ));
    InMux I__2500 (
            .O(N__11901),
            .I(N__11898));
    LocalMux I__2499 (
            .O(N__11898),
            .I(N__11895));
    Odrv4 I__2498 (
            .O(N__11895),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_2 ));
    InMux I__2497 (
            .O(N__11892),
            .I(N__11889));
    LocalMux I__2496 (
            .O(N__11889),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_3 ));
    InMux I__2495 (
            .O(N__11886),
            .I(N__11883));
    LocalMux I__2494 (
            .O(N__11883),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_4 ));
    InMux I__2493 (
            .O(N__11880),
            .I(N__11877));
    LocalMux I__2492 (
            .O(N__11877),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_5 ));
    InMux I__2491 (
            .O(N__11874),
            .I(N__11871));
    LocalMux I__2490 (
            .O(N__11871),
            .I(N__11868));
    Odrv4 I__2489 (
            .O(N__11868),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_6 ));
    InMux I__2488 (
            .O(N__11865),
            .I(N__11862));
    LocalMux I__2487 (
            .O(N__11862),
            .I(N__11859));
    Span4Mux_h I__2486 (
            .O(N__11859),
            .I(N__11856));
    Odrv4 I__2485 (
            .O(N__11856),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_7 ));
    CEMux I__2484 (
            .O(N__11853),
            .I(N__11849));
    CEMux I__2483 (
            .O(N__11852),
            .I(N__11845));
    LocalMux I__2482 (
            .O(N__11849),
            .I(N__11842));
    CEMux I__2481 (
            .O(N__11848),
            .I(N__11839));
    LocalMux I__2480 (
            .O(N__11845),
            .I(N__11835));
    Span4Mux_s2_v I__2479 (
            .O(N__11842),
            .I(N__11829));
    LocalMux I__2478 (
            .O(N__11839),
            .I(N__11829));
    InMux I__2477 (
            .O(N__11838),
            .I(N__11826));
    Span4Mux_v I__2476 (
            .O(N__11835),
            .I(N__11823));
    CEMux I__2475 (
            .O(N__11834),
            .I(N__11820));
    Span4Mux_v I__2474 (
            .O(N__11829),
            .I(N__11815));
    LocalMux I__2473 (
            .O(N__11826),
            .I(N__11815));
    Span4Mux_h I__2472 (
            .O(N__11823),
            .I(N__11812));
    LocalMux I__2471 (
            .O(N__11820),
            .I(N__11809));
    Span4Mux_h I__2470 (
            .O(N__11815),
            .I(N__11806));
    Odrv4 I__2469 (
            .O(N__11812),
            .I(\DUT.fifo_tx_inst.rFifoData_awe0 ));
    Odrv12 I__2468 (
            .O(N__11809),
            .I(\DUT.fifo_tx_inst.rFifoData_awe0 ));
    Odrv4 I__2467 (
            .O(N__11806),
            .I(\DUT.fifo_tx_inst.rFifoData_awe0 ));
    InMux I__2466 (
            .O(N__11799),
            .I(N__11796));
    LocalMux I__2465 (
            .O(N__11796),
            .I(N__11793));
    Odrv4 I__2464 (
            .O(N__11793),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_5 ));
    CascadeMux I__2463 (
            .O(N__11790),
            .I(N__11787));
    InMux I__2462 (
            .O(N__11787),
            .I(N__11784));
    LocalMux I__2461 (
            .O(N__11784),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_6 ));
    InMux I__2460 (
            .O(N__11781),
            .I(N__11778));
    LocalMux I__2459 (
            .O(N__11778),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_7 ));
    CascadeMux I__2458 (
            .O(N__11775),
            .I(N__11772));
    InMux I__2457 (
            .O(N__11772),
            .I(N__11769));
    LocalMux I__2456 (
            .O(N__11769),
            .I(N__11766));
    Odrv4 I__2455 (
            .O(N__11766),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_2 ));
    CascadeMux I__2454 (
            .O(N__11763),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_ ));
    InMux I__2453 (
            .O(N__11760),
            .I(N__11757));
    LocalMux I__2452 (
            .O(N__11757),
            .I(N__11754));
    Odrv4 I__2451 (
            .O(N__11754),
            .I(\DUT.rFifoDatarx_2 ));
    InMux I__2450 (
            .O(N__11751),
            .I(N__11748));
    LocalMux I__2449 (
            .O(N__11748),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_2 ));
    InMux I__2448 (
            .O(N__11745),
            .I(N__11732));
    InMux I__2447 (
            .O(N__11744),
            .I(N__11732));
    InMux I__2446 (
            .O(N__11743),
            .I(N__11732));
    InMux I__2445 (
            .O(N__11742),
            .I(N__11723));
    InMux I__2444 (
            .O(N__11741),
            .I(N__11716));
    InMux I__2443 (
            .O(N__11740),
            .I(N__11716));
    InMux I__2442 (
            .O(N__11739),
            .I(N__11716));
    LocalMux I__2441 (
            .O(N__11732),
            .I(N__11713));
    InMux I__2440 (
            .O(N__11731),
            .I(N__11708));
    InMux I__2439 (
            .O(N__11730),
            .I(N__11708));
    InMux I__2438 (
            .O(N__11729),
            .I(N__11699));
    InMux I__2437 (
            .O(N__11728),
            .I(N__11699));
    InMux I__2436 (
            .O(N__11727),
            .I(N__11699));
    InMux I__2435 (
            .O(N__11726),
            .I(N__11699));
    LocalMux I__2434 (
            .O(N__11723),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__2433 (
            .O(N__11716),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    Odrv4 I__2432 (
            .O(N__11713),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__2431 (
            .O(N__11708),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__2430 (
            .O(N__11699),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    InMux I__2429 (
            .O(N__11688),
            .I(N__11685));
    LocalMux I__2428 (
            .O(N__11685),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_3 ));
    CascadeMux I__2427 (
            .O(N__11682),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ));
    CascadeMux I__2426 (
            .O(N__11679),
            .I(N__11670));
    CascadeMux I__2425 (
            .O(N__11678),
            .I(N__11667));
    CascadeMux I__2424 (
            .O(N__11677),
            .I(N__11659));
    CascadeMux I__2423 (
            .O(N__11676),
            .I(N__11651));
    InMux I__2422 (
            .O(N__11675),
            .I(N__11638));
    InMux I__2421 (
            .O(N__11674),
            .I(N__11638));
    InMux I__2420 (
            .O(N__11673),
            .I(N__11638));
    InMux I__2419 (
            .O(N__11670),
            .I(N__11638));
    InMux I__2418 (
            .O(N__11667),
            .I(N__11638));
    InMux I__2417 (
            .O(N__11666),
            .I(N__11638));
    CascadeMux I__2416 (
            .O(N__11665),
            .I(N__11632));
    InMux I__2415 (
            .O(N__11664),
            .I(N__11619));
    InMux I__2414 (
            .O(N__11663),
            .I(N__11619));
    InMux I__2413 (
            .O(N__11662),
            .I(N__11619));
    InMux I__2412 (
            .O(N__11659),
            .I(N__11619));
    InMux I__2411 (
            .O(N__11658),
            .I(N__11619));
    InMux I__2410 (
            .O(N__11657),
            .I(N__11619));
    InMux I__2409 (
            .O(N__11656),
            .I(N__11610));
    InMux I__2408 (
            .O(N__11655),
            .I(N__11610));
    InMux I__2407 (
            .O(N__11654),
            .I(N__11610));
    InMux I__2406 (
            .O(N__11651),
            .I(N__11610));
    LocalMux I__2405 (
            .O(N__11638),
            .I(N__11607));
    InMux I__2404 (
            .O(N__11637),
            .I(N__11598));
    InMux I__2403 (
            .O(N__11636),
            .I(N__11598));
    InMux I__2402 (
            .O(N__11635),
            .I(N__11598));
    InMux I__2401 (
            .O(N__11632),
            .I(N__11598));
    LocalMux I__2400 (
            .O(N__11619),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__2399 (
            .O(N__11610),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    Odrv4 I__2398 (
            .O(N__11607),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__2397 (
            .O(N__11598),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    InMux I__2396 (
            .O(N__11589),
            .I(N__11586));
    LocalMux I__2395 (
            .O(N__11586),
            .I(N__11583));
    Odrv12 I__2394 (
            .O(N__11583),
            .I(\DUT.rFifoDatarx_3 ));
    InMux I__2393 (
            .O(N__11580),
            .I(N__11577));
    LocalMux I__2392 (
            .O(N__11577),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_3 ));
    CascadeMux I__2391 (
            .O(N__11574),
            .I(N__11569));
    CascadeMux I__2390 (
            .O(N__11573),
            .I(N__11565));
    CascadeMux I__2389 (
            .O(N__11572),
            .I(N__11559));
    InMux I__2388 (
            .O(N__11569),
            .I(N__11552));
    InMux I__2387 (
            .O(N__11568),
            .I(N__11552));
    InMux I__2386 (
            .O(N__11565),
            .I(N__11552));
    InMux I__2385 (
            .O(N__11564),
            .I(N__11549));
    InMux I__2384 (
            .O(N__11563),
            .I(N__11539));
    InMux I__2383 (
            .O(N__11562),
            .I(N__11539));
    InMux I__2382 (
            .O(N__11559),
            .I(N__11536));
    LocalMux I__2381 (
            .O(N__11552),
            .I(N__11533));
    LocalMux I__2380 (
            .O(N__11549),
            .I(N__11530));
    InMux I__2379 (
            .O(N__11548),
            .I(N__11523));
    InMux I__2378 (
            .O(N__11547),
            .I(N__11523));
    InMux I__2377 (
            .O(N__11546),
            .I(N__11523));
    InMux I__2376 (
            .O(N__11545),
            .I(N__11520));
    InMux I__2375 (
            .O(N__11544),
            .I(N__11517));
    LocalMux I__2374 (
            .O(N__11539),
            .I(N__11510));
    LocalMux I__2373 (
            .O(N__11536),
            .I(N__11510));
    Span4Mux_h I__2372 (
            .O(N__11533),
            .I(N__11510));
    Odrv12 I__2371 (
            .O(N__11530),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_5 ));
    LocalMux I__2370 (
            .O(N__11523),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_5 ));
    LocalMux I__2369 (
            .O(N__11520),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_5 ));
    LocalMux I__2368 (
            .O(N__11517),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_5 ));
    Odrv4 I__2367 (
            .O(N__11510),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_5 ));
    CascadeMux I__2366 (
            .O(N__11499),
            .I(N__11494));
    InMux I__2365 (
            .O(N__11498),
            .I(N__11484));
    CascadeMux I__2364 (
            .O(N__11497),
            .I(N__11481));
    InMux I__2363 (
            .O(N__11494),
            .I(N__11475));
    InMux I__2362 (
            .O(N__11493),
            .I(N__11475));
    InMux I__2361 (
            .O(N__11492),
            .I(N__11468));
    InMux I__2360 (
            .O(N__11491),
            .I(N__11468));
    InMux I__2359 (
            .O(N__11490),
            .I(N__11468));
    InMux I__2358 (
            .O(N__11489),
            .I(N__11462));
    InMux I__2357 (
            .O(N__11488),
            .I(N__11462));
    CascadeMux I__2356 (
            .O(N__11487),
            .I(N__11459));
    LocalMux I__2355 (
            .O(N__11484),
            .I(N__11456));
    InMux I__2354 (
            .O(N__11481),
            .I(N__11452));
    InMux I__2353 (
            .O(N__11480),
            .I(N__11449));
    LocalMux I__2352 (
            .O(N__11475),
            .I(N__11444));
    LocalMux I__2351 (
            .O(N__11468),
            .I(N__11444));
    CascadeMux I__2350 (
            .O(N__11467),
            .I(N__11441));
    LocalMux I__2349 (
            .O(N__11462),
            .I(N__11438));
    InMux I__2348 (
            .O(N__11459),
            .I(N__11435));
    Span4Mux_v I__2347 (
            .O(N__11456),
            .I(N__11432));
    InMux I__2346 (
            .O(N__11455),
            .I(N__11429));
    LocalMux I__2345 (
            .O(N__11452),
            .I(N__11426));
    LocalMux I__2344 (
            .O(N__11449),
            .I(N__11421));
    Span4Mux_v I__2343 (
            .O(N__11444),
            .I(N__11421));
    InMux I__2342 (
            .O(N__11441),
            .I(N__11418));
    Span4Mux_v I__2341 (
            .O(N__11438),
            .I(N__11415));
    LocalMux I__2340 (
            .O(N__11435),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_4 ));
    Odrv4 I__2339 (
            .O(N__11432),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_4 ));
    LocalMux I__2338 (
            .O(N__11429),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_4 ));
    Odrv4 I__2337 (
            .O(N__11426),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_4 ));
    Odrv4 I__2336 (
            .O(N__11421),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_4 ));
    LocalMux I__2335 (
            .O(N__11418),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_4 ));
    Odrv4 I__2334 (
            .O(N__11415),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_4 ));
    InMux I__2333 (
            .O(N__11400),
            .I(N__11394));
    InMux I__2332 (
            .O(N__11399),
            .I(N__11389));
    InMux I__2331 (
            .O(N__11398),
            .I(N__11384));
    InMux I__2330 (
            .O(N__11397),
            .I(N__11384));
    LocalMux I__2329 (
            .O(N__11394),
            .I(N__11381));
    CascadeMux I__2328 (
            .O(N__11393),
            .I(N__11374));
    InMux I__2327 (
            .O(N__11392),
            .I(N__11371));
    LocalMux I__2326 (
            .O(N__11389),
            .I(N__11368));
    LocalMux I__2325 (
            .O(N__11384),
            .I(N__11363));
    Span4Mux_h I__2324 (
            .O(N__11381),
            .I(N__11363));
    InMux I__2323 (
            .O(N__11380),
            .I(N__11356));
    InMux I__2322 (
            .O(N__11379),
            .I(N__11356));
    InMux I__2321 (
            .O(N__11378),
            .I(N__11356));
    InMux I__2320 (
            .O(N__11377),
            .I(N__11353));
    InMux I__2319 (
            .O(N__11374),
            .I(N__11350));
    LocalMux I__2318 (
            .O(N__11371),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_1 ));
    Odrv4 I__2317 (
            .O(N__11368),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_1 ));
    Odrv4 I__2316 (
            .O(N__11363),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_1 ));
    LocalMux I__2315 (
            .O(N__11356),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_1 ));
    LocalMux I__2314 (
            .O(N__11353),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_1 ));
    LocalMux I__2313 (
            .O(N__11350),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_1 ));
    InMux I__2312 (
            .O(N__11337),
            .I(N__11333));
    CascadeMux I__2311 (
            .O(N__11336),
            .I(N__11329));
    LocalMux I__2310 (
            .O(N__11333),
            .I(N__11326));
    InMux I__2309 (
            .O(N__11332),
            .I(N__11323));
    InMux I__2308 (
            .O(N__11329),
            .I(N__11318));
    Span4Mux_v I__2307 (
            .O(N__11326),
            .I(N__11313));
    LocalMux I__2306 (
            .O(N__11323),
            .I(N__11313));
    InMux I__2305 (
            .O(N__11322),
            .I(N__11308));
    InMux I__2304 (
            .O(N__11321),
            .I(N__11308));
    LocalMux I__2303 (
            .O(N__11318),
            .I(\DUT.uart_inst0.recv_stateZ0Z_3 ));
    Odrv4 I__2302 (
            .O(N__11313),
            .I(\DUT.uart_inst0.recv_stateZ0Z_3 ));
    LocalMux I__2301 (
            .O(N__11308),
            .I(\DUT.uart_inst0.recv_stateZ0Z_3 ));
    InMux I__2300 (
            .O(N__11301),
            .I(N__11298));
    LocalMux I__2299 (
            .O(N__11298),
            .I(N__11295));
    Span4Mux_v I__2298 (
            .O(N__11295),
            .I(N__11292));
    Odrv4 I__2297 (
            .O(N__11292),
            .I(\DUT.uart_inst0.m6_e_2 ));
    CascadeMux I__2296 (
            .O(N__11289),
            .I(\DUT.uart_inst0.m6_e_3_cascade_ ));
    InMux I__2295 (
            .O(N__11286),
            .I(N__11282));
    InMux I__2294 (
            .O(N__11285),
            .I(N__11279));
    LocalMux I__2293 (
            .O(N__11282),
            .I(N__11276));
    LocalMux I__2292 (
            .O(N__11279),
            .I(\DUT.uart_inst0.N_15_mux ));
    Odrv4 I__2291 (
            .O(N__11276),
            .I(\DUT.uart_inst0.N_15_mux ));
    InMux I__2290 (
            .O(N__11271),
            .I(N__11268));
    LocalMux I__2289 (
            .O(N__11268),
            .I(\DUT.uart_inst0.N_18_mux_1 ));
    CascadeMux I__2288 (
            .O(N__11265),
            .I(N__11258));
    InMux I__2287 (
            .O(N__11264),
            .I(N__11251));
    InMux I__2286 (
            .O(N__11263),
            .I(N__11251));
    InMux I__2285 (
            .O(N__11262),
            .I(N__11246));
    InMux I__2284 (
            .O(N__11261),
            .I(N__11246));
    InMux I__2283 (
            .O(N__11258),
            .I(N__11241));
    InMux I__2282 (
            .O(N__11257),
            .I(N__11238));
    InMux I__2281 (
            .O(N__11256),
            .I(N__11235));
    LocalMux I__2280 (
            .O(N__11251),
            .I(N__11230));
    LocalMux I__2279 (
            .O(N__11246),
            .I(N__11230));
    InMux I__2278 (
            .O(N__11245),
            .I(N__11225));
    InMux I__2277 (
            .O(N__11244),
            .I(N__11225));
    LocalMux I__2276 (
            .O(N__11241),
            .I(N__11221));
    LocalMux I__2275 (
            .O(N__11238),
            .I(N__11213));
    LocalMux I__2274 (
            .O(N__11235),
            .I(N__11213));
    Span4Mux_h I__2273 (
            .O(N__11230),
            .I(N__11208));
    LocalMux I__2272 (
            .O(N__11225),
            .I(N__11208));
    CascadeMux I__2271 (
            .O(N__11224),
            .I(N__11205));
    Span4Mux_v I__2270 (
            .O(N__11221),
            .I(N__11202));
    InMux I__2269 (
            .O(N__11220),
            .I(N__11197));
    InMux I__2268 (
            .O(N__11219),
            .I(N__11197));
    InMux I__2267 (
            .O(N__11218),
            .I(N__11194));
    Span4Mux_v I__2266 (
            .O(N__11213),
            .I(N__11189));
    Span4Mux_v I__2265 (
            .O(N__11208),
            .I(N__11189));
    InMux I__2264 (
            .O(N__11205),
            .I(N__11186));
    Odrv4 I__2263 (
            .O(N__11202),
            .I(\DUT.uart_inst0.rx_countdownZ1Z_3 ));
    LocalMux I__2262 (
            .O(N__11197),
            .I(\DUT.uart_inst0.rx_countdownZ1Z_3 ));
    LocalMux I__2261 (
            .O(N__11194),
            .I(\DUT.uart_inst0.rx_countdownZ1Z_3 ));
    Odrv4 I__2260 (
            .O(N__11189),
            .I(\DUT.uart_inst0.rx_countdownZ1Z_3 ));
    LocalMux I__2259 (
            .O(N__11186),
            .I(\DUT.uart_inst0.rx_countdownZ1Z_3 ));
    InMux I__2258 (
            .O(N__11175),
            .I(N__11170));
    InMux I__2257 (
            .O(N__11174),
            .I(N__11167));
    InMux I__2256 (
            .O(N__11173),
            .I(N__11164));
    LocalMux I__2255 (
            .O(N__11170),
            .I(\DUT.uart_inst0.recv_stateZ0Z_4 ));
    LocalMux I__2254 (
            .O(N__11167),
            .I(\DUT.uart_inst0.recv_stateZ0Z_4 ));
    LocalMux I__2253 (
            .O(N__11164),
            .I(\DUT.uart_inst0.recv_stateZ0Z_4 ));
    InMux I__2252 (
            .O(N__11157),
            .I(N__11150));
    CascadeMux I__2251 (
            .O(N__11156),
            .I(N__11146));
    InMux I__2250 (
            .O(N__11155),
            .I(N__11141));
    InMux I__2249 (
            .O(N__11154),
            .I(N__11141));
    InMux I__2248 (
            .O(N__11153),
            .I(N__11136));
    LocalMux I__2247 (
            .O(N__11150),
            .I(N__11133));
    InMux I__2246 (
            .O(N__11149),
            .I(N__11128));
    InMux I__2245 (
            .O(N__11146),
            .I(N__11128));
    LocalMux I__2244 (
            .O(N__11141),
            .I(N__11125));
    InMux I__2243 (
            .O(N__11140),
            .I(N__11120));
    InMux I__2242 (
            .O(N__11139),
            .I(N__11120));
    LocalMux I__2241 (
            .O(N__11136),
            .I(N__11109));
    Span4Mux_v I__2240 (
            .O(N__11133),
            .I(N__11109));
    LocalMux I__2239 (
            .O(N__11128),
            .I(N__11109));
    Span4Mux_h I__2238 (
            .O(N__11125),
            .I(N__11104));
    LocalMux I__2237 (
            .O(N__11120),
            .I(N__11104));
    InMux I__2236 (
            .O(N__11119),
            .I(N__11095));
    InMux I__2235 (
            .O(N__11118),
            .I(N__11095));
    InMux I__2234 (
            .O(N__11117),
            .I(N__11095));
    InMux I__2233 (
            .O(N__11116),
            .I(N__11095));
    Span4Mux_h I__2232 (
            .O(N__11109),
            .I(N__11092));
    Odrv4 I__2231 (
            .O(N__11104),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_2 ));
    LocalMux I__2230 (
            .O(N__11095),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_2 ));
    Odrv4 I__2229 (
            .O(N__11092),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_2 ));
    CascadeMux I__2228 (
            .O(N__11085),
            .I(N__11082));
    InMux I__2227 (
            .O(N__11082),
            .I(N__11079));
    LocalMux I__2226 (
            .O(N__11079),
            .I(N__11076));
    Odrv4 I__2225 (
            .O(N__11076),
            .I(\DUT.uart_inst0.G_19_0_a5_2 ));
    CascadeMux I__2224 (
            .O(N__11073),
            .I(N__11070));
    InMux I__2223 (
            .O(N__11070),
            .I(N__11067));
    LocalMux I__2222 (
            .O(N__11067),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_0 ));
    InMux I__2221 (
            .O(N__11064),
            .I(N__11061));
    LocalMux I__2220 (
            .O(N__11061),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_1 ));
    CascadeMux I__2219 (
            .O(N__11058),
            .I(N__11055));
    InMux I__2218 (
            .O(N__11055),
            .I(N__11052));
    LocalMux I__2217 (
            .O(N__11052),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_4 ));
    InMux I__2216 (
            .O(N__11049),
            .I(N__11043));
    InMux I__2215 (
            .O(N__11048),
            .I(N__11043));
    LocalMux I__2214 (
            .O(N__11043),
            .I(\DUT.fifo_rx_inst.N_77_mux ));
    InMux I__2213 (
            .O(N__11040),
            .I(N__11036));
    InMux I__2212 (
            .O(N__11039),
            .I(N__11032));
    LocalMux I__2211 (
            .O(N__11036),
            .I(N__11029));
    InMux I__2210 (
            .O(N__11035),
            .I(N__11026));
    LocalMux I__2209 (
            .O(N__11032),
            .I(N__11023));
    Odrv4 I__2208 (
            .O(N__11029),
            .I(\DUT.uart_inst0.g1_0 ));
    LocalMux I__2207 (
            .O(N__11026),
            .I(\DUT.uart_inst0.g1_0 ));
    Odrv4 I__2206 (
            .O(N__11023),
            .I(\DUT.uart_inst0.g1_0 ));
    CascadeMux I__2205 (
            .O(N__11016),
            .I(N__11006));
    CascadeMux I__2204 (
            .O(N__11015),
            .I(N__11001));
    CascadeMux I__2203 (
            .O(N__11014),
            .I(N__10998));
    InMux I__2202 (
            .O(N__11013),
            .I(N__10990));
    InMux I__2201 (
            .O(N__11012),
            .I(N__10985));
    InMux I__2200 (
            .O(N__11011),
            .I(N__10985));
    InMux I__2199 (
            .O(N__11010),
            .I(N__10976));
    InMux I__2198 (
            .O(N__11009),
            .I(N__10976));
    InMux I__2197 (
            .O(N__11006),
            .I(N__10976));
    InMux I__2196 (
            .O(N__11005),
            .I(N__10976));
    InMux I__2195 (
            .O(N__11004),
            .I(N__10961));
    InMux I__2194 (
            .O(N__11001),
            .I(N__10961));
    InMux I__2193 (
            .O(N__10998),
            .I(N__10961));
    InMux I__2192 (
            .O(N__10997),
            .I(N__10961));
    InMux I__2191 (
            .O(N__10996),
            .I(N__10961));
    InMux I__2190 (
            .O(N__10995),
            .I(N__10961));
    InMux I__2189 (
            .O(N__10994),
            .I(N__10961));
    CascadeMux I__2188 (
            .O(N__10993),
            .I(N__10956));
    LocalMux I__2187 (
            .O(N__10990),
            .I(N__10949));
    LocalMux I__2186 (
            .O(N__10985),
            .I(N__10946));
    LocalMux I__2185 (
            .O(N__10976),
            .I(N__10941));
    LocalMux I__2184 (
            .O(N__10961),
            .I(N__10941));
    InMux I__2183 (
            .O(N__10960),
            .I(N__10928));
    InMux I__2182 (
            .O(N__10959),
            .I(N__10928));
    InMux I__2181 (
            .O(N__10956),
            .I(N__10928));
    InMux I__2180 (
            .O(N__10955),
            .I(N__10928));
    InMux I__2179 (
            .O(N__10954),
            .I(N__10928));
    InMux I__2178 (
            .O(N__10953),
            .I(N__10928));
    InMux I__2177 (
            .O(N__10952),
            .I(N__10922));
    Span4Mux_h I__2176 (
            .O(N__10949),
            .I(N__10919));
    Span4Mux_h I__2175 (
            .O(N__10946),
            .I(N__10916));
    Span4Mux_v I__2174 (
            .O(N__10941),
            .I(N__10913));
    LocalMux I__2173 (
            .O(N__10928),
            .I(N__10910));
    InMux I__2172 (
            .O(N__10927),
            .I(N__10903));
    InMux I__2171 (
            .O(N__10926),
            .I(N__10903));
    InMux I__2170 (
            .O(N__10925),
            .I(N__10903));
    LocalMux I__2169 (
            .O(N__10922),
            .I(\DUT.uart_inst0.recv_stateZ0Z_0 ));
    Odrv4 I__2168 (
            .O(N__10919),
            .I(\DUT.uart_inst0.recv_stateZ0Z_0 ));
    Odrv4 I__2167 (
            .O(N__10916),
            .I(\DUT.uart_inst0.recv_stateZ0Z_0 ));
    Odrv4 I__2166 (
            .O(N__10913),
            .I(\DUT.uart_inst0.recv_stateZ0Z_0 ));
    Odrv4 I__2165 (
            .O(N__10910),
            .I(\DUT.uart_inst0.recv_stateZ0Z_0 ));
    LocalMux I__2164 (
            .O(N__10903),
            .I(\DUT.uart_inst0.recv_stateZ0Z_0 ));
    CascadeMux I__2163 (
            .O(N__10890),
            .I(N__10886));
    InMux I__2162 (
            .O(N__10889),
            .I(N__10883));
    InMux I__2161 (
            .O(N__10886),
            .I(N__10880));
    LocalMux I__2160 (
            .O(N__10883),
            .I(N__10873));
    LocalMux I__2159 (
            .O(N__10880),
            .I(N__10870));
    InMux I__2158 (
            .O(N__10879),
            .I(N__10865));
    InMux I__2157 (
            .O(N__10878),
            .I(N__10865));
    InMux I__2156 (
            .O(N__10877),
            .I(N__10860));
    InMux I__2155 (
            .O(N__10876),
            .I(N__10860));
    Odrv4 I__2154 (
            .O(N__10873),
            .I(\DUT.uart_inst0.recv_stateZ0Z_5 ));
    Odrv4 I__2153 (
            .O(N__10870),
            .I(\DUT.uart_inst0.recv_stateZ0Z_5 ));
    LocalMux I__2152 (
            .O(N__10865),
            .I(\DUT.uart_inst0.recv_stateZ0Z_5 ));
    LocalMux I__2151 (
            .O(N__10860),
            .I(\DUT.uart_inst0.recv_stateZ0Z_5 ));
    CascadeMux I__2150 (
            .O(N__10851),
            .I(N__10848));
    InMux I__2149 (
            .O(N__10848),
            .I(N__10845));
    LocalMux I__2148 (
            .O(N__10845),
            .I(N__10842));
    Span4Mux_v I__2147 (
            .O(N__10842),
            .I(N__10839));
    Odrv4 I__2146 (
            .O(N__10839),
            .I(\DUT.uart_inst0.rx_countdown_8_i_a2_0_2 ));
    InMux I__2145 (
            .O(N__10836),
            .I(N__10833));
    LocalMux I__2144 (
            .O(N__10833),
            .I(\DUT.uart_inst0.m10_e_3 ));
    InMux I__2143 (
            .O(N__10830),
            .I(N__10827));
    LocalMux I__2142 (
            .O(N__10827),
            .I(\DUT.uart_inst0.m10_e_2 ));
    InMux I__2141 (
            .O(N__10824),
            .I(N__10818));
    CascadeMux I__2140 (
            .O(N__10823),
            .I(N__10815));
    IoInMux I__2139 (
            .O(N__10822),
            .I(N__10809));
    InMux I__2138 (
            .O(N__10821),
            .I(N__10806));
    LocalMux I__2137 (
            .O(N__10818),
            .I(N__10803));
    InMux I__2136 (
            .O(N__10815),
            .I(N__10800));
    InMux I__2135 (
            .O(N__10814),
            .I(N__10795));
    InMux I__2134 (
            .O(N__10813),
            .I(N__10795));
    InMux I__2133 (
            .O(N__10812),
            .I(N__10792));
    LocalMux I__2132 (
            .O(N__10809),
            .I(N__10788));
    LocalMux I__2131 (
            .O(N__10806),
            .I(N__10784));
    Span4Mux_v I__2130 (
            .O(N__10803),
            .I(N__10779));
    LocalMux I__2129 (
            .O(N__10800),
            .I(N__10779));
    LocalMux I__2128 (
            .O(N__10795),
            .I(N__10776));
    LocalMux I__2127 (
            .O(N__10792),
            .I(N__10773));
    InMux I__2126 (
            .O(N__10791),
            .I(N__10770));
    Span4Mux_s1_v I__2125 (
            .O(N__10788),
            .I(N__10767));
    InMux I__2124 (
            .O(N__10787),
            .I(N__10764));
    Span4Mux_v I__2123 (
            .O(N__10784),
            .I(N__10759));
    Span4Mux_v I__2122 (
            .O(N__10779),
            .I(N__10759));
    Span4Mux_h I__2121 (
            .O(N__10776),
            .I(N__10752));
    Span4Mux_v I__2120 (
            .O(N__10773),
            .I(N__10752));
    LocalMux I__2119 (
            .O(N__10770),
            .I(N__10752));
    Span4Mux_v I__2118 (
            .O(N__10767),
            .I(N__10749));
    LocalMux I__2117 (
            .O(N__10764),
            .I(N__10746));
    Sp12to4 I__2116 (
            .O(N__10759),
            .I(N__10743));
    Span4Mux_v I__2115 (
            .O(N__10752),
            .I(N__10740));
    Sp12to4 I__2114 (
            .O(N__10749),
            .I(N__10735));
    Span12Mux_s5_v I__2113 (
            .O(N__10746),
            .I(N__10735));
    Span12Mux_h I__2112 (
            .O(N__10743),
            .I(N__10730));
    Sp12to4 I__2111 (
            .O(N__10740),
            .I(N__10730));
    Span12Mux_h I__2110 (
            .O(N__10735),
            .I(N__10727));
    Span12Mux_h I__2109 (
            .O(N__10730),
            .I(N__10724));
    Span12Mux_v I__2108 (
            .O(N__10727),
            .I(N__10721));
    Span12Mux_v I__2107 (
            .O(N__10724),
            .I(N__10718));
    Odrv12 I__2106 (
            .O(N__10721),
            .I(wPllLocked));
    Odrv12 I__2105 (
            .O(N__10718),
            .I(wPllLocked));
    CascadeMux I__2104 (
            .O(N__10713),
            .I(\DUT.uart_inst0.N_20_mux_cascade_ ));
    InMux I__2103 (
            .O(N__10710),
            .I(N__10703));
    CascadeMux I__2102 (
            .O(N__10709),
            .I(N__10696));
    InMux I__2101 (
            .O(N__10708),
            .I(N__10687));
    InMux I__2100 (
            .O(N__10707),
            .I(N__10687));
    CascadeMux I__2099 (
            .O(N__10706),
            .I(N__10679));
    LocalMux I__2098 (
            .O(N__10703),
            .I(N__10672));
    InMux I__2097 (
            .O(N__10702),
            .I(N__10667));
    InMux I__2096 (
            .O(N__10701),
            .I(N__10667));
    InMux I__2095 (
            .O(N__10700),
            .I(N__10664));
    InMux I__2094 (
            .O(N__10699),
            .I(N__10659));
    InMux I__2093 (
            .O(N__10696),
            .I(N__10659));
    InMux I__2092 (
            .O(N__10695),
            .I(N__10656));
    InMux I__2091 (
            .O(N__10694),
            .I(N__10653));
    InMux I__2090 (
            .O(N__10693),
            .I(N__10648));
    InMux I__2089 (
            .O(N__10692),
            .I(N__10648));
    LocalMux I__2088 (
            .O(N__10687),
            .I(N__10645));
    InMux I__2087 (
            .O(N__10686),
            .I(N__10642));
    InMux I__2086 (
            .O(N__10685),
            .I(N__10637));
    InMux I__2085 (
            .O(N__10684),
            .I(N__10637));
    InMux I__2084 (
            .O(N__10683),
            .I(N__10632));
    InMux I__2083 (
            .O(N__10682),
            .I(N__10632));
    InMux I__2082 (
            .O(N__10679),
            .I(N__10627));
    InMux I__2081 (
            .O(N__10678),
            .I(N__10627));
    InMux I__2080 (
            .O(N__10677),
            .I(N__10622));
    InMux I__2079 (
            .O(N__10676),
            .I(N__10622));
    InMux I__2078 (
            .O(N__10675),
            .I(N__10619));
    Span4Mux_v I__2077 (
            .O(N__10672),
            .I(N__10608));
    LocalMux I__2076 (
            .O(N__10667),
            .I(N__10608));
    LocalMux I__2075 (
            .O(N__10664),
            .I(N__10608));
    LocalMux I__2074 (
            .O(N__10659),
            .I(N__10608));
    LocalMux I__2073 (
            .O(N__10656),
            .I(N__10608));
    LocalMux I__2072 (
            .O(N__10653),
            .I(N__10603));
    LocalMux I__2071 (
            .O(N__10648),
            .I(N__10603));
    Span4Mux_v I__2070 (
            .O(N__10645),
            .I(N__10600));
    LocalMux I__2069 (
            .O(N__10642),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    LocalMux I__2068 (
            .O(N__10637),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    LocalMux I__2067 (
            .O(N__10632),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    LocalMux I__2066 (
            .O(N__10627),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    LocalMux I__2065 (
            .O(N__10622),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    LocalMux I__2064 (
            .O(N__10619),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    Odrv4 I__2063 (
            .O(N__10608),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    Odrv4 I__2062 (
            .O(N__10603),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    Odrv4 I__2061 (
            .O(N__10600),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    CascadeMux I__2060 (
            .O(N__10581),
            .I(\DUT.uart_inst0.m7_3_cascade_ ));
    InMux I__2059 (
            .O(N__10578),
            .I(N__10575));
    LocalMux I__2058 (
            .O(N__10575),
            .I(N__10572));
    Odrv12 I__2057 (
            .O(N__10572),
            .I(\DUT.uart_inst0.N_28_mux ));
    CascadeMux I__2056 (
            .O(N__10569),
            .I(N__10552));
    CascadeMux I__2055 (
            .O(N__10568),
            .I(N__10549));
    CascadeMux I__2054 (
            .O(N__10567),
            .I(N__10544));
    InMux I__2053 (
            .O(N__10566),
            .I(N__10537));
    InMux I__2052 (
            .O(N__10565),
            .I(N__10537));
    InMux I__2051 (
            .O(N__10564),
            .I(N__10537));
    CascadeMux I__2050 (
            .O(N__10563),
            .I(N__10532));
    CascadeMux I__2049 (
            .O(N__10562),
            .I(N__10528));
    CascadeMux I__2048 (
            .O(N__10561),
            .I(N__10523));
    CascadeMux I__2047 (
            .O(N__10560),
            .I(N__10520));
    CascadeMux I__2046 (
            .O(N__10559),
            .I(N__10514));
    CascadeMux I__2045 (
            .O(N__10558),
            .I(N__10510));
    CascadeMux I__2044 (
            .O(N__10557),
            .I(N__10506));
    InMux I__2043 (
            .O(N__10556),
            .I(N__10499));
    InMux I__2042 (
            .O(N__10555),
            .I(N__10494));
    InMux I__2041 (
            .O(N__10552),
            .I(N__10494));
    InMux I__2040 (
            .O(N__10549),
            .I(N__10491));
    InMux I__2039 (
            .O(N__10548),
            .I(N__10488));
    InMux I__2038 (
            .O(N__10547),
            .I(N__10483));
    InMux I__2037 (
            .O(N__10544),
            .I(N__10483));
    LocalMux I__2036 (
            .O(N__10537),
            .I(N__10479));
    InMux I__2035 (
            .O(N__10536),
            .I(N__10474));
    InMux I__2034 (
            .O(N__10535),
            .I(N__10474));
    InMux I__2033 (
            .O(N__10532),
            .I(N__10463));
    InMux I__2032 (
            .O(N__10531),
            .I(N__10463));
    InMux I__2031 (
            .O(N__10528),
            .I(N__10463));
    InMux I__2030 (
            .O(N__10527),
            .I(N__10463));
    InMux I__2029 (
            .O(N__10526),
            .I(N__10463));
    InMux I__2028 (
            .O(N__10523),
            .I(N__10456));
    InMux I__2027 (
            .O(N__10520),
            .I(N__10456));
    InMux I__2026 (
            .O(N__10519),
            .I(N__10456));
    InMux I__2025 (
            .O(N__10518),
            .I(N__10453));
    InMux I__2024 (
            .O(N__10517),
            .I(N__10450));
    InMux I__2023 (
            .O(N__10514),
            .I(N__10443));
    InMux I__2022 (
            .O(N__10513),
            .I(N__10443));
    InMux I__2021 (
            .O(N__10510),
            .I(N__10443));
    InMux I__2020 (
            .O(N__10509),
            .I(N__10430));
    InMux I__2019 (
            .O(N__10506),
            .I(N__10430));
    InMux I__2018 (
            .O(N__10505),
            .I(N__10430));
    InMux I__2017 (
            .O(N__10504),
            .I(N__10430));
    InMux I__2016 (
            .O(N__10503),
            .I(N__10430));
    InMux I__2015 (
            .O(N__10502),
            .I(N__10430));
    LocalMux I__2014 (
            .O(N__10499),
            .I(N__10425));
    LocalMux I__2013 (
            .O(N__10494),
            .I(N__10425));
    LocalMux I__2012 (
            .O(N__10491),
            .I(N__10417));
    LocalMux I__2011 (
            .O(N__10488),
            .I(N__10417));
    LocalMux I__2010 (
            .O(N__10483),
            .I(N__10417));
    CascadeMux I__2009 (
            .O(N__10482),
            .I(N__10414));
    Span4Mux_v I__2008 (
            .O(N__10479),
            .I(N__10409));
    LocalMux I__2007 (
            .O(N__10474),
            .I(N__10409));
    LocalMux I__2006 (
            .O(N__10463),
            .I(N__10406));
    LocalMux I__2005 (
            .O(N__10456),
            .I(N__10403));
    LocalMux I__2004 (
            .O(N__10453),
            .I(N__10400));
    LocalMux I__2003 (
            .O(N__10450),
            .I(N__10393));
    LocalMux I__2002 (
            .O(N__10443),
            .I(N__10393));
    LocalMux I__2001 (
            .O(N__10430),
            .I(N__10393));
    Span4Mux_v I__2000 (
            .O(N__10425),
            .I(N__10390));
    InMux I__1999 (
            .O(N__10424),
            .I(N__10387));
    Span4Mux_v I__1998 (
            .O(N__10417),
            .I(N__10384));
    InMux I__1997 (
            .O(N__10414),
            .I(N__10381));
    Span4Mux_h I__1996 (
            .O(N__10409),
            .I(N__10376));
    Span4Mux_h I__1995 (
            .O(N__10406),
            .I(N__10376));
    Span4Mux_h I__1994 (
            .O(N__10403),
            .I(N__10369));
    Span4Mux_v I__1993 (
            .O(N__10400),
            .I(N__10369));
    Span4Mux_h I__1992 (
            .O(N__10393),
            .I(N__10369));
    Sp12to4 I__1991 (
            .O(N__10390),
            .I(N__10360));
    LocalMux I__1990 (
            .O(N__10387),
            .I(N__10360));
    Sp12to4 I__1989 (
            .O(N__10384),
            .I(N__10360));
    LocalMux I__1988 (
            .O(N__10381),
            .I(N__10360));
    Span4Mux_h I__1987 (
            .O(N__10376),
            .I(N__10357));
    Span4Mux_h I__1986 (
            .O(N__10369),
            .I(N__10354));
    Span12Mux_h I__1985 (
            .O(N__10360),
            .I(N__10351));
    Span4Mux_v I__1984 (
            .O(N__10357),
            .I(N__10348));
    Span4Mux_v I__1983 (
            .O(N__10354),
            .I(N__10345));
    Odrv12 I__1982 (
            .O(N__10351),
            .I(P1A1_c));
    Odrv4 I__1981 (
            .O(N__10348),
            .I(P1A1_c));
    Odrv4 I__1980 (
            .O(N__10345),
            .I(P1A1_c));
    CascadeMux I__1979 (
            .O(N__10338),
            .I(N__10335));
    InMux I__1978 (
            .O(N__10335),
            .I(N__10332));
    LocalMux I__1977 (
            .O(N__10332),
            .I(\DUT.uart_inst0.m2_e_0 ));
    InMux I__1976 (
            .O(N__10329),
            .I(N__10326));
    LocalMux I__1975 (
            .O(N__10326),
            .I(N__10323));
    Span4Mux_v I__1974 (
            .O(N__10323),
            .I(N__10320));
    Odrv4 I__1973 (
            .O(N__10320),
            .I(\DUT.uart_inst0.G_19_0_1 ));
    CascadeMux I__1972 (
            .O(N__10317),
            .I(\DUT.uart_inst0.G_19_0_a5_0_4_cascade_ ));
    InMux I__1971 (
            .O(N__10314),
            .I(N__10310));
    InMux I__1970 (
            .O(N__10313),
            .I(N__10307));
    LocalMux I__1969 (
            .O(N__10310),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_2_0_2 ));
    LocalMux I__1968 (
            .O(N__10307),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_2_0_2 ));
    InMux I__1967 (
            .O(N__10302),
            .I(N__10299));
    LocalMux I__1966 (
            .O(N__10299),
            .I(\DUT.uart_inst0.G_8_i_a3_1 ));
    InMux I__1965 (
            .O(N__10296),
            .I(N__10293));
    LocalMux I__1964 (
            .O(N__10293),
            .I(N__10286));
    InMux I__1963 (
            .O(N__10292),
            .I(N__10283));
    InMux I__1962 (
            .O(N__10291),
            .I(N__10278));
    InMux I__1961 (
            .O(N__10290),
            .I(N__10278));
    InMux I__1960 (
            .O(N__10289),
            .I(N__10268));
    Span4Mux_h I__1959 (
            .O(N__10286),
            .I(N__10261));
    LocalMux I__1958 (
            .O(N__10283),
            .I(N__10261));
    LocalMux I__1957 (
            .O(N__10278),
            .I(N__10261));
    InMux I__1956 (
            .O(N__10277),
            .I(N__10258));
    InMux I__1955 (
            .O(N__10276),
            .I(N__10253));
    InMux I__1954 (
            .O(N__10275),
            .I(N__10253));
    InMux I__1953 (
            .O(N__10274),
            .I(N__10246));
    InMux I__1952 (
            .O(N__10273),
            .I(N__10246));
    InMux I__1951 (
            .O(N__10272),
            .I(N__10246));
    InMux I__1950 (
            .O(N__10271),
            .I(N__10243));
    LocalMux I__1949 (
            .O(N__10268),
            .I(DUT_uart_inst0_rx_countdown_3_s1_4));
    Odrv4 I__1948 (
            .O(N__10261),
            .I(DUT_uart_inst0_rx_countdown_3_s1_4));
    LocalMux I__1947 (
            .O(N__10258),
            .I(DUT_uart_inst0_rx_countdown_3_s1_4));
    LocalMux I__1946 (
            .O(N__10253),
            .I(DUT_uart_inst0_rx_countdown_3_s1_4));
    LocalMux I__1945 (
            .O(N__10246),
            .I(DUT_uart_inst0_rx_countdown_3_s1_4));
    LocalMux I__1944 (
            .O(N__10243),
            .I(DUT_uart_inst0_rx_countdown_3_s1_4));
    InMux I__1943 (
            .O(N__10230),
            .I(N__10225));
    InMux I__1942 (
            .O(N__10229),
            .I(N__10222));
    InMux I__1941 (
            .O(N__10228),
            .I(N__10211));
    LocalMux I__1940 (
            .O(N__10225),
            .I(N__10206));
    LocalMux I__1939 (
            .O(N__10222),
            .I(N__10206));
    InMux I__1938 (
            .O(N__10221),
            .I(N__10201));
    InMux I__1937 (
            .O(N__10220),
            .I(N__10201));
    InMux I__1936 (
            .O(N__10219),
            .I(N__10198));
    InMux I__1935 (
            .O(N__10218),
            .I(N__10193));
    InMux I__1934 (
            .O(N__10217),
            .I(N__10193));
    InMux I__1933 (
            .O(N__10216),
            .I(N__10190));
    InMux I__1932 (
            .O(N__10215),
            .I(N__10185));
    InMux I__1931 (
            .O(N__10214),
            .I(N__10185));
    LocalMux I__1930 (
            .O(N__10211),
            .I(DUT_uart_inst0_rx_countdown_3_s1_5));
    Odrv4 I__1929 (
            .O(N__10206),
            .I(DUT_uart_inst0_rx_countdown_3_s1_5));
    LocalMux I__1928 (
            .O(N__10201),
            .I(DUT_uart_inst0_rx_countdown_3_s1_5));
    LocalMux I__1927 (
            .O(N__10198),
            .I(DUT_uart_inst0_rx_countdown_3_s1_5));
    LocalMux I__1926 (
            .O(N__10193),
            .I(DUT_uart_inst0_rx_countdown_3_s1_5));
    LocalMux I__1925 (
            .O(N__10190),
            .I(DUT_uart_inst0_rx_countdown_3_s1_5));
    LocalMux I__1924 (
            .O(N__10185),
            .I(DUT_uart_inst0_rx_countdown_3_s1_5));
    InMux I__1923 (
            .O(N__10170),
            .I(N__10165));
    CascadeMux I__1922 (
            .O(N__10169),
            .I(N__10160));
    CascadeMux I__1921 (
            .O(N__10168),
            .I(N__10154));
    LocalMux I__1920 (
            .O(N__10165),
            .I(N__10148));
    InMux I__1919 (
            .O(N__10164),
            .I(N__10143));
    InMux I__1918 (
            .O(N__10163),
            .I(N__10143));
    InMux I__1917 (
            .O(N__10160),
            .I(N__10139));
    InMux I__1916 (
            .O(N__10159),
            .I(N__10136));
    InMux I__1915 (
            .O(N__10158),
            .I(N__10129));
    InMux I__1914 (
            .O(N__10157),
            .I(N__10129));
    InMux I__1913 (
            .O(N__10154),
            .I(N__10129));
    InMux I__1912 (
            .O(N__10153),
            .I(N__10122));
    InMux I__1911 (
            .O(N__10152),
            .I(N__10122));
    InMux I__1910 (
            .O(N__10151),
            .I(N__10122));
    Span4Mux_h I__1909 (
            .O(N__10148),
            .I(N__10117));
    LocalMux I__1908 (
            .O(N__10143),
            .I(N__10117));
    InMux I__1907 (
            .O(N__10142),
            .I(N__10114));
    LocalMux I__1906 (
            .O(N__10139),
            .I(DUT_uart_inst0_rx_countdown_3_s1_3));
    LocalMux I__1905 (
            .O(N__10136),
            .I(DUT_uart_inst0_rx_countdown_3_s1_3));
    LocalMux I__1904 (
            .O(N__10129),
            .I(DUT_uart_inst0_rx_countdown_3_s1_3));
    LocalMux I__1903 (
            .O(N__10122),
            .I(DUT_uart_inst0_rx_countdown_3_s1_3));
    Odrv4 I__1902 (
            .O(N__10117),
            .I(DUT_uart_inst0_rx_countdown_3_s1_3));
    LocalMux I__1901 (
            .O(N__10114),
            .I(DUT_uart_inst0_rx_countdown_3_s1_3));
    InMux I__1900 (
            .O(N__10101),
            .I(N__10094));
    CascadeMux I__1899 (
            .O(N__10100),
            .I(N__10090));
    InMux I__1898 (
            .O(N__10099),
            .I(N__10087));
    InMux I__1897 (
            .O(N__10098),
            .I(N__10082));
    InMux I__1896 (
            .O(N__10097),
            .I(N__10082));
    LocalMux I__1895 (
            .O(N__10094),
            .I(N__10077));
    InMux I__1894 (
            .O(N__10093),
            .I(N__10072));
    InMux I__1893 (
            .O(N__10090),
            .I(N__10072));
    LocalMux I__1892 (
            .O(N__10087),
            .I(N__10066));
    LocalMux I__1891 (
            .O(N__10082),
            .I(N__10066));
    InMux I__1890 (
            .O(N__10081),
            .I(N__10061));
    InMux I__1889 (
            .O(N__10080),
            .I(N__10058));
    Span4Mux_v I__1888 (
            .O(N__10077),
            .I(N__10052));
    LocalMux I__1887 (
            .O(N__10072),
            .I(N__10052));
    InMux I__1886 (
            .O(N__10071),
            .I(N__10046));
    Span4Mux_v I__1885 (
            .O(N__10066),
            .I(N__10043));
    InMux I__1884 (
            .O(N__10065),
            .I(N__10038));
    InMux I__1883 (
            .O(N__10064),
            .I(N__10038));
    LocalMux I__1882 (
            .O(N__10061),
            .I(N__10033));
    LocalMux I__1881 (
            .O(N__10058),
            .I(N__10033));
    InMux I__1880 (
            .O(N__10057),
            .I(N__10030));
    Span4Mux_h I__1879 (
            .O(N__10052),
            .I(N__10027));
    InMux I__1878 (
            .O(N__10051),
            .I(N__10022));
    InMux I__1877 (
            .O(N__10050),
            .I(N__10022));
    InMux I__1876 (
            .O(N__10049),
            .I(N__10019));
    LocalMux I__1875 (
            .O(N__10046),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    Odrv4 I__1874 (
            .O(N__10043),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    LocalMux I__1873 (
            .O(N__10038),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    Odrv4 I__1872 (
            .O(N__10033),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    LocalMux I__1871 (
            .O(N__10030),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    Odrv4 I__1870 (
            .O(N__10027),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    LocalMux I__1869 (
            .O(N__10022),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    LocalMux I__1868 (
            .O(N__10019),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    CascadeMux I__1867 (
            .O(N__10002),
            .I(N__9998));
    InMux I__1866 (
            .O(N__10001),
            .I(N__9992));
    InMux I__1865 (
            .O(N__9998),
            .I(N__9989));
    InMux I__1864 (
            .O(N__9997),
            .I(N__9986));
    CascadeMux I__1863 (
            .O(N__9996),
            .I(N__9978));
    CascadeMux I__1862 (
            .O(N__9995),
            .I(N__9974));
    LocalMux I__1861 (
            .O(N__9992),
            .I(N__9969));
    LocalMux I__1860 (
            .O(N__9989),
            .I(N__9969));
    LocalMux I__1859 (
            .O(N__9986),
            .I(N__9966));
    InMux I__1858 (
            .O(N__9985),
            .I(N__9963));
    InMux I__1857 (
            .O(N__9984),
            .I(N__9958));
    InMux I__1856 (
            .O(N__9983),
            .I(N__9958));
    InMux I__1855 (
            .O(N__9982),
            .I(N__9955));
    InMux I__1854 (
            .O(N__9981),
            .I(N__9948));
    InMux I__1853 (
            .O(N__9978),
            .I(N__9948));
    InMux I__1852 (
            .O(N__9977),
            .I(N__9948));
    InMux I__1851 (
            .O(N__9974),
            .I(N__9945));
    Span4Mux_v I__1850 (
            .O(N__9969),
            .I(N__9940));
    Span4Mux_v I__1849 (
            .O(N__9966),
            .I(N__9940));
    LocalMux I__1848 (
            .O(N__9963),
            .I(DUT_uart_inst0_rx_countdown_3_s1_2));
    LocalMux I__1847 (
            .O(N__9958),
            .I(DUT_uart_inst0_rx_countdown_3_s1_2));
    LocalMux I__1846 (
            .O(N__9955),
            .I(DUT_uart_inst0_rx_countdown_3_s1_2));
    LocalMux I__1845 (
            .O(N__9948),
            .I(DUT_uart_inst0_rx_countdown_3_s1_2));
    LocalMux I__1844 (
            .O(N__9945),
            .I(DUT_uart_inst0_rx_countdown_3_s1_2));
    Odrv4 I__1843 (
            .O(N__9940),
            .I(DUT_uart_inst0_rx_countdown_3_s1_2));
    InMux I__1842 (
            .O(N__9927),
            .I(N__9922));
    InMux I__1841 (
            .O(N__9926),
            .I(N__9914));
    InMux I__1840 (
            .O(N__9925),
            .I(N__9914));
    LocalMux I__1839 (
            .O(N__9922),
            .I(N__9910));
    CascadeMux I__1838 (
            .O(N__9921),
            .I(N__9904));
    CascadeMux I__1837 (
            .O(N__9920),
            .I(N__9900));
    InMux I__1836 (
            .O(N__9919),
            .I(N__9896));
    LocalMux I__1835 (
            .O(N__9914),
            .I(N__9893));
    InMux I__1834 (
            .O(N__9913),
            .I(N__9890));
    Span4Mux_v I__1833 (
            .O(N__9910),
            .I(N__9887));
    InMux I__1832 (
            .O(N__9909),
            .I(N__9884));
    InMux I__1831 (
            .O(N__9908),
            .I(N__9881));
    InMux I__1830 (
            .O(N__9907),
            .I(N__9878));
    InMux I__1829 (
            .O(N__9904),
            .I(N__9873));
    InMux I__1828 (
            .O(N__9903),
            .I(N__9873));
    InMux I__1827 (
            .O(N__9900),
            .I(N__9868));
    InMux I__1826 (
            .O(N__9899),
            .I(N__9868));
    LocalMux I__1825 (
            .O(N__9896),
            .I(N__9861));
    Span4Mux_h I__1824 (
            .O(N__9893),
            .I(N__9861));
    LocalMux I__1823 (
            .O(N__9890),
            .I(N__9861));
    Odrv4 I__1822 (
            .O(N__9887),
            .I(DUT_uart_inst0_rx_countdown_3_s1_1));
    LocalMux I__1821 (
            .O(N__9884),
            .I(DUT_uart_inst0_rx_countdown_3_s1_1));
    LocalMux I__1820 (
            .O(N__9881),
            .I(DUT_uart_inst0_rx_countdown_3_s1_1));
    LocalMux I__1819 (
            .O(N__9878),
            .I(DUT_uart_inst0_rx_countdown_3_s1_1));
    LocalMux I__1818 (
            .O(N__9873),
            .I(DUT_uart_inst0_rx_countdown_3_s1_1));
    LocalMux I__1817 (
            .O(N__9868),
            .I(DUT_uart_inst0_rx_countdown_3_s1_1));
    Odrv4 I__1816 (
            .O(N__9861),
            .I(DUT_uart_inst0_rx_countdown_3_s1_1));
    InMux I__1815 (
            .O(N__9846),
            .I(N__9843));
    LocalMux I__1814 (
            .O(N__9843),
            .I(\DUT.uart_inst0.G_19_0_a5_4 ));
    InMux I__1813 (
            .O(N__9840),
            .I(N__9833));
    InMux I__1812 (
            .O(N__9839),
            .I(N__9833));
    InMux I__1811 (
            .O(N__9838),
            .I(N__9830));
    LocalMux I__1810 (
            .O(N__9833),
            .I(N__9827));
    LocalMux I__1809 (
            .O(N__9830),
            .I(N__9822));
    Span4Mux_h I__1808 (
            .O(N__9827),
            .I(N__9822));
    Odrv4 I__1807 (
            .O(N__9822),
            .I(\DUT.uart_inst0.N_44 ));
    InMux I__1806 (
            .O(N__9819),
            .I(N__9816));
    LocalMux I__1805 (
            .O(N__9816),
            .I(N__9813));
    Span4Mux_h I__1804 (
            .O(N__9813),
            .I(N__9810));
    Odrv4 I__1803 (
            .O(N__9810),
            .I(\DUT.uart_inst0.g1_i_a4_1_5 ));
    CascadeMux I__1802 (
            .O(N__9807),
            .I(N__9804));
    InMux I__1801 (
            .O(N__9804),
            .I(N__9801));
    LocalMux I__1800 (
            .O(N__9801),
            .I(\DUT.uart_inst0.g1_i_a4_1_3 ));
    CascadeMux I__1799 (
            .O(N__9798),
            .I(\DUT.uart_inst0.N_78_cascade_ ));
    CascadeMux I__1798 (
            .O(N__9795),
            .I(\DUT.uart_inst0.N_10_mux_cascade_ ));
    InMux I__1797 (
            .O(N__9792),
            .I(N__9789));
    LocalMux I__1796 (
            .O(N__9789),
            .I(\DUT.uart_inst0.P6_mux ));
    CascadeMux I__1795 (
            .O(N__9786),
            .I(\DUT.uart_inst0.G_19_0_a5_0_2_cascade_ ));
    CEMux I__1794 (
            .O(N__9783),
            .I(N__9780));
    LocalMux I__1793 (
            .O(N__9780),
            .I(N__9777));
    Span4Mux_v I__1792 (
            .O(N__9777),
            .I(N__9774));
    Odrv4 I__1791 (
            .O(N__9774),
            .I(\DUT.uart_inst0.rx_bits_remaining_2_sqmuxa ));
    InMux I__1790 (
            .O(N__9771),
            .I(N__9768));
    LocalMux I__1789 (
            .O(N__9768),
            .I(\DUT.uart_inst0.m6_2 ));
    CascadeMux I__1788 (
            .O(N__9765),
            .I(N__9761));
    InMux I__1787 (
            .O(N__9764),
            .I(N__9758));
    InMux I__1786 (
            .O(N__9761),
            .I(N__9755));
    LocalMux I__1785 (
            .O(N__9758),
            .I(N__9749));
    LocalMux I__1784 (
            .O(N__9755),
            .I(N__9749));
    InMux I__1783 (
            .O(N__9754),
            .I(N__9746));
    Span4Mux_v I__1782 (
            .O(N__9749),
            .I(N__9743));
    LocalMux I__1781 (
            .O(N__9746),
            .I(N__9740));
    Odrv4 I__1780 (
            .O(N__9743),
            .I(G_114));
    Odrv12 I__1779 (
            .O(N__9740),
            .I(G_114));
    InMux I__1778 (
            .O(N__9735),
            .I(N__9732));
    LocalMux I__1777 (
            .O(N__9732),
            .I(N__9727));
    InMux I__1776 (
            .O(N__9731),
            .I(N__9724));
    InMux I__1775 (
            .O(N__9730),
            .I(N__9721));
    Odrv4 I__1774 (
            .O(N__9727),
            .I(G_113));
    LocalMux I__1773 (
            .O(N__9724),
            .I(G_113));
    LocalMux I__1772 (
            .O(N__9721),
            .I(G_113));
    CascadeMux I__1771 (
            .O(N__9714),
            .I(\fifo_inst.ftdi_input_inst.un1_rWrStateZ0Z_1_cascade_ ));
    CascadeMux I__1770 (
            .O(N__9711),
            .I(N__9708));
    InMux I__1769 (
            .O(N__9708),
            .I(N__9705));
    LocalMux I__1768 (
            .O(N__9705),
            .I(N__9701));
    InMux I__1767 (
            .O(N__9704),
            .I(N__9698));
    Odrv4 I__1766 (
            .O(N__9701),
            .I(G_118));
    LocalMux I__1765 (
            .O(N__9698),
            .I(G_118));
    CascadeMux I__1764 (
            .O(N__9693),
            .I(G_118_cascade_));
    InMux I__1763 (
            .O(N__9690),
            .I(N__9687));
    LocalMux I__1762 (
            .O(N__9687),
            .I(G_119));
    CascadeMux I__1761 (
            .O(N__9684),
            .I(N__9681));
    InMux I__1760 (
            .O(N__9681),
            .I(N__9678));
    LocalMux I__1759 (
            .O(N__9678),
            .I(N__9673));
    InMux I__1758 (
            .O(N__9677),
            .I(N__9670));
    InMux I__1757 (
            .O(N__9676),
            .I(N__9667));
    Odrv12 I__1756 (
            .O(N__9673),
            .I(G_116));
    LocalMux I__1755 (
            .O(N__9670),
            .I(G_116));
    LocalMux I__1754 (
            .O(N__9667),
            .I(G_116));
    InMux I__1753 (
            .O(N__9660),
            .I(N__9654));
    InMux I__1752 (
            .O(N__9659),
            .I(N__9654));
    LocalMux I__1751 (
            .O(N__9654),
            .I(\fifo_inst.ftdi_input_inst.un1_rWrStateZ0Z_1 ));
    CascadeMux I__1750 (
            .O(N__9651),
            .I(G_116_cascade_));
    CascadeMux I__1749 (
            .O(N__9648),
            .I(N__9645));
    InMux I__1748 (
            .O(N__9645),
            .I(N__9642));
    LocalMux I__1747 (
            .O(N__9642),
            .I(N__9637));
    InMux I__1746 (
            .O(N__9641),
            .I(N__9634));
    InMux I__1745 (
            .O(N__9640),
            .I(N__9631));
    Odrv12 I__1744 (
            .O(N__9637),
            .I(G_117));
    LocalMux I__1743 (
            .O(N__9634),
            .I(G_117));
    LocalMux I__1742 (
            .O(N__9631),
            .I(G_117));
    CascadeMux I__1741 (
            .O(N__9624),
            .I(N__9621));
    InMux I__1740 (
            .O(N__9621),
            .I(N__9618));
    LocalMux I__1739 (
            .O(N__9618),
            .I(N__9615));
    Odrv4 I__1738 (
            .O(N__9615),
            .I(\DUT.rFifoDataror_1 ));
    CascadeMux I__1737 (
            .O(N__9612),
            .I(\DUT.rFifoDataror_1_cascade_ ));
    InMux I__1736 (
            .O(N__9609),
            .I(N__9606));
    LocalMux I__1735 (
            .O(N__9606),
            .I(N__9602));
    InMux I__1734 (
            .O(N__9605),
            .I(N__9599));
    Odrv4 I__1733 (
            .O(N__9602),
            .I(\DUT.rFifoDataror_0_0 ));
    LocalMux I__1732 (
            .O(N__9599),
            .I(\DUT.rFifoDataror_0_0 ));
    InMux I__1731 (
            .O(N__9594),
            .I(N__9573));
    InMux I__1730 (
            .O(N__9593),
            .I(N__9573));
    InMux I__1729 (
            .O(N__9592),
            .I(N__9573));
    InMux I__1728 (
            .O(N__9591),
            .I(N__9573));
    InMux I__1727 (
            .O(N__9590),
            .I(N__9573));
    InMux I__1726 (
            .O(N__9589),
            .I(N__9573));
    InMux I__1725 (
            .O(N__9588),
            .I(N__9573));
    LocalMux I__1724 (
            .O(N__9573),
            .I(\DUT.rFifoDataror_0 ));
    InMux I__1723 (
            .O(N__9570),
            .I(N__9566));
    SRMux I__1722 (
            .O(N__9569),
            .I(N__9563));
    LocalMux I__1721 (
            .O(N__9566),
            .I(N__9560));
    LocalMux I__1720 (
            .O(N__9563),
            .I(N__9557));
    Span4Mux_s3_v I__1719 (
            .O(N__9560),
            .I(N__9551));
    Span4Mux_h I__1718 (
            .O(N__9557),
            .I(N__9551));
    InMux I__1717 (
            .O(N__9556),
            .I(N__9548));
    Odrv4 I__1716 (
            .O(N__9551),
            .I(G_115));
    LocalMux I__1715 (
            .O(N__9548),
            .I(G_115));
    InMux I__1714 (
            .O(N__9543),
            .I(N__9540));
    LocalMux I__1713 (
            .O(N__9540),
            .I(\DUT.rFifoDatarx_5 ));
    InMux I__1712 (
            .O(N__9537),
            .I(N__9534));
    LocalMux I__1711 (
            .O(N__9534),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_5 ));
    InMux I__1710 (
            .O(N__9531),
            .I(N__9528));
    LocalMux I__1709 (
            .O(N__9528),
            .I(N__9525));
    Odrv12 I__1708 (
            .O(N__9525),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_6 ));
    CascadeMux I__1707 (
            .O(N__9522),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_ ));
    InMux I__1706 (
            .O(N__9519),
            .I(N__9516));
    LocalMux I__1705 (
            .O(N__9516),
            .I(\DUT.rFifoDatarx_6 ));
    InMux I__1704 (
            .O(N__9513),
            .I(N__9508));
    InMux I__1703 (
            .O(N__9512),
            .I(N__9505));
    CascadeMux I__1702 (
            .O(N__9511),
            .I(N__9502));
    LocalMux I__1701 (
            .O(N__9508),
            .I(N__9497));
    LocalMux I__1700 (
            .O(N__9505),
            .I(N__9497));
    InMux I__1699 (
            .O(N__9502),
            .I(N__9492));
    Span4Mux_h I__1698 (
            .O(N__9497),
            .I(N__9489));
    InMux I__1697 (
            .O(N__9496),
            .I(N__9484));
    InMux I__1696 (
            .O(N__9495),
            .I(N__9484));
    LocalMux I__1695 (
            .O(N__9492),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_1 ));
    Odrv4 I__1694 (
            .O(N__9489),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_1 ));
    LocalMux I__1693 (
            .O(N__9484),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_1 ));
    InMux I__1692 (
            .O(N__9477),
            .I(N__9473));
    InMux I__1691 (
            .O(N__9476),
            .I(N__9470));
    LocalMux I__1690 (
            .O(N__9473),
            .I(N__9464));
    LocalMux I__1689 (
            .O(N__9470),
            .I(N__9464));
    CascadeMux I__1688 (
            .O(N__9469),
            .I(N__9461));
    Span4Mux_h I__1687 (
            .O(N__9464),
            .I(N__9458));
    InMux I__1686 (
            .O(N__9461),
            .I(N__9452));
    Span4Mux_v I__1685 (
            .O(N__9458),
            .I(N__9449));
    InMux I__1684 (
            .O(N__9457),
            .I(N__9442));
    InMux I__1683 (
            .O(N__9456),
            .I(N__9442));
    InMux I__1682 (
            .O(N__9455),
            .I(N__9442));
    LocalMux I__1681 (
            .O(N__9452),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_0 ));
    Odrv4 I__1680 (
            .O(N__9449),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_0 ));
    LocalMux I__1679 (
            .O(N__9442),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_0 ));
    CascadeMux I__1678 (
            .O(N__9435),
            .I(N__9431));
    CascadeMux I__1677 (
            .O(N__9434),
            .I(N__9426));
    InMux I__1676 (
            .O(N__9431),
            .I(N__9422));
    InMux I__1675 (
            .O(N__9430),
            .I(N__9417));
    InMux I__1674 (
            .O(N__9429),
            .I(N__9417));
    InMux I__1673 (
            .O(N__9426),
            .I(N__9413));
    InMux I__1672 (
            .O(N__9425),
            .I(N__9409));
    LocalMux I__1671 (
            .O(N__9422),
            .I(N__9403));
    LocalMux I__1670 (
            .O(N__9417),
            .I(N__9403));
    InMux I__1669 (
            .O(N__9416),
            .I(N__9400));
    LocalMux I__1668 (
            .O(N__9413),
            .I(N__9394));
    CascadeMux I__1667 (
            .O(N__9412),
            .I(N__9391));
    LocalMux I__1666 (
            .O(N__9409),
            .I(N__9388));
    InMux I__1665 (
            .O(N__9408),
            .I(N__9385));
    Span4Mux_h I__1664 (
            .O(N__9403),
            .I(N__9382));
    LocalMux I__1663 (
            .O(N__9400),
            .I(N__9379));
    InMux I__1662 (
            .O(N__9399),
            .I(N__9374));
    InMux I__1661 (
            .O(N__9398),
            .I(N__9374));
    InMux I__1660 (
            .O(N__9397),
            .I(N__9369));
    Span4Mux_v I__1659 (
            .O(N__9394),
            .I(N__9366));
    InMux I__1658 (
            .O(N__9391),
            .I(N__9363));
    Span4Mux_h I__1657 (
            .O(N__9388),
            .I(N__9360));
    LocalMux I__1656 (
            .O(N__9385),
            .I(N__9351));
    Span4Mux_v I__1655 (
            .O(N__9382),
            .I(N__9351));
    Span4Mux_s2_v I__1654 (
            .O(N__9379),
            .I(N__9351));
    LocalMux I__1653 (
            .O(N__9374),
            .I(N__9351));
    InMux I__1652 (
            .O(N__9373),
            .I(N__9346));
    InMux I__1651 (
            .O(N__9372),
            .I(N__9346));
    LocalMux I__1650 (
            .O(N__9369),
            .I(\DUT.rTransmitZ0 ));
    Odrv4 I__1649 (
            .O(N__9366),
            .I(\DUT.rTransmitZ0 ));
    LocalMux I__1648 (
            .O(N__9363),
            .I(\DUT.rTransmitZ0 ));
    Odrv4 I__1647 (
            .O(N__9360),
            .I(\DUT.rTransmitZ0 ));
    Odrv4 I__1646 (
            .O(N__9351),
            .I(\DUT.rTransmitZ0 ));
    LocalMux I__1645 (
            .O(N__9346),
            .I(\DUT.rTransmitZ0 ));
    InMux I__1644 (
            .O(N__9333),
            .I(N__9329));
    InMux I__1643 (
            .O(N__9332),
            .I(N__9326));
    LocalMux I__1642 (
            .O(N__9329),
            .I(N__9320));
    LocalMux I__1641 (
            .O(N__9326),
            .I(N__9320));
    InMux I__1640 (
            .O(N__9325),
            .I(N__9314));
    Span4Mux_h I__1639 (
            .O(N__9320),
            .I(N__9311));
    InMux I__1638 (
            .O(N__9319),
            .I(N__9304));
    InMux I__1637 (
            .O(N__9318),
            .I(N__9304));
    InMux I__1636 (
            .O(N__9317),
            .I(N__9304));
    LocalMux I__1635 (
            .O(N__9314),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_2 ));
    Odrv4 I__1634 (
            .O(N__9311),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_2 ));
    LocalMux I__1633 (
            .O(N__9304),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_2 ));
    CascadeMux I__1632 (
            .O(N__9297),
            .I(\DUT.fifo_tx_inst.rReadPtr11_cascade_ ));
    CascadeMux I__1631 (
            .O(N__9294),
            .I(\DUT.fifo_tx_inst.un1_i11_2_i_cascade_ ));
    InMux I__1630 (
            .O(N__9291),
            .I(N__9285));
    InMux I__1629 (
            .O(N__9290),
            .I(N__9285));
    LocalMux I__1628 (
            .O(N__9285),
            .I(\DUT.fifo_tx_inst.rReadPtr11 ));
    InMux I__1627 (
            .O(N__9282),
            .I(N__9279));
    LocalMux I__1626 (
            .O(N__9279),
            .I(\DUT.fifo_tx_inst.un1_i11_2_i ));
    CascadeMux I__1625 (
            .O(N__9276),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ));
    InMux I__1624 (
            .O(N__9273),
            .I(N__9270));
    LocalMux I__1623 (
            .O(N__9270),
            .I(N__9267));
    Odrv4 I__1622 (
            .O(N__9267),
            .I(\DUT.rFifoDatarx_0 ));
    InMux I__1621 (
            .O(N__9264),
            .I(N__9261));
    LocalMux I__1620 (
            .O(N__9261),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_0 ));
    InMux I__1619 (
            .O(N__9258),
            .I(N__9255));
    LocalMux I__1618 (
            .O(N__9255),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_1 ));
    CascadeMux I__1617 (
            .O(N__9252),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1_cascade_ ));
    InMux I__1616 (
            .O(N__9249),
            .I(N__9246));
    LocalMux I__1615 (
            .O(N__9246),
            .I(\DUT.rFifoDatarx_1 ));
    CascadeMux I__1614 (
            .O(N__9243),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_ ));
    InMux I__1613 (
            .O(N__9240),
            .I(N__9237));
    LocalMux I__1612 (
            .O(N__9237),
            .I(\DUT.rFifoDatarx_4 ));
    InMux I__1611 (
            .O(N__9234),
            .I(N__9231));
    LocalMux I__1610 (
            .O(N__9231),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_4 ));
    CascadeMux I__1609 (
            .O(N__9228),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ));
    InMux I__1608 (
            .O(N__9225),
            .I(N__9222));
    LocalMux I__1607 (
            .O(N__9222),
            .I(N__9219));
    Odrv4 I__1606 (
            .O(N__9219),
            .I(\DUT.uart_inst0.N_19 ));
    InMux I__1605 (
            .O(N__9216),
            .I(N__9213));
    LocalMux I__1604 (
            .O(N__9213),
            .I(\DUT.uart_inst0.G_8_i_a3_0_0 ));
    CascadeMux I__1603 (
            .O(N__9210),
            .I(N__9207));
    InMux I__1602 (
            .O(N__9207),
            .I(N__9204));
    LocalMux I__1601 (
            .O(N__9204),
            .I(N__9201));
    Span4Mux_h I__1600 (
            .O(N__9201),
            .I(N__9198));
    Odrv4 I__1599 (
            .O(N__9198),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_1_1_2 ));
    CascadeMux I__1598 (
            .O(N__9195),
            .I(N__9174));
    CascadeMux I__1597 (
            .O(N__9194),
            .I(N__9171));
    CascadeMux I__1596 (
            .O(N__9193),
            .I(N__9168));
    CascadeMux I__1595 (
            .O(N__9192),
            .I(N__9165));
    CascadeMux I__1594 (
            .O(N__9191),
            .I(N__9162));
    CascadeMux I__1593 (
            .O(N__9190),
            .I(N__9159));
    CascadeMux I__1592 (
            .O(N__9189),
            .I(N__9156));
    CascadeMux I__1591 (
            .O(N__9188),
            .I(N__9153));
    CascadeMux I__1590 (
            .O(N__9187),
            .I(N__9150));
    CascadeMux I__1589 (
            .O(N__9186),
            .I(N__9147));
    CascadeMux I__1588 (
            .O(N__9185),
            .I(N__9144));
    CascadeMux I__1587 (
            .O(N__9184),
            .I(N__9141));
    CascadeMux I__1586 (
            .O(N__9183),
            .I(N__9138));
    CascadeMux I__1585 (
            .O(N__9182),
            .I(N__9135));
    CascadeMux I__1584 (
            .O(N__9181),
            .I(N__9132));
    CascadeMux I__1583 (
            .O(N__9180),
            .I(N__9129));
    SRMux I__1582 (
            .O(N__9179),
            .I(N__9121));
    InMux I__1581 (
            .O(N__9178),
            .I(N__9116));
    InMux I__1580 (
            .O(N__9177),
            .I(N__9116));
    InMux I__1579 (
            .O(N__9174),
            .I(N__9110));
    InMux I__1578 (
            .O(N__9171),
            .I(N__9101));
    InMux I__1577 (
            .O(N__9168),
            .I(N__9101));
    InMux I__1576 (
            .O(N__9165),
            .I(N__9101));
    InMux I__1575 (
            .O(N__9162),
            .I(N__9101));
    InMux I__1574 (
            .O(N__9159),
            .I(N__9094));
    InMux I__1573 (
            .O(N__9156),
            .I(N__9094));
    InMux I__1572 (
            .O(N__9153),
            .I(N__9094));
    InMux I__1571 (
            .O(N__9150),
            .I(N__9085));
    InMux I__1570 (
            .O(N__9147),
            .I(N__9085));
    InMux I__1569 (
            .O(N__9144),
            .I(N__9085));
    InMux I__1568 (
            .O(N__9141),
            .I(N__9085));
    InMux I__1567 (
            .O(N__9138),
            .I(N__9076));
    InMux I__1566 (
            .O(N__9135),
            .I(N__9076));
    InMux I__1565 (
            .O(N__9132),
            .I(N__9076));
    InMux I__1564 (
            .O(N__9129),
            .I(N__9076));
    CascadeMux I__1563 (
            .O(N__9128),
            .I(N__9073));
    CascadeMux I__1562 (
            .O(N__9127),
            .I(N__9070));
    CascadeMux I__1561 (
            .O(N__9126),
            .I(N__9067));
    CascadeMux I__1560 (
            .O(N__9125),
            .I(N__9064));
    CascadeMux I__1559 (
            .O(N__9124),
            .I(N__9061));
    LocalMux I__1558 (
            .O(N__9121),
            .I(N__9051));
    LocalMux I__1557 (
            .O(N__9116),
            .I(N__9048));
    InMux I__1556 (
            .O(N__9115),
            .I(N__9041));
    InMux I__1555 (
            .O(N__9114),
            .I(N__9041));
    InMux I__1554 (
            .O(N__9113),
            .I(N__9041));
    LocalMux I__1553 (
            .O(N__9110),
            .I(N__9034));
    LocalMux I__1552 (
            .O(N__9101),
            .I(N__9034));
    LocalMux I__1551 (
            .O(N__9094),
            .I(N__9034));
    LocalMux I__1550 (
            .O(N__9085),
            .I(N__9029));
    LocalMux I__1549 (
            .O(N__9076),
            .I(N__9029));
    InMux I__1548 (
            .O(N__9073),
            .I(N__9024));
    InMux I__1547 (
            .O(N__9070),
            .I(N__9024));
    InMux I__1546 (
            .O(N__9067),
            .I(N__9017));
    InMux I__1545 (
            .O(N__9064),
            .I(N__9017));
    InMux I__1544 (
            .O(N__9061),
            .I(N__9017));
    CascadeMux I__1543 (
            .O(N__9060),
            .I(N__9014));
    CascadeMux I__1542 (
            .O(N__9059),
            .I(N__9011));
    CascadeMux I__1541 (
            .O(N__9058),
            .I(N__9008));
    CascadeMux I__1540 (
            .O(N__9057),
            .I(N__9005));
    CascadeMux I__1539 (
            .O(N__9056),
            .I(N__9002));
    CascadeMux I__1538 (
            .O(N__9055),
            .I(N__8999));
    CascadeMux I__1537 (
            .O(N__9054),
            .I(N__8996));
    Span4Mux_v I__1536 (
            .O(N__9051),
            .I(N__8993));
    Span4Mux_h I__1535 (
            .O(N__9048),
            .I(N__8990));
    LocalMux I__1534 (
            .O(N__9041),
            .I(N__8987));
    Span4Mux_v I__1533 (
            .O(N__9034),
            .I(N__8978));
    Span4Mux_v I__1532 (
            .O(N__9029),
            .I(N__8978));
    LocalMux I__1531 (
            .O(N__9024),
            .I(N__8978));
    LocalMux I__1530 (
            .O(N__9017),
            .I(N__8978));
    InMux I__1529 (
            .O(N__9014),
            .I(N__8971));
    InMux I__1528 (
            .O(N__9011),
            .I(N__8971));
    InMux I__1527 (
            .O(N__9008),
            .I(N__8971));
    InMux I__1526 (
            .O(N__9005),
            .I(N__8962));
    InMux I__1525 (
            .O(N__9002),
            .I(N__8962));
    InMux I__1524 (
            .O(N__8999),
            .I(N__8962));
    InMux I__1523 (
            .O(N__8996),
            .I(N__8962));
    Span4Mux_h I__1522 (
            .O(N__8993),
            .I(N__8955));
    Span4Mux_v I__1521 (
            .O(N__8990),
            .I(N__8955));
    Span4Mux_v I__1520 (
            .O(N__8987),
            .I(N__8955));
    Span4Mux_v I__1519 (
            .O(N__8978),
            .I(N__8948));
    LocalMux I__1518 (
            .O(N__8971),
            .I(N__8948));
    LocalMux I__1517 (
            .O(N__8962),
            .I(N__8948));
    Odrv4 I__1516 (
            .O(N__8955),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__1515 (
            .O(N__8948),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__1514 (
            .O(N__8943),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_ ));
    InMux I__1513 (
            .O(N__8940),
            .I(N__8937));
    LocalMux I__1512 (
            .O(N__8937),
            .I(\DUT.rFifoDatarx_7 ));
    InMux I__1511 (
            .O(N__8934),
            .I(N__8931));
    LocalMux I__1510 (
            .O(N__8931),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_7 ));
    InMux I__1509 (
            .O(N__8928),
            .I(N__8925));
    LocalMux I__1508 (
            .O(N__8925),
            .I(\DUT.uart_inst0.m6_1 ));
    InMux I__1507 (
            .O(N__8922),
            .I(N__8916));
    InMux I__1506 (
            .O(N__8921),
            .I(N__8916));
    LocalMux I__1505 (
            .O(N__8916),
            .I(\DUT.uart_inst0.N_7 ));
    InMux I__1504 (
            .O(N__8913),
            .I(N__8910));
    LocalMux I__1503 (
            .O(N__8910),
            .I(\DUT.uart_inst0.recv_state_srsts_1_5 ));
    InMux I__1502 (
            .O(N__8907),
            .I(N__8902));
    InMux I__1501 (
            .O(N__8906),
            .I(N__8897));
    InMux I__1500 (
            .O(N__8905),
            .I(N__8897));
    LocalMux I__1499 (
            .O(N__8902),
            .I(N__8894));
    LocalMux I__1498 (
            .O(N__8897),
            .I(N__8891));
    Span4Mux_v I__1497 (
            .O(N__8894),
            .I(N__8888));
    Odrv4 I__1496 (
            .O(N__8891),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_2_2 ));
    Odrv4 I__1495 (
            .O(N__8888),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_2_2 ));
    CascadeMux I__1494 (
            .O(N__8883),
            .I(\DUT.uart_inst0.recv_state_srsts_1_5_cascade_ ));
    InMux I__1493 (
            .O(N__8880),
            .I(N__8877));
    LocalMux I__1492 (
            .O(N__8877),
            .I(\DUT.uart_inst0.recv_state_srsts_1_4 ));
    InMux I__1491 (
            .O(N__8874),
            .I(N__8870));
    InMux I__1490 (
            .O(N__8873),
            .I(N__8860));
    LocalMux I__1489 (
            .O(N__8870),
            .I(N__8857));
    InMux I__1488 (
            .O(N__8869),
            .I(N__8854));
    InMux I__1487 (
            .O(N__8868),
            .I(N__8847));
    InMux I__1486 (
            .O(N__8867),
            .I(N__8847));
    InMux I__1485 (
            .O(N__8866),
            .I(N__8847));
    InMux I__1484 (
            .O(N__8865),
            .I(N__8840));
    InMux I__1483 (
            .O(N__8864),
            .I(N__8840));
    InMux I__1482 (
            .O(N__8863),
            .I(N__8840));
    LocalMux I__1481 (
            .O(N__8860),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    Odrv4 I__1480 (
            .O(N__8857),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    LocalMux I__1479 (
            .O(N__8854),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    LocalMux I__1478 (
            .O(N__8847),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    LocalMux I__1477 (
            .O(N__8840),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    CascadeMux I__1476 (
            .O(N__8829),
            .I(\DUT.uart_inst0.N_43_cascade_ ));
    CEMux I__1475 (
            .O(N__8826),
            .I(N__8822));
    CEMux I__1474 (
            .O(N__8825),
            .I(N__8819));
    LocalMux I__1473 (
            .O(N__8822),
            .I(N__8816));
    LocalMux I__1472 (
            .O(N__8819),
            .I(\DUT.uart_inst0.recv_state_RNIL139CZ0Z_1 ));
    Odrv4 I__1471 (
            .O(N__8816),
            .I(\DUT.uart_inst0.recv_state_RNIL139CZ0Z_1 ));
    CascadeMux I__1470 (
            .O(N__8811),
            .I(\DUT.uart_inst0.m3_e_1_cascade_ ));
    CascadeMux I__1469 (
            .O(N__8808),
            .I(N__8805));
    InMux I__1468 (
            .O(N__8805),
            .I(N__8802));
    LocalMux I__1467 (
            .O(N__8802),
            .I(N__8795));
    InMux I__1466 (
            .O(N__8801),
            .I(N__8792));
    InMux I__1465 (
            .O(N__8800),
            .I(N__8789));
    InMux I__1464 (
            .O(N__8799),
            .I(N__8780));
    InMux I__1463 (
            .O(N__8798),
            .I(N__8777));
    Span4Mux_h I__1462 (
            .O(N__8795),
            .I(N__8770));
    LocalMux I__1461 (
            .O(N__8792),
            .I(N__8770));
    LocalMux I__1460 (
            .O(N__8789),
            .I(N__8770));
    InMux I__1459 (
            .O(N__8788),
            .I(N__8765));
    InMux I__1458 (
            .O(N__8787),
            .I(N__8765));
    InMux I__1457 (
            .O(N__8786),
            .I(N__8762));
    InMux I__1456 (
            .O(N__8785),
            .I(N__8755));
    InMux I__1455 (
            .O(N__8784),
            .I(N__8755));
    InMux I__1454 (
            .O(N__8783),
            .I(N__8755));
    LocalMux I__1453 (
            .O(N__8780),
            .I(DUT_uart_inst0_recv_state_2));
    LocalMux I__1452 (
            .O(N__8777),
            .I(DUT_uart_inst0_recv_state_2));
    Odrv4 I__1451 (
            .O(N__8770),
            .I(DUT_uart_inst0_recv_state_2));
    LocalMux I__1450 (
            .O(N__8765),
            .I(DUT_uart_inst0_recv_state_2));
    LocalMux I__1449 (
            .O(N__8762),
            .I(DUT_uart_inst0_recv_state_2));
    LocalMux I__1448 (
            .O(N__8755),
            .I(DUT_uart_inst0_recv_state_2));
    InMux I__1447 (
            .O(N__8742),
            .I(N__8732));
    InMux I__1446 (
            .O(N__8741),
            .I(N__8732));
    InMux I__1445 (
            .O(N__8740),
            .I(N__8732));
    CascadeMux I__1444 (
            .O(N__8739),
            .I(N__8726));
    LocalMux I__1443 (
            .O(N__8732),
            .I(N__8723));
    InMux I__1442 (
            .O(N__8731),
            .I(N__8714));
    InMux I__1441 (
            .O(N__8730),
            .I(N__8714));
    InMux I__1440 (
            .O(N__8729),
            .I(N__8714));
    InMux I__1439 (
            .O(N__8726),
            .I(N__8714));
    Odrv12 I__1438 (
            .O(N__8723),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_2 ));
    LocalMux I__1437 (
            .O(N__8714),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_2 ));
    InMux I__1436 (
            .O(N__8709),
            .I(N__8704));
    InMux I__1435 (
            .O(N__8708),
            .I(N__8699));
    InMux I__1434 (
            .O(N__8707),
            .I(N__8699));
    LocalMux I__1433 (
            .O(N__8704),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_3 ));
    LocalMux I__1432 (
            .O(N__8699),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_3 ));
    CascadeMux I__1431 (
            .O(N__8694),
            .I(N__8689));
    InMux I__1430 (
            .O(N__8693),
            .I(N__8683));
    InMux I__1429 (
            .O(N__8692),
            .I(N__8683));
    InMux I__1428 (
            .O(N__8689),
            .I(N__8680));
    CascadeMux I__1427 (
            .O(N__8688),
            .I(N__8673));
    LocalMux I__1426 (
            .O(N__8683),
            .I(N__8668));
    LocalMux I__1425 (
            .O(N__8680),
            .I(N__8668));
    InMux I__1424 (
            .O(N__8679),
            .I(N__8663));
    InMux I__1423 (
            .O(N__8678),
            .I(N__8663));
    InMux I__1422 (
            .O(N__8677),
            .I(N__8656));
    InMux I__1421 (
            .O(N__8676),
            .I(N__8656));
    InMux I__1420 (
            .O(N__8673),
            .I(N__8656));
    Odrv4 I__1419 (
            .O(N__8668),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_1 ));
    LocalMux I__1418 (
            .O(N__8663),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_1 ));
    LocalMux I__1417 (
            .O(N__8656),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_1 ));
    InMux I__1416 (
            .O(N__8649),
            .I(N__8640));
    InMux I__1415 (
            .O(N__8648),
            .I(N__8640));
    InMux I__1414 (
            .O(N__8647),
            .I(N__8640));
    LocalMux I__1413 (
            .O(N__8640),
            .I(N__8634));
    InMux I__1412 (
            .O(N__8639),
            .I(N__8631));
    InMux I__1411 (
            .O(N__8638),
            .I(N__8626));
    InMux I__1410 (
            .O(N__8637),
            .I(N__8626));
    Odrv4 I__1409 (
            .O(N__8634),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_0 ));
    LocalMux I__1408 (
            .O(N__8631),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_0 ));
    LocalMux I__1407 (
            .O(N__8626),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_0 ));
    InMux I__1406 (
            .O(N__8619),
            .I(N__8616));
    LocalMux I__1405 (
            .O(N__8616),
            .I(N__8613));
    Span4Mux_v I__1404 (
            .O(N__8613),
            .I(N__8610));
    Odrv4 I__1403 (
            .O(N__8610),
            .I(\DUT.uart_inst0.recv_state_RNO_4Z0Z_2 ));
    CascadeMux I__1402 (
            .O(N__8607),
            .I(\DUT.uart_inst0.N_21_cascade_ ));
    CascadeMux I__1401 (
            .O(N__8604),
            .I(\DUT.uart_inst0.N_21_mux_cascade_ ));
    InMux I__1400 (
            .O(N__8601),
            .I(N__8598));
    LocalMux I__1399 (
            .O(N__8598),
            .I(\DUT.uart_inst0.N_19_mux ));
    CascadeMux I__1398 (
            .O(N__8595),
            .I(\DUT.uart_inst0.N_13_cascade_ ));
    InMux I__1397 (
            .O(N__8592),
            .I(N__8589));
    LocalMux I__1396 (
            .O(N__8589),
            .I(\DUT.uart_inst0.N_13_0 ));
    CascadeMux I__1395 (
            .O(N__8586),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_2_0_2_cascade_ ));
    InMux I__1394 (
            .O(N__8583),
            .I(N__8580));
    LocalMux I__1393 (
            .O(N__8580),
            .I(\DUT.fifo_tx_inst.un1_i11_i ));
    InMux I__1392 (
            .O(N__8577),
            .I(N__8574));
    LocalMux I__1391 (
            .O(N__8574),
            .I(N__8571));
    Odrv4 I__1390 (
            .O(N__8571),
            .I(\DUT.uart_inst0.g0_0 ));
    InMux I__1389 (
            .O(N__8568),
            .I(N__8565));
    LocalMux I__1388 (
            .O(N__8565),
            .I(\DUT.uart_inst0.N_49 ));
    InMux I__1387 (
            .O(N__8562),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_0_s1 ));
    InMux I__1386 (
            .O(N__8559),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_1_s1 ));
    InMux I__1385 (
            .O(N__8556),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_2_s1 ));
    InMux I__1384 (
            .O(N__8553),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_3_s1 ));
    InMux I__1383 (
            .O(N__8550),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_4_s1 ));
    InMux I__1382 (
            .O(N__8547),
            .I(N__8544));
    LocalMux I__1381 (
            .O(N__8544),
            .I(N__8540));
    InMux I__1380 (
            .O(N__8543),
            .I(N__8537));
    Span4Mux_s1_v I__1379 (
            .O(N__8540),
            .I(N__8533));
    LocalMux I__1378 (
            .O(N__8537),
            .I(N__8530));
    InMux I__1377 (
            .O(N__8536),
            .I(N__8527));
    Span4Mux_v I__1376 (
            .O(N__8533),
            .I(N__8524));
    Span12Mux_s8_v I__1375 (
            .O(N__8530),
            .I(N__8521));
    LocalMux I__1374 (
            .O(N__8527),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_0 ));
    Odrv4 I__1373 (
            .O(N__8524),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_0 ));
    Odrv12 I__1372 (
            .O(N__8521),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_0 ));
    SRMux I__1371 (
            .O(N__8514),
            .I(N__8510));
    SRMux I__1370 (
            .O(N__8513),
            .I(N__8506));
    LocalMux I__1369 (
            .O(N__8510),
            .I(N__8503));
    SRMux I__1368 (
            .O(N__8509),
            .I(N__8500));
    LocalMux I__1367 (
            .O(N__8506),
            .I(N__8497));
    Span4Mux_s1_v I__1366 (
            .O(N__8503),
            .I(N__8492));
    LocalMux I__1365 (
            .O(N__8500),
            .I(N__8492));
    Span4Mux_h I__1364 (
            .O(N__8497),
            .I(N__8489));
    Span4Mux_v I__1363 (
            .O(N__8492),
            .I(N__8486));
    Span4Mux_v I__1362 (
            .O(N__8489),
            .I(N__8483));
    Span4Mux_s1_v I__1361 (
            .O(N__8486),
            .I(N__8480));
    Odrv4 I__1360 (
            .O(N__8483),
            .I(\DUT.uart_inst0.N_20 ));
    Odrv4 I__1359 (
            .O(N__8480),
            .I(\DUT.uart_inst0.N_20 ));
    InMux I__1358 (
            .O(N__8475),
            .I(N__8472));
    LocalMux I__1357 (
            .O(N__8472),
            .I(N__8469));
    Span4Mux_h I__1356 (
            .O(N__8469),
            .I(N__8466));
    Odrv4 I__1355 (
            .O(N__8466),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO ));
    InMux I__1354 (
            .O(N__8463),
            .I(N__8459));
    CascadeMux I__1353 (
            .O(N__8462),
            .I(N__8455));
    LocalMux I__1352 (
            .O(N__8459),
            .I(N__8452));
    InMux I__1351 (
            .O(N__8458),
            .I(N__8447));
    InMux I__1350 (
            .O(N__8455),
            .I(N__8447));
    Odrv4 I__1349 (
            .O(N__8452),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_4 ));
    LocalMux I__1348 (
            .O(N__8447),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_4 ));
    CascadeMux I__1347 (
            .O(N__8442),
            .I(\DUT.uart_inst0.m6_3_cascade_ ));
    CascadeMux I__1346 (
            .O(N__8439),
            .I(\top_pll_inst.m12_1_1_cascade_ ));
    InMux I__1345 (
            .O(N__8436),
            .I(N__8433));
    LocalMux I__1344 (
            .O(N__8433),
            .I(\DUT.uart_inst0.G_30_1 ));
    CascadeMux I__1343 (
            .O(N__8430),
            .I(P18_mux_cascade_));
    InMux I__1342 (
            .O(N__8427),
            .I(N__8424));
    LocalMux I__1341 (
            .O(N__8424),
            .I(N__8421));
    Odrv4 I__1340 (
            .O(N__8421),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_11 ));
    InMux I__1339 (
            .O(N__8418),
            .I(N__8415));
    LocalMux I__1338 (
            .O(N__8415),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_10 ));
    CascadeMux I__1337 (
            .O(N__8412),
            .I(N__8409));
    InMux I__1336 (
            .O(N__8409),
            .I(N__8406));
    LocalMux I__1335 (
            .O(N__8406),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_12 ));
    InMux I__1334 (
            .O(N__8403),
            .I(N__8400));
    LocalMux I__1333 (
            .O(N__8400),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_13 ));
    CascadeMux I__1332 (
            .O(N__8397),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0_cascade_ ));
    InMux I__1331 (
            .O(N__8394),
            .I(N__8387));
    CascadeMux I__1330 (
            .O(N__8393),
            .I(N__8383));
    CascadeMux I__1329 (
            .O(N__8392),
            .I(N__8379));
    CascadeMux I__1328 (
            .O(N__8391),
            .I(N__8376));
    InMux I__1327 (
            .O(N__8390),
            .I(N__8373));
    LocalMux I__1326 (
            .O(N__8387),
            .I(N__8370));
    CascadeMux I__1325 (
            .O(N__8386),
            .I(N__8366));
    InMux I__1324 (
            .O(N__8383),
            .I(N__8358));
    InMux I__1323 (
            .O(N__8382),
            .I(N__8355));
    InMux I__1322 (
            .O(N__8379),
            .I(N__8352));
    InMux I__1321 (
            .O(N__8376),
            .I(N__8349));
    LocalMux I__1320 (
            .O(N__8373),
            .I(N__8344));
    Span4Mux_s2_v I__1319 (
            .O(N__8370),
            .I(N__8344));
    InMux I__1318 (
            .O(N__8369),
            .I(N__8341));
    InMux I__1317 (
            .O(N__8366),
            .I(N__8334));
    InMux I__1316 (
            .O(N__8365),
            .I(N__8334));
    InMux I__1315 (
            .O(N__8364),
            .I(N__8334));
    InMux I__1314 (
            .O(N__8363),
            .I(N__8327));
    InMux I__1313 (
            .O(N__8362),
            .I(N__8327));
    InMux I__1312 (
            .O(N__8361),
            .I(N__8327));
    LocalMux I__1311 (
            .O(N__8358),
            .I(\DUT.tx_state_1 ));
    LocalMux I__1310 (
            .O(N__8355),
            .I(\DUT.tx_state_1 ));
    LocalMux I__1309 (
            .O(N__8352),
            .I(\DUT.tx_state_1 ));
    LocalMux I__1308 (
            .O(N__8349),
            .I(\DUT.tx_state_1 ));
    Odrv4 I__1307 (
            .O(N__8344),
            .I(\DUT.tx_state_1 ));
    LocalMux I__1306 (
            .O(N__8341),
            .I(\DUT.tx_state_1 ));
    LocalMux I__1305 (
            .O(N__8334),
            .I(\DUT.tx_state_1 ));
    LocalMux I__1304 (
            .O(N__8327),
            .I(\DUT.tx_state_1 ));
    CascadeMux I__1303 (
            .O(N__8310),
            .I(\DUT.N_114_cascade_ ));
    CascadeMux I__1302 (
            .O(N__8307),
            .I(N__8304));
    InMux I__1301 (
            .O(N__8304),
            .I(N__8294));
    InMux I__1300 (
            .O(N__8303),
            .I(N__8289));
    InMux I__1299 (
            .O(N__8302),
            .I(N__8289));
    CascadeMux I__1298 (
            .O(N__8301),
            .I(N__8286));
    InMux I__1297 (
            .O(N__8300),
            .I(N__8283));
    CascadeMux I__1296 (
            .O(N__8299),
            .I(N__8280));
    CascadeMux I__1295 (
            .O(N__8298),
            .I(N__8274));
    CascadeMux I__1294 (
            .O(N__8297),
            .I(N__8269));
    LocalMux I__1293 (
            .O(N__8294),
            .I(N__8256));
    LocalMux I__1292 (
            .O(N__8289),
            .I(N__8253));
    InMux I__1291 (
            .O(N__8286),
            .I(N__8247));
    LocalMux I__1290 (
            .O(N__8283),
            .I(N__8244));
    InMux I__1289 (
            .O(N__8280),
            .I(N__8239));
    InMux I__1288 (
            .O(N__8279),
            .I(N__8239));
    InMux I__1287 (
            .O(N__8278),
            .I(N__8236));
    InMux I__1286 (
            .O(N__8277),
            .I(N__8233));
    InMux I__1285 (
            .O(N__8274),
            .I(N__8228));
    InMux I__1284 (
            .O(N__8273),
            .I(N__8228));
    InMux I__1283 (
            .O(N__8272),
            .I(N__8223));
    InMux I__1282 (
            .O(N__8269),
            .I(N__8223));
    InMux I__1281 (
            .O(N__8268),
            .I(N__8218));
    InMux I__1280 (
            .O(N__8267),
            .I(N__8218));
    InMux I__1279 (
            .O(N__8266),
            .I(N__8201));
    InMux I__1278 (
            .O(N__8265),
            .I(N__8201));
    InMux I__1277 (
            .O(N__8264),
            .I(N__8201));
    InMux I__1276 (
            .O(N__8263),
            .I(N__8201));
    InMux I__1275 (
            .O(N__8262),
            .I(N__8201));
    InMux I__1274 (
            .O(N__8261),
            .I(N__8201));
    InMux I__1273 (
            .O(N__8260),
            .I(N__8201));
    InMux I__1272 (
            .O(N__8259),
            .I(N__8201));
    Span4Mux_s3_v I__1271 (
            .O(N__8256),
            .I(N__8196));
    Span4Mux_h I__1270 (
            .O(N__8253),
            .I(N__8196));
    InMux I__1269 (
            .O(N__8252),
            .I(N__8189));
    InMux I__1268 (
            .O(N__8251),
            .I(N__8189));
    InMux I__1267 (
            .O(N__8250),
            .I(N__8189));
    LocalMux I__1266 (
            .O(N__8247),
            .I(N__8182));
    Span4Mux_s2_v I__1265 (
            .O(N__8244),
            .I(N__8182));
    LocalMux I__1264 (
            .O(N__8239),
            .I(N__8182));
    LocalMux I__1263 (
            .O(N__8236),
            .I(\DUT.tx_state_0 ));
    LocalMux I__1262 (
            .O(N__8233),
            .I(\DUT.tx_state_0 ));
    LocalMux I__1261 (
            .O(N__8228),
            .I(\DUT.tx_state_0 ));
    LocalMux I__1260 (
            .O(N__8223),
            .I(\DUT.tx_state_0 ));
    LocalMux I__1259 (
            .O(N__8218),
            .I(\DUT.tx_state_0 ));
    LocalMux I__1258 (
            .O(N__8201),
            .I(\DUT.tx_state_0 ));
    Odrv4 I__1257 (
            .O(N__8196),
            .I(\DUT.tx_state_0 ));
    LocalMux I__1256 (
            .O(N__8189),
            .I(\DUT.tx_state_0 ));
    Odrv4 I__1255 (
            .O(N__8182),
            .I(\DUT.tx_state_0 ));
    CascadeMux I__1254 (
            .O(N__8163),
            .I(N__8160));
    InMux I__1253 (
            .O(N__8160),
            .I(N__8157));
    LocalMux I__1252 (
            .O(N__8157),
            .I(N__8152));
    InMux I__1251 (
            .O(N__8156),
            .I(N__8149));
    InMux I__1250 (
            .O(N__8155),
            .I(N__8146));
    Odrv4 I__1249 (
            .O(N__8152),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_16 ));
    LocalMux I__1248 (
            .O(N__8149),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_16 ));
    LocalMux I__1247 (
            .O(N__8146),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_16 ));
    CascadeMux I__1246 (
            .O(N__8139),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_9_cascade_ ));
    CascadeMux I__1245 (
            .O(N__8136),
            .I(N__8133));
    InMux I__1244 (
            .O(N__8133),
            .I(N__8130));
    LocalMux I__1243 (
            .O(N__8130),
            .I(N__8125));
    InMux I__1242 (
            .O(N__8129),
            .I(N__8120));
    InMux I__1241 (
            .O(N__8128),
            .I(N__8120));
    Odrv4 I__1240 (
            .O(N__8125),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_1 ));
    LocalMux I__1239 (
            .O(N__8120),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_1 ));
    InMux I__1238 (
            .O(N__8115),
            .I(N__8112));
    LocalMux I__1237 (
            .O(N__8112),
            .I(N__8109));
    Odrv4 I__1236 (
            .O(N__8109),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO ));
    InMux I__1235 (
            .O(N__8106),
            .I(N__8103));
    LocalMux I__1234 (
            .O(N__8103),
            .I(N__8098));
    InMux I__1233 (
            .O(N__8102),
            .I(N__8093));
    InMux I__1232 (
            .O(N__8101),
            .I(N__8093));
    Odrv4 I__1231 (
            .O(N__8098),
            .I(\DUT.uart_inst0.rx_clk_dividerZ1Z_1 ));
    LocalMux I__1230 (
            .O(N__8093),
            .I(\DUT.uart_inst0.rx_clk_dividerZ1Z_1 ));
    InMux I__1229 (
            .O(N__8088),
            .I(N__8085));
    LocalMux I__1228 (
            .O(N__8085),
            .I(N__8082));
    Odrv4 I__1227 (
            .O(N__8082),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO ));
    InMux I__1226 (
            .O(N__8079),
            .I(N__8076));
    LocalMux I__1225 (
            .O(N__8076),
            .I(N__8071));
    InMux I__1224 (
            .O(N__8075),
            .I(N__8066));
    InMux I__1223 (
            .O(N__8074),
            .I(N__8066));
    Odrv4 I__1222 (
            .O(N__8071),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_2 ));
    LocalMux I__1221 (
            .O(N__8066),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_2 ));
    InMux I__1220 (
            .O(N__8061),
            .I(N__8058));
    LocalMux I__1219 (
            .O(N__8058),
            .I(N__8055));
    Odrv12 I__1218 (
            .O(N__8055),
            .I(\DUT.uart_inst0.rx_clk_divider_1_3 ));
    InMux I__1217 (
            .O(N__8052),
            .I(N__8049));
    LocalMux I__1216 (
            .O(N__8049),
            .I(N__8045));
    InMux I__1215 (
            .O(N__8048),
            .I(N__8042));
    Odrv4 I__1214 (
            .O(N__8045),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_3 ));
    LocalMux I__1213 (
            .O(N__8042),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_3 ));
    CascadeMux I__1212 (
            .O(N__8037),
            .I(N__8034));
    InMux I__1211 (
            .O(N__8034),
            .I(N__8031));
    LocalMux I__1210 (
            .O(N__8031),
            .I(\DUT.uart_inst0.tx_dataZ0Z_1 ));
    CascadeMux I__1209 (
            .O(N__8028),
            .I(N__8025));
    InMux I__1208 (
            .O(N__8025),
            .I(N__8022));
    LocalMux I__1207 (
            .O(N__8022),
            .I(\DUT.uart_inst0.tx_dataZ0Z_2 ));
    CascadeMux I__1206 (
            .O(N__8019),
            .I(N__8016));
    InMux I__1205 (
            .O(N__8016),
            .I(N__8013));
    LocalMux I__1204 (
            .O(N__8013),
            .I(N__8010));
    Odrv4 I__1203 (
            .O(N__8010),
            .I(\DUT.uart_inst0.tx_dataZ0Z_3 ));
    CascadeMux I__1202 (
            .O(N__8007),
            .I(N__8004));
    InMux I__1201 (
            .O(N__8004),
            .I(N__8001));
    LocalMux I__1200 (
            .O(N__8001),
            .I(\DUT.uart_inst0.tx_dataZ0Z_4 ));
    CascadeMux I__1199 (
            .O(N__7998),
            .I(N__7995));
    InMux I__1198 (
            .O(N__7995),
            .I(N__7992));
    LocalMux I__1197 (
            .O(N__7992),
            .I(\DUT.uart_inst0.tx_dataZ0Z_5 ));
    CascadeMux I__1196 (
            .O(N__7989),
            .I(N__7986));
    InMux I__1195 (
            .O(N__7986),
            .I(N__7983));
    LocalMux I__1194 (
            .O(N__7983),
            .I(\DUT.uart_inst0.tx_dataZ0Z_7 ));
    CascadeMux I__1193 (
            .O(N__7980),
            .I(N__7977));
    InMux I__1192 (
            .O(N__7977),
            .I(N__7974));
    LocalMux I__1191 (
            .O(N__7974),
            .I(\DUT.uart_inst0.tx_dataZ0Z_6 ));
    CEMux I__1190 (
            .O(N__7971),
            .I(N__7967));
    CEMux I__1189 (
            .O(N__7970),
            .I(N__7964));
    LocalMux I__1188 (
            .O(N__7967),
            .I(\DUT.uart_inst0.N_22_i ));
    LocalMux I__1187 (
            .O(N__7964),
            .I(\DUT.uart_inst0.N_22_i ));
    InMux I__1186 (
            .O(N__7959),
            .I(N__7950));
    InMux I__1185 (
            .O(N__7958),
            .I(N__7950));
    InMux I__1184 (
            .O(N__7957),
            .I(N__7950));
    LocalMux I__1183 (
            .O(N__7950),
            .I(\DUT.uart_inst0.N_102 ));
    InMux I__1182 (
            .O(N__7947),
            .I(N__7944));
    LocalMux I__1181 (
            .O(N__7944),
            .I(N__7941));
    Span4Mux_h I__1180 (
            .O(N__7941),
            .I(N__7938));
    Odrv4 I__1179 (
            .O(N__7938),
            .I(\DUT.uart_inst0.tx_state_0_sqmuxa_i_i_a3_0_1 ));
    CascadeMux I__1178 (
            .O(N__7935),
            .I(G_110_cascade_));
    InMux I__1177 (
            .O(N__7932),
            .I(N__7929));
    LocalMux I__1176 (
            .O(N__7929),
            .I(fifo_inst_ftdi_input_inst_oTxFull_0));
    InMux I__1175 (
            .O(N__7926),
            .I(N__7918));
    InMux I__1174 (
            .O(N__7925),
            .I(N__7918));
    InMux I__1173 (
            .O(N__7924),
            .I(N__7913));
    InMux I__1172 (
            .O(N__7923),
            .I(N__7913));
    LocalMux I__1171 (
            .O(N__7918),
            .I(G_108));
    LocalMux I__1170 (
            .O(N__7913),
            .I(G_108));
    InMux I__1169 (
            .O(N__7908),
            .I(N__7905));
    LocalMux I__1168 (
            .O(N__7905),
            .I(\fifo_inst.ftdi_input_inst.SUMZ0Z_3 ));
    InMux I__1167 (
            .O(N__7902),
            .I(N__7893));
    InMux I__1166 (
            .O(N__7901),
            .I(N__7893));
    InMux I__1165 (
            .O(N__7900),
            .I(N__7886));
    InMux I__1164 (
            .O(N__7899),
            .I(N__7886));
    InMux I__1163 (
            .O(N__7898),
            .I(N__7886));
    LocalMux I__1162 (
            .O(N__7893),
            .I(G_109));
    LocalMux I__1161 (
            .O(N__7886),
            .I(G_109));
    CascadeMux I__1160 (
            .O(N__7881),
            .I(N__7875));
    CascadeMux I__1159 (
            .O(N__7880),
            .I(N__7872));
    CascadeMux I__1158 (
            .O(N__7879),
            .I(N__7869));
    InMux I__1157 (
            .O(N__7878),
            .I(N__7863));
    InMux I__1156 (
            .O(N__7875),
            .I(N__7863));
    InMux I__1155 (
            .O(N__7872),
            .I(N__7856));
    InMux I__1154 (
            .O(N__7869),
            .I(N__7856));
    InMux I__1153 (
            .O(N__7868),
            .I(N__7856));
    LocalMux I__1152 (
            .O(N__7863),
            .I(G_110));
    LocalMux I__1151 (
            .O(N__7856),
            .I(G_110));
    CascadeMux I__1150 (
            .O(N__7851),
            .I(N__7848));
    InMux I__1149 (
            .O(N__7848),
            .I(N__7840));
    InMux I__1148 (
            .O(N__7847),
            .I(N__7840));
    InMux I__1147 (
            .O(N__7846),
            .I(N__7835));
    InMux I__1146 (
            .O(N__7845),
            .I(N__7835));
    LocalMux I__1145 (
            .O(N__7840),
            .I(G_111));
    LocalMux I__1144 (
            .O(N__7835),
            .I(G_111));
    InMux I__1143 (
            .O(N__7830),
            .I(N__7821));
    InMux I__1142 (
            .O(N__7829),
            .I(N__7821));
    InMux I__1141 (
            .O(N__7828),
            .I(N__7814));
    InMux I__1140 (
            .O(N__7827),
            .I(N__7814));
    InMux I__1139 (
            .O(N__7826),
            .I(N__7814));
    LocalMux I__1138 (
            .O(N__7821),
            .I(G_112));
    LocalMux I__1137 (
            .O(N__7814),
            .I(G_112));
    InMux I__1136 (
            .O(N__7809),
            .I(N__7806));
    LocalMux I__1135 (
            .O(N__7806),
            .I(N__7803));
    Span4Mux_h I__1134 (
            .O(N__7803),
            .I(N__7800));
    Odrv4 I__1133 (
            .O(N__7800),
            .I(\fifo_inst.ftdi_input_inst.un2_oPacketAvail_iZ0 ));
    InMux I__1132 (
            .O(N__7797),
            .I(N__7794));
    LocalMux I__1131 (
            .O(N__7794),
            .I(N__7791));
    Span4Mux_h I__1130 (
            .O(N__7791),
            .I(N__7787));
    InMux I__1129 (
            .O(N__7790),
            .I(N__7784));
    Odrv4 I__1128 (
            .O(N__7787),
            .I(\DUT.uart_inst0.tx_dataZ0Z_0 ));
    LocalMux I__1127 (
            .O(N__7784),
            .I(\DUT.uart_inst0.tx_dataZ0Z_0 ));
    IoInMux I__1126 (
            .O(N__7779),
            .I(N__7775));
    CascadeMux I__1125 (
            .O(N__7778),
            .I(N__7772));
    LocalMux I__1124 (
            .O(N__7775),
            .I(N__7769));
    InMux I__1123 (
            .O(N__7772),
            .I(N__7765));
    Span4Mux_s3_v I__1122 (
            .O(N__7769),
            .I(N__7762));
    InMux I__1121 (
            .O(N__7768),
            .I(N__7759));
    LocalMux I__1120 (
            .O(N__7765),
            .I(N__7755));
    Span4Mux_h I__1119 (
            .O(N__7762),
            .I(N__7752));
    LocalMux I__1118 (
            .O(N__7759),
            .I(N__7749));
    InMux I__1117 (
            .O(N__7758),
            .I(N__7746));
    Span4Mux_v I__1116 (
            .O(N__7755),
            .I(N__7743));
    Odrv4 I__1115 (
            .O(N__7752),
            .I(P1A7_c));
    Odrv4 I__1114 (
            .O(N__7749),
            .I(P1A7_c));
    LocalMux I__1113 (
            .O(N__7746),
            .I(P1A7_c));
    Odrv4 I__1112 (
            .O(N__7743),
            .I(P1A7_c));
    InMux I__1111 (
            .O(N__7734),
            .I(N__7731));
    LocalMux I__1110 (
            .O(N__7731),
            .I(N__7728));
    Odrv12 I__1109 (
            .O(N__7728),
            .I(\DUT.uart_inst0.N_116 ));
    CascadeMux I__1108 (
            .O(N__7725),
            .I(\DUT.uart_inst0.m13_2_cascade_ ));
    InMux I__1107 (
            .O(N__7722),
            .I(N__7719));
    LocalMux I__1106 (
            .O(N__7719),
            .I(\DUT.uart_inst0.m13_3 ));
    CascadeMux I__1105 (
            .O(N__7716),
            .I(\DUT.uart_inst0.P19_mux_cascade_ ));
    InMux I__1104 (
            .O(N__7713),
            .I(N__7710));
    LocalMux I__1103 (
            .O(N__7710),
            .I(N__7707));
    Odrv4 I__1102 (
            .O(N__7707),
            .I(\DUT.uart_inst0.g0_0_1 ));
    IoInMux I__1101 (
            .O(N__7704),
            .I(N__7701));
    LocalMux I__1100 (
            .O(N__7701),
            .I(N__7698));
    Span4Mux_s1_v I__1099 (
            .O(N__7698),
            .I(N__7695));
    Odrv4 I__1098 (
            .O(N__7695),
            .I(N_1257_i));
    CascadeMux I__1097 (
            .O(N__7692),
            .I(G_111_cascade_));
    CascadeMux I__1096 (
            .O(N__7689),
            .I(\fifo_inst.ftdi_input_inst.SUMZ0Z_2_cascade_ ));
    InMux I__1095 (
            .O(N__7686),
            .I(N__7683));
    LocalMux I__1094 (
            .O(N__7683),
            .I(\DUT.uart_inst0.g0_0_0_a3_0_4 ));
    CascadeMux I__1093 (
            .O(N__7680),
            .I(\DUT.uart_inst0.g0_0_0_a3_4_cascade_ ));
    InMux I__1092 (
            .O(N__7677),
            .I(N__7674));
    LocalMux I__1091 (
            .O(N__7674),
            .I(\DUT.uart_inst0.g0_0_0_a3_3 ));
    CascadeMux I__1090 (
            .O(N__7671),
            .I(\DUT.fifo_tx_inst.un1_i11_i_cascade_ ));
    CascadeMux I__1089 (
            .O(N__7668),
            .I(\DUT.fifo_rx_inst.N_57_cascade_ ));
    InMux I__1088 (
            .O(N__7665),
            .I(N__7659));
    InMux I__1087 (
            .O(N__7664),
            .I(N__7659));
    LocalMux I__1086 (
            .O(N__7659),
            .I(\DUT.fifo_rx_inst.un1_i11_i ));
    CascadeMux I__1085 (
            .O(N__7656),
            .I(\DUT.uart_inst0.N_21_0_cascade_ ));
    InMux I__1084 (
            .O(N__7653),
            .I(N__7650));
    LocalMux I__1083 (
            .O(N__7650),
            .I(\DUT.uart_inst0.N_21_mux_0 ));
    InMux I__1082 (
            .O(N__7647),
            .I(N__7644));
    LocalMux I__1081 (
            .O(N__7644),
            .I(\DUT.uart_inst0.m5_1 ));
    InMux I__1080 (
            .O(N__7641),
            .I(N__7638));
    LocalMux I__1079 (
            .O(N__7638),
            .I(\DUT.uart_inst0.N_6 ));
    CascadeMux I__1078 (
            .O(N__7635),
            .I(\DUT.uart_inst0.N_6_cascade_ ));
    InMux I__1077 (
            .O(N__7632),
            .I(N__7629));
    LocalMux I__1076 (
            .O(N__7629),
            .I(N__7626));
    Odrv4 I__1075 (
            .O(N__7626),
            .I(\DUT.uart_inst0.N_18 ));
    InMux I__1074 (
            .O(N__7623),
            .I(N__7620));
    LocalMux I__1073 (
            .O(N__7620),
            .I(\DUT.uart_inst0.N_18_mux_0 ));
    InMux I__1072 (
            .O(N__7617),
            .I(N__7614));
    LocalMux I__1071 (
            .O(N__7614),
            .I(N__7611));
    Span4Mux_h I__1070 (
            .O(N__7611),
            .I(N__7608));
    Odrv4 I__1069 (
            .O(N__7608),
            .I(\DUT.uart_inst0.N_30 ));
    CascadeMux I__1068 (
            .O(N__7605),
            .I(N__7602));
    InMux I__1067 (
            .O(N__7602),
            .I(N__7599));
    LocalMux I__1066 (
            .O(N__7599),
            .I(N__7596));
    Odrv4 I__1065 (
            .O(N__7596),
            .I(\DUT.uart_inst0.g1_i_a4_0_4 ));
    CascadeMux I__1064 (
            .O(N__7593),
            .I(\DUT.uart_inst0.g1_i_a4_0_5_cascade_ ));
    CascadeMux I__1063 (
            .O(N__7590),
            .I(\DUT.uart_inst0.m7_e_1_cascade_ ));
    CascadeMux I__1062 (
            .O(N__7587),
            .I(\DUT.uart_inst0.m7_e_3_cascade_ ));
    CascadeMux I__1061 (
            .O(N__7584),
            .I(\DUT.uart_inst0.m9_1_cascade_ ));
    InMux I__1060 (
            .O(N__7581),
            .I(N__7578));
    LocalMux I__1059 (
            .O(N__7578),
            .I(\DUT.uart_inst0.N_11_mux ));
    InMux I__1058 (
            .O(N__7575),
            .I(N__7572));
    LocalMux I__1057 (
            .O(N__7572),
            .I(\DUT.uart_inst0.N_66 ));
    CascadeMux I__1056 (
            .O(N__7569),
            .I(N__7566));
    InMux I__1055 (
            .O(N__7566),
            .I(N__7563));
    LocalMux I__1054 (
            .O(N__7563),
            .I(N__7560));
    Span4Mux_h I__1053 (
            .O(N__7560),
            .I(N__7557));
    Odrv4 I__1052 (
            .O(N__7557),
            .I(\DUT.uart_inst0.m4_e_0 ));
    InMux I__1051 (
            .O(N__7554),
            .I(N__7551));
    LocalMux I__1050 (
            .O(N__7551),
            .I(\DUT.uart_inst0.m4_e_3 ));
    CascadeMux I__1049 (
            .O(N__7548),
            .I(N__7545));
    InMux I__1048 (
            .O(N__7545),
            .I(N__7542));
    LocalMux I__1047 (
            .O(N__7542),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO ));
    InMux I__1046 (
            .O(N__7539),
            .I(N__7534));
    InMux I__1045 (
            .O(N__7538),
            .I(N__7531));
    InMux I__1044 (
            .O(N__7537),
            .I(N__7528));
    LocalMux I__1043 (
            .O(N__7534),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_11 ));
    LocalMux I__1042 (
            .O(N__7531),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_11 ));
    LocalMux I__1041 (
            .O(N__7528),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_11 ));
    InMux I__1040 (
            .O(N__7521),
            .I(N__7518));
    LocalMux I__1039 (
            .O(N__7518),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO ));
    CascadeMux I__1038 (
            .O(N__7515),
            .I(N__7512));
    InMux I__1037 (
            .O(N__7512),
            .I(N__7507));
    InMux I__1036 (
            .O(N__7511),
            .I(N__7504));
    InMux I__1035 (
            .O(N__7510),
            .I(N__7501));
    LocalMux I__1034 (
            .O(N__7507),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_7 ));
    LocalMux I__1033 (
            .O(N__7504),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_7 ));
    LocalMux I__1032 (
            .O(N__7501),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_7 ));
    InMux I__1031 (
            .O(N__7494),
            .I(N__7491));
    LocalMux I__1030 (
            .O(N__7491),
            .I(\DUT.uart_inst0.rx_clk_divider_1_5 ));
    InMux I__1029 (
            .O(N__7488),
            .I(N__7484));
    InMux I__1028 (
            .O(N__7487),
            .I(N__7481));
    LocalMux I__1027 (
            .O(N__7484),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_5 ));
    LocalMux I__1026 (
            .O(N__7481),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_5 ));
    InMux I__1025 (
            .O(N__7476),
            .I(N__7473));
    LocalMux I__1024 (
            .O(N__7473),
            .I(\DUT.uart_inst0.rx_clk_divider_1_6 ));
    InMux I__1023 (
            .O(N__7470),
            .I(N__7466));
    InMux I__1022 (
            .O(N__7469),
            .I(N__7463));
    LocalMux I__1021 (
            .O(N__7466),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_6 ));
    LocalMux I__1020 (
            .O(N__7463),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_6 ));
    InMux I__1019 (
            .O(N__7458),
            .I(N__7455));
    LocalMux I__1018 (
            .O(N__7455),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO ));
    CascadeMux I__1017 (
            .O(N__7452),
            .I(N__7447));
    InMux I__1016 (
            .O(N__7451),
            .I(N__7444));
    InMux I__1015 (
            .O(N__7450),
            .I(N__7439));
    InMux I__1014 (
            .O(N__7447),
            .I(N__7439));
    LocalMux I__1013 (
            .O(N__7444),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_8 ));
    LocalMux I__1012 (
            .O(N__7439),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_8 ));
    InMux I__1011 (
            .O(N__7434),
            .I(N__7431));
    LocalMux I__1010 (
            .O(N__7431),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO ));
    CascadeMux I__1009 (
            .O(N__7428),
            .I(N__7423));
    InMux I__1008 (
            .O(N__7427),
            .I(N__7420));
    InMux I__1007 (
            .O(N__7426),
            .I(N__7417));
    InMux I__1006 (
            .O(N__7423),
            .I(N__7414));
    LocalMux I__1005 (
            .O(N__7420),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_12 ));
    LocalMux I__1004 (
            .O(N__7417),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_12 ));
    LocalMux I__1003 (
            .O(N__7414),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_12 ));
    InMux I__1002 (
            .O(N__7407),
            .I(N__7404));
    LocalMux I__1001 (
            .O(N__7404),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO ));
    CascadeMux I__1000 (
            .O(N__7401),
            .I(N__7398));
    InMux I__999 (
            .O(N__7398),
            .I(N__7394));
    InMux I__998 (
            .O(N__7397),
            .I(N__7391));
    LocalMux I__997 (
            .O(N__7394),
            .I(\DUT.uart_inst0.tx_countdown_30_5 ));
    LocalMux I__996 (
            .O(N__7391),
            .I(\DUT.uart_inst0.tx_countdown_30_5 ));
    InMux I__995 (
            .O(N__7386),
            .I(N__7383));
    LocalMux I__994 (
            .O(N__7383),
            .I(N__7380));
    Odrv4 I__993 (
            .O(N__7380),
            .I(\DUT.uart_inst0.tx_countdown_7_m1_0_a3_0_2 ));
    CascadeMux I__992 (
            .O(N__7377),
            .I(N__7374));
    InMux I__991 (
            .O(N__7374),
            .I(N__7371));
    LocalMux I__990 (
            .O(N__7371),
            .I(\DUT.uart_inst0.N_113 ));
    InMux I__989 (
            .O(N__7368),
            .I(N__7358));
    InMux I__988 (
            .O(N__7367),
            .I(N__7358));
    InMux I__987 (
            .O(N__7366),
            .I(N__7351));
    InMux I__986 (
            .O(N__7365),
            .I(N__7351));
    InMux I__985 (
            .O(N__7364),
            .I(N__7351));
    InMux I__984 (
            .O(N__7363),
            .I(N__7348));
    LocalMux I__983 (
            .O(N__7358),
            .I(N__7345));
    LocalMux I__982 (
            .O(N__7351),
            .I(N__7342));
    LocalMux I__981 (
            .O(N__7348),
            .I(\DUT.uart_inst0.tx_countdown_7_sm0_0 ));
    Odrv4 I__980 (
            .O(N__7345),
            .I(\DUT.uart_inst0.tx_countdown_7_sm0_0 ));
    Odrv4 I__979 (
            .O(N__7342),
            .I(\DUT.uart_inst0.tx_countdown_7_sm0_0 ));
    CascadeMux I__978 (
            .O(N__7335),
            .I(N__7332));
    InMux I__977 (
            .O(N__7332),
            .I(N__7328));
    CascadeMux I__976 (
            .O(N__7331),
            .I(N__7325));
    LocalMux I__975 (
            .O(N__7328),
            .I(N__7322));
    InMux I__974 (
            .O(N__7325),
            .I(N__7314));
    Span4Mux_s2_v I__973 (
            .O(N__7322),
            .I(N__7311));
    InMux I__972 (
            .O(N__7321),
            .I(N__7308));
    InMux I__971 (
            .O(N__7320),
            .I(N__7303));
    InMux I__970 (
            .O(N__7319),
            .I(N__7303));
    InMux I__969 (
            .O(N__7318),
            .I(N__7298));
    InMux I__968 (
            .O(N__7317),
            .I(N__7298));
    LocalMux I__967 (
            .O(N__7314),
            .I(\DUT.uart_inst0.N_84 ));
    Odrv4 I__966 (
            .O(N__7311),
            .I(\DUT.uart_inst0.N_84 ));
    LocalMux I__965 (
            .O(N__7308),
            .I(\DUT.uart_inst0.N_84 ));
    LocalMux I__964 (
            .O(N__7303),
            .I(\DUT.uart_inst0.N_84 ));
    LocalMux I__963 (
            .O(N__7298),
            .I(\DUT.uart_inst0.N_84 ));
    CascadeMux I__962 (
            .O(N__7287),
            .I(N__7283));
    CascadeMux I__961 (
            .O(N__7286),
            .I(N__7280));
    InMux I__960 (
            .O(N__7283),
            .I(N__7277));
    InMux I__959 (
            .O(N__7280),
            .I(N__7274));
    LocalMux I__958 (
            .O(N__7277),
            .I(N__7271));
    LocalMux I__957 (
            .O(N__7274),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_17 ));
    Odrv4 I__956 (
            .O(N__7271),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_17 ));
    InMux I__955 (
            .O(N__7266),
            .I(N__7263));
    LocalMux I__954 (
            .O(N__7263),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO ));
    InMux I__953 (
            .O(N__7260),
            .I(N__7255));
    InMux I__952 (
            .O(N__7259),
            .I(N__7252));
    InMux I__951 (
            .O(N__7258),
            .I(N__7249));
    LocalMux I__950 (
            .O(N__7255),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_13 ));
    LocalMux I__949 (
            .O(N__7252),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_13 ));
    LocalMux I__948 (
            .O(N__7249),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_13 ));
    InMux I__947 (
            .O(N__7242),
            .I(N__7239));
    LocalMux I__946 (
            .O(N__7239),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO ));
    CascadeMux I__945 (
            .O(N__7236),
            .I(N__7233));
    InMux I__944 (
            .O(N__7233),
            .I(N__7228));
    InMux I__943 (
            .O(N__7232),
            .I(N__7225));
    InMux I__942 (
            .O(N__7231),
            .I(N__7222));
    LocalMux I__941 (
            .O(N__7228),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_14 ));
    LocalMux I__940 (
            .O(N__7225),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_14 ));
    LocalMux I__939 (
            .O(N__7222),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_14 ));
    InMux I__938 (
            .O(N__7215),
            .I(N__7212));
    LocalMux I__937 (
            .O(N__7212),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO ));
    InMux I__936 (
            .O(N__7209),
            .I(N__7204));
    InMux I__935 (
            .O(N__7208),
            .I(N__7199));
    InMux I__934 (
            .O(N__7207),
            .I(N__7199));
    LocalMux I__933 (
            .O(N__7204),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_15 ));
    LocalMux I__932 (
            .O(N__7199),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_15 ));
    CascadeMux I__931 (
            .O(N__7194),
            .I(N__7191));
    InMux I__930 (
            .O(N__7191),
            .I(N__7188));
    LocalMux I__929 (
            .O(N__7188),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO ));
    InMux I__928 (
            .O(N__7185),
            .I(N__7180));
    InMux I__927 (
            .O(N__7184),
            .I(N__7175));
    InMux I__926 (
            .O(N__7183),
            .I(N__7175));
    LocalMux I__925 (
            .O(N__7180),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_10 ));
    LocalMux I__924 (
            .O(N__7175),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_10 ));
    CascadeMux I__923 (
            .O(N__7170),
            .I(N__7167));
    InMux I__922 (
            .O(N__7167),
            .I(N__7164));
    LocalMux I__921 (
            .O(N__7164),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO ));
    InMux I__920 (
            .O(N__7161),
            .I(N__7156));
    InMux I__919 (
            .O(N__7160),
            .I(N__7151));
    InMux I__918 (
            .O(N__7159),
            .I(N__7151));
    LocalMux I__917 (
            .O(N__7156),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_9 ));
    LocalMux I__916 (
            .O(N__7151),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_9 ));
    CascadeMux I__915 (
            .O(N__7146),
            .I(\DUT.uart_inst0.N_218_cascade_ ));
    InMux I__914 (
            .O(N__7143),
            .I(N__7138));
    InMux I__913 (
            .O(N__7142),
            .I(N__7133));
    InMux I__912 (
            .O(N__7141),
            .I(N__7133));
    LocalMux I__911 (
            .O(N__7138),
            .I(\DUT.uart_inst0.N_109 ));
    LocalMux I__910 (
            .O(N__7133),
            .I(\DUT.uart_inst0.N_109 ));
    InMux I__909 (
            .O(N__7128),
            .I(N__7115));
    InMux I__908 (
            .O(N__7127),
            .I(N__7115));
    InMux I__907 (
            .O(N__7126),
            .I(N__7110));
    InMux I__906 (
            .O(N__7125),
            .I(N__7110));
    InMux I__905 (
            .O(N__7124),
            .I(N__7105));
    InMux I__904 (
            .O(N__7123),
            .I(N__7105));
    InMux I__903 (
            .O(N__7122),
            .I(N__7098));
    InMux I__902 (
            .O(N__7121),
            .I(N__7098));
    InMux I__901 (
            .O(N__7120),
            .I(N__7098));
    LocalMux I__900 (
            .O(N__7115),
            .I(N__7095));
    LocalMux I__899 (
            .O(N__7110),
            .I(N__7088));
    LocalMux I__898 (
            .O(N__7105),
            .I(N__7088));
    LocalMux I__897 (
            .O(N__7098),
            .I(N__7088));
    Odrv4 I__896 (
            .O(N__7095),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_1 ));
    Odrv4 I__895 (
            .O(N__7088),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_1 ));
    CascadeMux I__894 (
            .O(N__7083),
            .I(N__7077));
    InMux I__893 (
            .O(N__7082),
            .I(N__7073));
    CascadeMux I__892 (
            .O(N__7081),
            .I(N__7066));
    InMux I__891 (
            .O(N__7080),
            .I(N__7061));
    InMux I__890 (
            .O(N__7077),
            .I(N__7061));
    InMux I__889 (
            .O(N__7076),
            .I(N__7058));
    LocalMux I__888 (
            .O(N__7073),
            .I(N__7055));
    InMux I__887 (
            .O(N__7072),
            .I(N__7048));
    InMux I__886 (
            .O(N__7071),
            .I(N__7048));
    InMux I__885 (
            .O(N__7070),
            .I(N__7048));
    InMux I__884 (
            .O(N__7069),
            .I(N__7043));
    InMux I__883 (
            .O(N__7066),
            .I(N__7043));
    LocalMux I__882 (
            .O(N__7061),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_0 ));
    LocalMux I__881 (
            .O(N__7058),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_0 ));
    Odrv4 I__880 (
            .O(N__7055),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_0 ));
    LocalMux I__879 (
            .O(N__7048),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_0 ));
    LocalMux I__878 (
            .O(N__7043),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_0 ));
    InMux I__877 (
            .O(N__7032),
            .I(N__7029));
    LocalMux I__876 (
            .O(N__7029),
            .I(N__7025));
    InMux I__875 (
            .O(N__7028),
            .I(N__7022));
    Odrv4 I__874 (
            .O(N__7025),
            .I(\DUT.uart_inst0.N_120 ));
    LocalMux I__873 (
            .O(N__7022),
            .I(\DUT.uart_inst0.N_120 ));
    CascadeMux I__872 (
            .O(N__7017),
            .I(\DUT.uart_inst0.tx_countdown_RNO_1Z0Z_3_cascade_ ));
    InMux I__871 (
            .O(N__7014),
            .I(N__7005));
    InMux I__870 (
            .O(N__7013),
            .I(N__7002));
    InMux I__869 (
            .O(N__7012),
            .I(N__6989));
    InMux I__868 (
            .O(N__7011),
            .I(N__6989));
    InMux I__867 (
            .O(N__7010),
            .I(N__6989));
    InMux I__866 (
            .O(N__7009),
            .I(N__6989));
    InMux I__865 (
            .O(N__7008),
            .I(N__6986));
    LocalMux I__864 (
            .O(N__7005),
            .I(N__6983));
    LocalMux I__863 (
            .O(N__7002),
            .I(N__6980));
    InMux I__862 (
            .O(N__7001),
            .I(N__6971));
    InMux I__861 (
            .O(N__7000),
            .I(N__6971));
    InMux I__860 (
            .O(N__6999),
            .I(N__6971));
    InMux I__859 (
            .O(N__6998),
            .I(N__6971));
    LocalMux I__858 (
            .O(N__6989),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0 ));
    LocalMux I__857 (
            .O(N__6986),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0 ));
    Odrv4 I__856 (
            .O(N__6983),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0 ));
    Odrv4 I__855 (
            .O(N__6980),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0 ));
    LocalMux I__854 (
            .O(N__6971),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0 ));
    InMux I__853 (
            .O(N__6960),
            .I(N__6951));
    InMux I__852 (
            .O(N__6959),
            .I(N__6951));
    InMux I__851 (
            .O(N__6958),
            .I(N__6951));
    LocalMux I__850 (
            .O(N__6951),
            .I(\DUT.uart_inst0.N_164 ));
    CascadeMux I__849 (
            .O(N__6948),
            .I(\DUT.uart_inst0.N_164_cascade_ ));
    InMux I__848 (
            .O(N__6945),
            .I(N__6942));
    LocalMux I__847 (
            .O(N__6942),
            .I(\DUT.uart_inst0.tx_countdown_RNO_0Z0Z_3 ));
    CascadeMux I__846 (
            .O(N__6939),
            .I(N__6935));
    InMux I__845 (
            .O(N__6938),
            .I(N__6928));
    InMux I__844 (
            .O(N__6935),
            .I(N__6928));
    InMux I__843 (
            .O(N__6934),
            .I(N__6923));
    InMux I__842 (
            .O(N__6933),
            .I(N__6923));
    LocalMux I__841 (
            .O(N__6928),
            .I(N__6918));
    LocalMux I__840 (
            .O(N__6923),
            .I(N__6918));
    Odrv4 I__839 (
            .O(N__6918),
            .I(\DUT.uart_inst0.tx_state_ns_i_i_o2_a0_2_0 ));
    InMux I__838 (
            .O(N__6915),
            .I(N__6912));
    LocalMux I__837 (
            .O(N__6912),
            .I(N__6905));
    InMux I__836 (
            .O(N__6911),
            .I(N__6900));
    InMux I__835 (
            .O(N__6910),
            .I(N__6900));
    InMux I__834 (
            .O(N__6909),
            .I(N__6895));
    InMux I__833 (
            .O(N__6908),
            .I(N__6895));
    Span4Mux_v I__832 (
            .O(N__6905),
            .I(N__6888));
    LocalMux I__831 (
            .O(N__6900),
            .I(N__6888));
    LocalMux I__830 (
            .O(N__6895),
            .I(N__6888));
    Odrv4 I__829 (
            .O(N__6888),
            .I(\DUT.uart_inst0.N_159 ));
    InMux I__828 (
            .O(N__6885),
            .I(N__6882));
    LocalMux I__827 (
            .O(N__6882),
            .I(N__6875));
    InMux I__826 (
            .O(N__6881),
            .I(N__6870));
    InMux I__825 (
            .O(N__6880),
            .I(N__6870));
    InMux I__824 (
            .O(N__6879),
            .I(N__6867));
    InMux I__823 (
            .O(N__6878),
            .I(N__6864));
    Span4Mux_s1_v I__822 (
            .O(N__6875),
            .I(N__6859));
    LocalMux I__821 (
            .O(N__6870),
            .I(N__6859));
    LocalMux I__820 (
            .O(N__6867),
            .I(\DUT.uart_inst0.N_100 ));
    LocalMux I__819 (
            .O(N__6864),
            .I(\DUT.uart_inst0.N_100 ));
    Odrv4 I__818 (
            .O(N__6859),
            .I(\DUT.uart_inst0.N_100 ));
    InMux I__817 (
            .O(N__6852),
            .I(N__6849));
    LocalMux I__816 (
            .O(N__6849),
            .I(\DUT.uart_inst0.N_163 ));
    InMux I__815 (
            .O(N__6846),
            .I(N__6843));
    LocalMux I__814 (
            .O(N__6843),
            .I(N__6839));
    InMux I__813 (
            .O(N__6842),
            .I(N__6832));
    Span4Mux_s2_v I__812 (
            .O(N__6839),
            .I(N__6829));
    InMux I__811 (
            .O(N__6838),
            .I(N__6824));
    InMux I__810 (
            .O(N__6837),
            .I(N__6824));
    InMux I__809 (
            .O(N__6836),
            .I(N__6819));
    InMux I__808 (
            .O(N__6835),
            .I(N__6819));
    LocalMux I__807 (
            .O(N__6832),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_5 ));
    Odrv4 I__806 (
            .O(N__6829),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_5 ));
    LocalMux I__805 (
            .O(N__6824),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_5 ));
    LocalMux I__804 (
            .O(N__6819),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_5 ));
    CascadeMux I__803 (
            .O(N__6810),
            .I(N__6807));
    InMux I__802 (
            .O(N__6807),
            .I(N__6802));
    InMux I__801 (
            .O(N__6806),
            .I(N__6797));
    InMux I__800 (
            .O(N__6805),
            .I(N__6797));
    LocalMux I__799 (
            .O(N__6802),
            .I(\DUT.uart_inst0.tx_countdown_0_c3 ));
    LocalMux I__798 (
            .O(N__6797),
            .I(\DUT.uart_inst0.tx_countdown_0_c3 ));
    InMux I__797 (
            .O(N__6792),
            .I(N__6785));
    CascadeMux I__796 (
            .O(N__6791),
            .I(N__6781));
    CascadeMux I__795 (
            .O(N__6790),
            .I(N__6775));
    CascadeMux I__794 (
            .O(N__6789),
            .I(N__6772));
    InMux I__793 (
            .O(N__6788),
            .I(N__6769));
    LocalMux I__792 (
            .O(N__6785),
            .I(N__6766));
    InMux I__791 (
            .O(N__6784),
            .I(N__6759));
    InMux I__790 (
            .O(N__6781),
            .I(N__6759));
    InMux I__789 (
            .O(N__6780),
            .I(N__6759));
    InMux I__788 (
            .O(N__6779),
            .I(N__6750));
    InMux I__787 (
            .O(N__6778),
            .I(N__6750));
    InMux I__786 (
            .O(N__6775),
            .I(N__6750));
    InMux I__785 (
            .O(N__6772),
            .I(N__6750));
    LocalMux I__784 (
            .O(N__6769),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_3 ));
    Odrv4 I__783 (
            .O(N__6766),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_3 ));
    LocalMux I__782 (
            .O(N__6759),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_3 ));
    LocalMux I__781 (
            .O(N__6750),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_3 ));
    CascadeMux I__780 (
            .O(N__6741),
            .I(N__6737));
    InMux I__779 (
            .O(N__6740),
            .I(N__6734));
    InMux I__778 (
            .O(N__6737),
            .I(N__6725));
    LocalMux I__777 (
            .O(N__6734),
            .I(N__6722));
    InMux I__776 (
            .O(N__6733),
            .I(N__6713));
    InMux I__775 (
            .O(N__6732),
            .I(N__6713));
    InMux I__774 (
            .O(N__6731),
            .I(N__6713));
    InMux I__773 (
            .O(N__6730),
            .I(N__6713));
    InMux I__772 (
            .O(N__6729),
            .I(N__6708));
    InMux I__771 (
            .O(N__6728),
            .I(N__6708));
    LocalMux I__770 (
            .O(N__6725),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_4 ));
    Odrv4 I__769 (
            .O(N__6722),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_4 ));
    LocalMux I__768 (
            .O(N__6713),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_4 ));
    LocalMux I__767 (
            .O(N__6708),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_4 ));
    CascadeMux I__766 (
            .O(N__6699),
            .I(\DUT.uart_inst0.N_160_cascade_ ));
    InMux I__765 (
            .O(N__6696),
            .I(N__6688));
    InMux I__764 (
            .O(N__6695),
            .I(N__6688));
    InMux I__763 (
            .O(N__6694),
            .I(N__6683));
    InMux I__762 (
            .O(N__6693),
            .I(N__6683));
    LocalMux I__761 (
            .O(N__6688),
            .I(\DUT.uart_inst0.tx_countdown_0_ac0_1 ));
    LocalMux I__760 (
            .O(N__6683),
            .I(\DUT.uart_inst0.tx_countdown_0_ac0_1 ));
    InMux I__759 (
            .O(N__6678),
            .I(N__6675));
    LocalMux I__758 (
            .O(N__6675),
            .I(\DUT.uart_inst0.N_154 ));
    CascadeMux I__757 (
            .O(N__6672),
            .I(N__6666));
    InMux I__756 (
            .O(N__6671),
            .I(N__6662));
    InMux I__755 (
            .O(N__6670),
            .I(N__6657));
    InMux I__754 (
            .O(N__6669),
            .I(N__6657));
    InMux I__753 (
            .O(N__6666),
            .I(N__6654));
    InMux I__752 (
            .O(N__6665),
            .I(N__6651));
    LocalMux I__751 (
            .O(N__6662),
            .I(N__6648));
    LocalMux I__750 (
            .O(N__6657),
            .I(N__6645));
    LocalMux I__749 (
            .O(N__6654),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_3 ));
    LocalMux I__748 (
            .O(N__6651),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_3 ));
    Odrv4 I__747 (
            .O(N__6648),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_3 ));
    Odrv4 I__746 (
            .O(N__6645),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_3 ));
    InMux I__745 (
            .O(N__6636),
            .I(N__6633));
    LocalMux I__744 (
            .O(N__6633),
            .I(\DUT.uart_inst0.N_72 ));
    InMux I__743 (
            .O(N__6630),
            .I(N__6626));
    InMux I__742 (
            .O(N__6629),
            .I(N__6623));
    LocalMux I__741 (
            .O(N__6626),
            .I(\DUT.uart_inst0.N_99 ));
    LocalMux I__740 (
            .O(N__6623),
            .I(\DUT.uart_inst0.N_99 ));
    InMux I__739 (
            .O(N__6618),
            .I(N__6615));
    LocalMux I__738 (
            .O(N__6615),
            .I(N__6612));
    Span4Mux_s3_v I__737 (
            .O(N__6612),
            .I(N__6609));
    Odrv4 I__736 (
            .O(N__6609),
            .I(\DUT.uart_inst0.tx_countdown_RNO_0Z0Z_1 ));
    SRMux I__735 (
            .O(N__6606),
            .I(N__6602));
    SRMux I__734 (
            .O(N__6605),
            .I(N__6599));
    LocalMux I__733 (
            .O(N__6602),
            .I(N__6594));
    LocalMux I__732 (
            .O(N__6599),
            .I(N__6594));
    Span4Mux_v I__731 (
            .O(N__6594),
            .I(N__6591));
    Span4Mux_h I__730 (
            .O(N__6591),
            .I(N__6588));
    Odrv4 I__729 (
            .O(N__6588),
            .I(\DUT.uart_inst0.N_88_i ));
    CascadeMux I__728 (
            .O(N__6585),
            .I(N__6581));
    InMux I__727 (
            .O(N__6584),
            .I(N__6577));
    InMux I__726 (
            .O(N__6581),
            .I(N__6574));
    InMux I__725 (
            .O(N__6580),
            .I(N__6571));
    LocalMux I__724 (
            .O(N__6577),
            .I(\DUT.uart_inst0.N_160 ));
    LocalMux I__723 (
            .O(N__6574),
            .I(\DUT.uart_inst0.N_160 ));
    LocalMux I__722 (
            .O(N__6571),
            .I(\DUT.uart_inst0.N_160 ));
    InMux I__721 (
            .O(N__6564),
            .I(N__6561));
    LocalMux I__720 (
            .O(N__6561),
            .I(\DUT.uart_inst0.N_218 ));
    InMux I__719 (
            .O(N__6558),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_8 ));
    InMux I__718 (
            .O(N__6555),
            .I(N__6551));
    InMux I__717 (
            .O(N__6554),
            .I(N__6548));
    LocalMux I__716 (
            .O(N__6551),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_10 ));
    LocalMux I__715 (
            .O(N__6548),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_10 ));
    InMux I__714 (
            .O(N__6543),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_9 ));
    CascadeMux I__713 (
            .O(N__6540),
            .I(N__6536));
    InMux I__712 (
            .O(N__6539),
            .I(N__6533));
    InMux I__711 (
            .O(N__6536),
            .I(N__6530));
    LocalMux I__710 (
            .O(N__6533),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_11 ));
    LocalMux I__709 (
            .O(N__6530),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_11 ));
    InMux I__708 (
            .O(N__6525),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_10 ));
    InMux I__707 (
            .O(N__6522),
            .I(N__6518));
    InMux I__706 (
            .O(N__6521),
            .I(N__6515));
    LocalMux I__705 (
            .O(N__6518),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_12 ));
    LocalMux I__704 (
            .O(N__6515),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_12 ));
    InMux I__703 (
            .O(N__6510),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_11 ));
    InMux I__702 (
            .O(N__6507),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_12 ));
    CascadeMux I__701 (
            .O(N__6504),
            .I(N__6500));
    InMux I__700 (
            .O(N__6503),
            .I(N__6497));
    InMux I__699 (
            .O(N__6500),
            .I(N__6494));
    LocalMux I__698 (
            .O(N__6497),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_13 ));
    LocalMux I__697 (
            .O(N__6494),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_13 ));
    InMux I__696 (
            .O(N__6489),
            .I(N__6486));
    LocalMux I__695 (
            .O(N__6486),
            .I(N__6480));
    InMux I__694 (
            .O(N__6485),
            .I(N__6473));
    InMux I__693 (
            .O(N__6484),
            .I(N__6473));
    InMux I__692 (
            .O(N__6483),
            .I(N__6473));
    Odrv4 I__691 (
            .O(N__6480),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_2 ));
    LocalMux I__690 (
            .O(N__6473),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_2 ));
    InMux I__689 (
            .O(N__6468),
            .I(N__6465));
    LocalMux I__688 (
            .O(N__6465),
            .I(N__6461));
    InMux I__687 (
            .O(N__6464),
            .I(N__6455));
    Span4Mux_v I__686 (
            .O(N__6461),
            .I(N__6452));
    InMux I__685 (
            .O(N__6460),
            .I(N__6445));
    InMux I__684 (
            .O(N__6459),
            .I(N__6445));
    InMux I__683 (
            .O(N__6458),
            .I(N__6445));
    LocalMux I__682 (
            .O(N__6455),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_1 ));
    Odrv4 I__681 (
            .O(N__6452),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_1 ));
    LocalMux I__680 (
            .O(N__6445),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_1 ));
    InMux I__679 (
            .O(N__6438),
            .I(N__6435));
    LocalMux I__678 (
            .O(N__6435),
            .I(N__6432));
    Odrv4 I__677 (
            .O(N__6432),
            .I(\DUT.uart_inst0.m9_e_0_3 ));
    InMux I__676 (
            .O(N__6429),
            .I(N__6423));
    CascadeMux I__675 (
            .O(N__6428),
            .I(N__6418));
    CascadeMux I__674 (
            .O(N__6427),
            .I(N__6415));
    InMux I__673 (
            .O(N__6426),
            .I(N__6412));
    LocalMux I__672 (
            .O(N__6423),
            .I(N__6409));
    InMux I__671 (
            .O(N__6422),
            .I(N__6400));
    InMux I__670 (
            .O(N__6421),
            .I(N__6400));
    InMux I__669 (
            .O(N__6418),
            .I(N__6400));
    InMux I__668 (
            .O(N__6415),
            .I(N__6400));
    LocalMux I__667 (
            .O(N__6412),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_0 ));
    Odrv4 I__666 (
            .O(N__6409),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_0 ));
    LocalMux I__665 (
            .O(N__6400),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_0 ));
    InMux I__664 (
            .O(N__6393),
            .I(N__6390));
    LocalMux I__663 (
            .O(N__6390),
            .I(\DUT.uart_inst0.m9_e_0_0 ));
    InMux I__662 (
            .O(N__6387),
            .I(N__6383));
    InMux I__661 (
            .O(N__6386),
            .I(N__6380));
    LocalMux I__660 (
            .O(N__6383),
            .I(\DUT.uart_inst0.N_152 ));
    LocalMux I__659 (
            .O(N__6380),
            .I(\DUT.uart_inst0.N_152 ));
    CascadeMux I__658 (
            .O(N__6375),
            .I(\DUT.uart_inst0.tx_state_0_sqmuxa_i_i_a3_c_cascade_ ));
    InMux I__657 (
            .O(N__6372),
            .I(N__6368));
    InMux I__656 (
            .O(N__6371),
            .I(N__6365));
    LocalMux I__655 (
            .O(N__6368),
            .I(N__6362));
    LocalMux I__654 (
            .O(N__6365),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_1 ));
    Odrv4 I__653 (
            .O(N__6362),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_1 ));
    InMux I__652 (
            .O(N__6357),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_0 ));
    CascadeMux I__651 (
            .O(N__6354),
            .I(N__6350));
    InMux I__650 (
            .O(N__6353),
            .I(N__6347));
    InMux I__649 (
            .O(N__6350),
            .I(N__6344));
    LocalMux I__648 (
            .O(N__6347),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_2 ));
    LocalMux I__647 (
            .O(N__6344),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_2 ));
    InMux I__646 (
            .O(N__6339),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_1 ));
    InMux I__645 (
            .O(N__6336),
            .I(N__6332));
    InMux I__644 (
            .O(N__6335),
            .I(N__6329));
    LocalMux I__643 (
            .O(N__6332),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_3 ));
    LocalMux I__642 (
            .O(N__6329),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_3 ));
    InMux I__641 (
            .O(N__6324),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_2 ));
    InMux I__640 (
            .O(N__6321),
            .I(N__6317));
    InMux I__639 (
            .O(N__6320),
            .I(N__6314));
    LocalMux I__638 (
            .O(N__6317),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_4 ));
    LocalMux I__637 (
            .O(N__6314),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_4 ));
    InMux I__636 (
            .O(N__6309),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_3 ));
    InMux I__635 (
            .O(N__6306),
            .I(N__6302));
    InMux I__634 (
            .O(N__6305),
            .I(N__6299));
    LocalMux I__633 (
            .O(N__6302),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_5 ));
    LocalMux I__632 (
            .O(N__6299),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_5 ));
    InMux I__631 (
            .O(N__6294),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_4 ));
    InMux I__630 (
            .O(N__6291),
            .I(N__6287));
    InMux I__629 (
            .O(N__6290),
            .I(N__6284));
    LocalMux I__628 (
            .O(N__6287),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_6 ));
    LocalMux I__627 (
            .O(N__6284),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_6 ));
    InMux I__626 (
            .O(N__6279),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_5 ));
    InMux I__625 (
            .O(N__6276),
            .I(N__6272));
    InMux I__624 (
            .O(N__6275),
            .I(N__6269));
    LocalMux I__623 (
            .O(N__6272),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_7 ));
    LocalMux I__622 (
            .O(N__6269),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_7 ));
    InMux I__621 (
            .O(N__6264),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_6 ));
    InMux I__620 (
            .O(N__6261),
            .I(N__6257));
    InMux I__619 (
            .O(N__6260),
            .I(N__6254));
    LocalMux I__618 (
            .O(N__6257),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_8 ));
    LocalMux I__617 (
            .O(N__6254),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_8 ));
    InMux I__616 (
            .O(N__6249),
            .I(bfn_14_3_0_));
    InMux I__615 (
            .O(N__6246),
            .I(N__6242));
    InMux I__614 (
            .O(N__6245),
            .I(N__6239));
    LocalMux I__613 (
            .O(N__6242),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_9 ));
    LocalMux I__612 (
            .O(N__6239),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_9 ));
    CascadeMux I__611 (
            .O(N__6234),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_1_2_cascade_ ));
    InMux I__610 (
            .O(N__6231),
            .I(N__6228));
    LocalMux I__609 (
            .O(N__6228),
            .I(\DUT.uart_inst0.N_67 ));
    CascadeMux I__608 (
            .O(N__6225),
            .I(\DUT.uart_inst0.g0_0_0_a3_0_3_cascade_ ));
    InMux I__607 (
            .O(N__6222),
            .I(N__6219));
    LocalMux I__606 (
            .O(N__6219),
            .I(\DUT.uart_inst0.N_159_0 ));
    InMux I__605 (
            .O(N__6216),
            .I(N__6213));
    LocalMux I__604 (
            .O(N__6213),
            .I(\DUT.uart_inst0.N_4 ));
    InMux I__603 (
            .O(N__6210),
            .I(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0 ));
    InMux I__602 (
            .O(N__6207),
            .I(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1 ));
    InMux I__601 (
            .O(N__6204),
            .I(N__6201));
    LocalMux I__600 (
            .O(N__6201),
            .I(\DUT.fifo_tx_inst.rFifoCount_RNISSQ21Z0Z_1 ));
    CascadeMux I__599 (
            .O(N__6198),
            .I(\DUT.fifo_tx_inst.N_108_cascade_ ));
    InMux I__598 (
            .O(N__6195),
            .I(N__6192));
    LocalMux I__597 (
            .O(N__6192),
            .I(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0 ));
    InMux I__596 (
            .O(N__6189),
            .I(N__6184));
    InMux I__595 (
            .O(N__6188),
            .I(N__6179));
    InMux I__594 (
            .O(N__6187),
            .I(N__6179));
    LocalMux I__593 (
            .O(N__6184),
            .I(\DUT.fifo_tx_inst.N_108 ));
    LocalMux I__592 (
            .O(N__6179),
            .I(\DUT.fifo_tx_inst.N_108 ));
    CascadeMux I__591 (
            .O(N__6174),
            .I(N__6170));
    CascadeMux I__590 (
            .O(N__6173),
            .I(N__6167));
    InMux I__589 (
            .O(N__6170),
            .I(N__6159));
    InMux I__588 (
            .O(N__6167),
            .I(N__6159));
    InMux I__587 (
            .O(N__6166),
            .I(N__6159));
    LocalMux I__586 (
            .O(N__6159),
            .I(rTxWriteZ0));
    CascadeMux I__585 (
            .O(N__6156),
            .I(\DUT.fifo_tx_inst.N_104_cascade_ ));
    InMux I__584 (
            .O(N__6153),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_9 ));
    InMux I__583 (
            .O(N__6150),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_10 ));
    InMux I__582 (
            .O(N__6147),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_11 ));
    InMux I__581 (
            .O(N__6144),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_12 ));
    InMux I__580 (
            .O(N__6141),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_13 ));
    InMux I__579 (
            .O(N__6138),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_14 ));
    InMux I__578 (
            .O(N__6135),
            .I(bfn_13_9_0_));
    InMux I__577 (
            .O(N__6132),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_16 ));
    InMux I__576 (
            .O(N__6129),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_0 ));
    InMux I__575 (
            .O(N__6126),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_1 ));
    InMux I__574 (
            .O(N__6123),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_2 ));
    InMux I__573 (
            .O(N__6120),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_3 ));
    InMux I__572 (
            .O(N__6117),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_4 ));
    InMux I__571 (
            .O(N__6114),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_5 ));
    InMux I__570 (
            .O(N__6111),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_6 ));
    InMux I__569 (
            .O(N__6108),
            .I(bfn_13_8_0_));
    InMux I__568 (
            .O(N__6105),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_8 ));
    CascadeMux I__567 (
            .O(N__6102),
            .I(\DUT.uart_inst0.tx_countdown_RNO_0Z0Z_4_cascade_ ));
    CascadeMux I__566 (
            .O(N__6099),
            .I(\DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0_cascade_ ));
    CascadeMux I__565 (
            .O(N__6096),
            .I(\DUT.uart_inst0.m25_e_3_cascade_ ));
    CascadeMux I__564 (
            .O(N__6093),
            .I(N__6090));
    InMux I__563 (
            .O(N__6090),
            .I(N__6087));
    LocalMux I__562 (
            .O(N__6087),
            .I(N__6084));
    Odrv4 I__561 (
            .O(N__6084),
            .I(\DUT.uart_inst0.m3_0 ));
    InMux I__560 (
            .O(N__6081),
            .I(N__6078));
    LocalMux I__559 (
            .O(N__6078),
            .I(\DUT.uart_inst0.N_5 ));
    CascadeMux I__558 (
            .O(N__6075),
            .I(\DUT.uart_inst0.tx_countdown_7_m1_0_o2_2_2_cascade_ ));
    CascadeMux I__557 (
            .O(N__6072),
            .I(\DUT.uart_inst0.tx_out_6_iv_0_a3_0_1_cascade_ ));
    CascadeMux I__556 (
            .O(N__6069),
            .I(\DUT.uart_inst0.tx_out_6_iv_0_1_cascade_ ));
    InMux I__555 (
            .O(N__6066),
            .I(N__6063));
    LocalMux I__554 (
            .O(N__6063),
            .I(\DUT.uart_inst0.N_119 ));
    CascadeMux I__553 (
            .O(N__6060),
            .I(\DUT.uart_inst0.g2_3_cascade_ ));
    InMux I__552 (
            .O(N__6057),
            .I(N__6054));
    LocalMux I__551 (
            .O(N__6054),
            .I(\DUT.uart_inst0.g2 ));
    InMux I__550 (
            .O(N__6051),
            .I(N__6048));
    LocalMux I__549 (
            .O(N__6048),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_9 ));
    InMux I__548 (
            .O(N__6045),
            .I(N__6042));
    LocalMux I__547 (
            .O(N__6042),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_8 ));
    CascadeMux I__546 (
            .O(N__6039),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_6_cascade_ ));
    InMux I__545 (
            .O(N__6036),
            .I(N__6033));
    LocalMux I__544 (
            .O(N__6033),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_7 ));
    CascadeMux I__543 (
            .O(N__6030),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0_cascade_ ));
    CascadeMux I__542 (
            .O(N__6027),
            .I(\DUT.uart_inst0.N_152_cascade_ ));
    CascadeMux I__541 (
            .O(N__6024),
            .I(\DUT.uart_inst0.N_6_0_cascade_ ));
    CascadeMux I__540 (
            .O(N__6021),
            .I(\DUT.uart_inst0.N_22_cascade_ ));
    CascadeMux I__539 (
            .O(N__6018),
            .I(N__6015));
    InMux I__538 (
            .O(N__6015),
            .I(N__6009));
    InMux I__537 (
            .O(N__6014),
            .I(N__6009));
    LocalMux I__536 (
            .O(N__6009),
            .I(\DUT.uart_inst0.N_22 ));
    IoInMux I__535 (
            .O(N__6006),
            .I(N__6003));
    LocalMux I__534 (
            .O(N__6003),
            .I(N__6000));
    IoSpan4Mux I__533 (
            .O(N__6000),
            .I(N__5997));
    Sp12to4 I__532 (
            .O(N__5997),
            .I(N__5994));
    Span12Mux_s7_v I__531 (
            .O(N__5994),
            .I(N__5991));
    Odrv12 I__530 (
            .O(N__5991),
            .I(wRamRdData_0));
    IoInMux I__529 (
            .O(N__5988),
            .I(N__5985));
    LocalMux I__528 (
            .O(N__5985),
            .I(N__5982));
    Span4Mux_s3_v I__527 (
            .O(N__5982),
            .I(N__5979));
    Span4Mux_v I__526 (
            .O(N__5979),
            .I(N__5976));
    Odrv4 I__525 (
            .O(N__5976),
            .I(wRamRdData_3));
    InMux I__524 (
            .O(N__5973),
            .I(N__5970));
    LocalMux I__523 (
            .O(N__5970),
            .I(\PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO ));
    IoInMux I__522 (
            .O(N__5967),
            .I(N__5964));
    LocalMux I__521 (
            .O(N__5964),
            .I(\top_pll_inst.wPllLocked_iso_i ));
    IoInMux I__520 (
            .O(N__5961),
            .I(N__5958));
    LocalMux I__519 (
            .O(N__5958),
            .I(N__5955));
    Span12Mux_s1_v I__518 (
            .O(N__5955),
            .I(N__5952));
    Odrv12 I__517 (
            .O(N__5952),
            .I(wRamRdData_4));
    IoInMux I__516 (
            .O(N__5949),
            .I(N__5946));
    LocalMux I__515 (
            .O(N__5946),
            .I(N__5943));
    Span12Mux_s9_v I__514 (
            .O(N__5943),
            .I(N__5940));
    Span12Mux_v I__513 (
            .O(N__5940),
            .I(N__5937));
    Odrv12 I__512 (
            .O(N__5937),
            .I(BTN_N_c));
    IoInMux I__511 (
            .O(N__5934),
            .I(N__5931));
    LocalMux I__510 (
            .O(N__5931),
            .I(N__5928));
    Span12Mux_s2_v I__509 (
            .O(N__5928),
            .I(N__5925));
    Span12Mux_v I__508 (
            .O(N__5925),
            .I(N__5922));
    Odrv12 I__507 (
            .O(N__5922),
            .I(wRamRdData_7));
    IoInMux I__506 (
            .O(N__5919),
            .I(N__5916));
    LocalMux I__505 (
            .O(N__5916),
            .I(N__5913));
    IoSpan4Mux I__504 (
            .O(N__5913),
            .I(N__5910));
    Sp12to4 I__503 (
            .O(N__5910),
            .I(N__5907));
    Span12Mux_s7_v I__502 (
            .O(N__5907),
            .I(N__5904));
    Odrv12 I__501 (
            .O(N__5904),
            .I(wRamRdData_1));
    IoInMux I__500 (
            .O(N__5901),
            .I(N__5898));
    LocalMux I__499 (
            .O(N__5898),
            .I(N__5895));
    Sp12to4 I__498 (
            .O(N__5895),
            .I(N__5892));
    Span12Mux_v I__497 (
            .O(N__5892),
            .I(N__5889));
    Odrv12 I__496 (
            .O(N__5889),
            .I(wRamRdData_6));
    IoInMux I__495 (
            .O(N__5886),
            .I(N__5883));
    LocalMux I__494 (
            .O(N__5883),
            .I(N__5880));
    Span4Mux_s3_v I__493 (
            .O(N__5880),
            .I(N__5877));
    Span4Mux_v I__492 (
            .O(N__5877),
            .I(N__5874));
    Odrv4 I__491 (
            .O(N__5874),
            .I(wRamRdData_2));
    IoInMux I__490 (
            .O(N__5871),
            .I(N__5868));
    LocalMux I__489 (
            .O(N__5868),
            .I(N__5865));
    Span12Mux_s6_v I__488 (
            .O(N__5865),
            .I(N__5862));
    Odrv12 I__487 (
            .O(N__5862),
            .I(wRamRdData_5));
    defparam IN_MUX_bfv_14_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_2_0_));
    defparam IN_MUX_bfv_14_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_3_0_ (
            .carryinitin(\DUT.uart_inst0.tx_clk_divider_cry_7 ),
            .carryinitout(bfn_14_3_0_));
    defparam IN_MUX_bfv_13_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_7_0_));
    defparam IN_MUX_bfv_13_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_8_0_ (
            .carryinitin(\DUT.uart_inst0.rx_clk_divider_1_cry_7 ),
            .carryinitout(bfn_13_8_0_));
    defparam IN_MUX_bfv_13_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_9_0_ (
            .carryinitin(\DUT.uart_inst0.rx_clk_divider_1_cry_15 ),
            .carryinitout(bfn_13_9_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_18_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_12_0_));
    defparam IN_MUX_bfv_15_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_9_0_));
    ICE_GB \top_pll_inst.top_pll_inst_RNISDA2_1  (
            .USERSIGNALTOGLOBALBUFFER(N__5967),
            .GLOBALBUFFEROUTPUT(wPllLocked_iso_i_g));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB \top_pll_inst.top_pll_inst_RNISDA2  (
            .USERSIGNALTOGLOBALBUFFER(N__10822),
            .GLOBALBUFFEROUTPUT(wPllLocked_g));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0 .C_ON=1'b0;
    defparam \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0 .SEQ_MODE=4'b0000;
    defparam \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5973),
            .lcout(wPllLocked),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.oPacketAvail_latch_LC_12_7_3 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.oPacketAvail_latch_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.oPacketAvail_latch_LC_12_7_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_inst.ftdi_input_inst.oPacketAvail_latch_LC_12_7_3  (
            .in0(N__14548),
            .in1(N__14588),
            .in2(_gnd_net_),
            .in3(N__7809),
            .lcout(G_120),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \top_pll_inst.top_pll_inst_RNISDA2_0_LC_12_30_3 .C_ON=1'b0;
    defparam \top_pll_inst.top_pll_inst_RNISDA2_0_LC_12_30_3 .SEQ_MODE=4'b0000;
    defparam \top_pll_inst.top_pll_inst_RNISDA2_0_LC_12_30_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \top_pll_inst.top_pll_inst_RNISDA2_0_LC_12_30_3  (
            .in0(N__14574),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\top_pll_inst.wPllLocked_iso_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_0_2_LC_13_2_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_0_2_LC_13_2_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_0_2_LC_13_2_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_0_2_LC_13_2_0  (
            .in0(N__6484),
            .in1(N__6459),
            .in2(N__6428),
            .in3(N__6670),
            .lcout(\DUT.uart_inst0.N_159_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNI92K37_0_LC_13_2_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNI92K37_0_LC_13_2_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNI92K37_0_LC_13_2_1 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \DUT.uart_inst0.tx_state_RNI92K37_0_LC_13_2_1  (
            .in0(N__6885),
            .in1(N__6057),
            .in2(N__8307),
            .in3(N__7014),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_6_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNINQKO8_1_LC_13_2_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNINQKO8_1_LC_13_2_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNINQKO8_1_LC_13_2_2 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \DUT.uart_inst0.tx_state_RNINQKO8_1_LC_13_2_2  (
            .in0(N__10787),
            .in1(N__8394),
            .in2(N__6024),
            .in3(N__6216),
            .lcout(\DUT.uart_inst0.N_22 ),
            .ltout(\DUT.uart_inst0.N_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_1_LC_13_2_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_1_LC_13_2_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_bits_remaining_1_LC_13_2_3 .LUT_INIT=16'b1111110000000011;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_1_LC_13_2_3  (
            .in0(_gnd_net_),
            .in1(N__6422),
            .in2(N__6021),
            .in3(N__6464),
            .lcout(\DUT.uart_inst0.tx_bits_remainingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15035),
            .ce(),
            .sr(N__6606));
    defparam \DUT.uart_inst0.tx_bits_remaining_2_LC_13_2_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_2_LC_13_2_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_bits_remaining_2_LC_13_2_4 .LUT_INIT=16'b1010101010101001;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_2_LC_13_2_4  (
            .in0(N__6485),
            .in1(N__6460),
            .in2(N__6018),
            .in3(N__6426),
            .lcout(\DUT.uart_inst0.tx_bits_remainingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15035),
            .ce(),
            .sr(N__6606));
    defparam \DUT.uart_inst0.tx_bits_remaining_0_LC_13_2_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_0_LC_13_2_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_bits_remaining_0_LC_13_2_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_0_LC_13_2_5  (
            .in0(_gnd_net_),
            .in1(N__6421),
            .in2(_gnd_net_),
            .in3(N__6014),
            .lcout(\DUT.uart_inst0.tx_bits_remainingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15035),
            .ce(),
            .sr(N__6606));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_2_LC_13_2_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_2_LC_13_2_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_2_LC_13_2_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_2_LC_13_2_6  (
            .in0(N__6483),
            .in1(N__6458),
            .in2(N__6427),
            .in3(N__6669),
            .lcout(\DUT.uart_inst0.N_159 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_RNI2V95_2_LC_13_3_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI2V95_2_LC_13_3_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI2V95_2_LC_13_3_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNI2V95_2_LC_13_3_0  (
            .in0(N__6320),
            .in1(N__6335),
            .in2(N__6354),
            .in3(N__6305),
            .lcout(\DUT.uart_inst0.un1_tx_clk_divider_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_13_LC_13_3_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_13_LC_13_3_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_13_LC_13_3_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_13_LC_13_3_1  (
            .in0(N__6521),
            .in1(N__6275),
            .in2(N__6504),
            .in3(N__6290),
            .lcout(\DUT.uart_inst0.un1_tx_clk_divider_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_8_LC_13_3_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_8_LC_13_3_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_8_LC_13_3_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_8_LC_13_3_2  (
            .in0(N__6554),
            .in1(N__6245),
            .in2(N__6540),
            .in3(N__6260),
            .lcout(\DUT.uart_inst0.un1_tx_clk_divider_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNI01HK1_5_LC_13_3_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNI01HK1_5_LC_13_3_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNI01HK1_5_LC_13_3_3 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNI01HK1_5_LC_13_3_3  (
            .in0(N__7127),
            .in1(N__6846),
            .in2(N__7335),
            .in3(N__7082),
            .lcout(),
            .ltout(\DUT.uart_inst0.g2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNIJKPE2_4_LC_13_3_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNIJKPE2_4_LC_13_3_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNIJKPE2_4_LC_13_3_4 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNIJKPE2_4_LC_13_3_4  (
            .in0(N__6740),
            .in1(_gnd_net_),
            .in2(N__6060),
            .in3(N__6792),
            .lcout(\DUT.uart_inst0.g2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_1_LC_13_3_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_1_LC_13_3_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_1_LC_13_3_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \DUT.uart_inst0.tx_countdown_1_LC_13_3_5  (
            .in0(N__7128),
            .in1(N__6618),
            .in2(_gnd_net_),
            .in3(N__7363),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15029),
            .ce(N__14421),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_RNIBPK2_0_LC_13_4_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNIBPK2_0_LC_13_4_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNIBPK2_0_LC_13_4_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNIBPK2_0_LC_13_4_0  (
            .in0(N__6372),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8543),
            .lcout(),
            .ltout(\DUT.uart_inst0.un1_tx_clk_divider_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_RNITC2S1_0_LC_13_4_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNITC2S1_0_LC_13_4_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNITC2S1_0_LC_13_4_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNITC2S1_0_LC_13_4_1  (
            .in0(N__6051),
            .in1(N__6045),
            .in2(N__6039),
            .in3(N__6036),
            .lcout(\DUT.uart_inst0.un1_tx_clk_divider_0 ),
            .ltout(\DUT.uart_inst0.un1_tx_clk_divider_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNI3MLP6_0_LC_13_4_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNI3MLP6_0_LC_13_4_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNI3MLP6_0_LC_13_4_2 .LUT_INIT=16'b0111111101110000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNI3MLP6_0_LC_13_4_2  (
            .in0(N__6695),
            .in1(N__6938),
            .in2(N__6030),
            .in3(N__6881),
            .lcout(\DUT.uart_inst0.N_109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_13_4_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_13_4_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_13_4_3 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_13_4_3  (
            .in0(N__7001),
            .in1(N__6636),
            .in2(N__6093),
            .in3(N__8303),
            .lcout(\DUT.uart_inst0.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNIMDQK4_0_0_LC_13_4_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNIMDQK4_0_0_LC_13_4_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNIMDQK4_0_0_LC_13_4_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \DUT.uart_inst0.tx_state_RNIMDQK4_0_0_LC_13_4_4  (
            .in0(N__8302),
            .in1(N__6880),
            .in2(_gnd_net_),
            .in3(N__6998),
            .lcout(\DUT.uart_inst0.N_152 ),
            .ltout(\DUT.uart_inst0.N_152_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNIBVOQB_1_LC_13_4_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNIBVOQB_1_LC_13_4_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNIBVOQB_1_LC_13_4_5 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \DUT.uart_inst0.tx_state_RNIBVOQB_1_LC_13_4_5  (
            .in0(N__7000),
            .in1(N__6629),
            .in2(N__6027),
            .in3(N__6678),
            .lcout(\DUT.uart_inst0.tx_countdown_7_sm0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_3_LC_13_4_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_3_LC_13_4_6 .SEQ_MODE=4'b1001;
    defparam \DUT.uart_inst0.tx_bits_remaining_3_LC_13_4_6 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_3_LC_13_4_6  (
            .in0(N__6081),
            .in1(N__6438),
            .in2(N__6672),
            .in3(N__6387),
            .lcout(\DUT.uart_inst0.tx_bits_remainingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15023),
            .ce(),
            .sr(N__6605));
    defparam \DUT.uart_inst0.tx_state_RNISP995_0_LC_13_4_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNISP995_0_LC_13_4_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNISP995_0_LC_13_4_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \DUT.uart_inst0.tx_state_RNISP995_0_LC_13_4_7  (
            .in0(N__6999),
            .in1(N__6696),
            .in2(N__6939),
            .in3(N__6580),
            .lcout(\DUT.uart_inst0.N_120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNIDD8Q_0_LC_13_5_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNIDD8Q_0_LC_13_5_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNIDD8Q_0_LC_13_5_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNIDD8Q_0_LC_13_5_0  (
            .in0(N__7121),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7071),
            .lcout(\DUT.uart_inst0.tx_countdown_0_ac0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_2_2_LC_13_5_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_2_2_LC_13_5_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_2_2_LC_13_5_1 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_2_2_LC_13_5_1  (
            .in0(N__7072),
            .in1(N__6788),
            .in2(N__6741),
            .in3(N__7122),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_countdown_7_m1_0_o2_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_2_LC_13_5_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_2_LC_13_5_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_2_LC_13_5_2 .LUT_INIT=16'b1111111110101000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_1_2_LC_13_5_2  (
            .in0(N__8273),
            .in1(N__7397),
            .in2(N__6075),
            .in3(N__6630),
            .lcout(\DUT.uart_inst0.N_113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNILLC71_2_LC_13_5_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNILLC71_2_LC_13_5_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNILLC71_2_LC_13_5_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNILLC71_2_LC_13_5_3  (
            .in0(N__7070),
            .in1(N__7120),
            .in2(_gnd_net_),
            .in3(N__7321),
            .lcout(\DUT.uart_inst0.tx_countdown_0_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_RNO_1_LC_13_5_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_RNO_1_LC_13_5_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_out_RNO_1_LC_13_5_4 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \DUT.uart_inst0.tx_out_RNO_1_LC_13_5_4  (
            .in0(N__6911),
            .in1(N__7797),
            .in2(N__8298),
            .in3(N__8390),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_out_6_iv_0_a3_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_RNO_0_LC_13_5_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_RNO_0_LC_13_5_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_out_RNO_0_LC_13_5_5 .LUT_INIT=16'b1110111011111110;
    LogicCell40 \DUT.uart_inst0.tx_out_RNO_0_LC_13_5_5  (
            .in0(N__7734),
            .in1(N__6066),
            .in2(N__6072),
            .in3(N__7141),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_out_6_iv_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_LC_13_5_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_LC_13_5_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_out_LC_13_5_6 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \DUT.uart_inst0.tx_out_LC_13_5_6  (
            .in0(N__7142),
            .in1(N__7768),
            .in2(N__6069),
            .in3(N__8272),
            .lcout(P1A7_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15017),
            .ce(N__14428),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_RNO_3_LC_13_5_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_RNO_3_LC_13_5_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_out_RNO_3_LC_13_5_7 .LUT_INIT=16'b1100010000000100;
    LogicCell40 \DUT.uart_inst0.tx_out_RNO_3_LC_13_5_7  (
            .in0(N__9425),
            .in1(N__7758),
            .in2(N__8297),
            .in3(N__6910),
            .lcout(\DUT.uart_inst0.N_119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_0_LC_13_6_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_0_LC_13_6_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_0_LC_13_6_0 .LUT_INIT=16'b0100010000100010;
    LogicCell40 \DUT.uart_inst0.tx_countdown_0_LC_13_6_0  (
            .in0(N__6959),
            .in1(N__7069),
            .in2(_gnd_net_),
            .in3(N__7364),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15012),
            .ce(N__14435),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_4_LC_13_6_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_4_LC_13_6_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_4_LC_13_6_1 .LUT_INIT=16'b1100100100000000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_0_4_LC_13_6_1  (
            .in0(N__6784),
            .in1(N__6732),
            .in2(N__6810),
            .in3(N__6958),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_countdown_RNO_0Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_4_LC_13_6_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_4_LC_13_6_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_4_LC_13_6_2 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_4_LC_13_6_2  (
            .in0(N__6733),
            .in1(_gnd_net_),
            .in2(N__6102),
            .in3(N__7365),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15012),
            .ce(N__14435),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNI34HK1_5_LC_13_6_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNI34HK1_5_LC_13_6_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNI34HK1_5_LC_13_6_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNI34HK1_5_LC_13_6_3  (
            .in0(N__6837),
            .in1(N__6730),
            .in2(N__7081),
            .in3(N__7319),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNIJKPE2_1_LC_13_6_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNIJKPE2_1_LC_13_6_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNIJKPE2_1_LC_13_6_4 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNIJKPE2_1_LC_13_6_4  (
            .in0(_gnd_net_),
            .in1(N__6780),
            .in2(N__6099),
            .in3(N__7123),
            .lcout(\DUT.uart_inst0.N_100 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_5_3_LC_13_6_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_5_3_LC_13_6_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_5_3_LC_13_6_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNO_5_3_LC_13_6_5  (
            .in0(N__6838),
            .in1(N__7320),
            .in2(N__6791),
            .in3(N__6731),
            .lcout(),
            .ltout(\DUT.uart_inst0.m25_e_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_3_3_LC_13_6_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_3_3_LC_13_6_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_3_3_LC_13_6_6 .LUT_INIT=16'b1100110001001100;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNO_3_3_LC_13_6_6  (
            .in0(N__7076),
            .in1(N__6671),
            .in2(N__6096),
            .in3(N__7124),
            .lcout(\DUT.uart_inst0.m3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_5_LC_13_6_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_5_LC_13_6_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_5_LC_13_6_7 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_5_LC_13_6_7  (
            .in0(N__7366),
            .in1(N__6960),
            .in2(N__7401),
            .in3(N__6842),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15012),
            .ce(N__14435),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_13_7_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_13_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_13_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8136),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_7_0_),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_13_7_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_13_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_13_7_1  (
            .in0(_gnd_net_),
            .in1(N__8106),
            .in2(N__9180),
            .in3(N__6129),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_0 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_13_7_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_13_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_13_7_2  (
            .in0(_gnd_net_),
            .in1(N__8079),
            .in2(N__9188),
            .in3(N__6126),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_1 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_3_LC_13_7_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_3_LC_13_7_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_3_LC_13_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNO_0_3_LC_13_7_3  (
            .in0(_gnd_net_),
            .in1(N__8052),
            .in2(N__9182),
            .in3(N__6123),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_3 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_2 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_13_7_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_13_7_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_13_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_13_7_4  (
            .in0(_gnd_net_),
            .in1(N__8463),
            .in2(N__9189),
            .in3(N__6120),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_3 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_5_LC_13_7_5 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_5_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_5_LC_13_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNO_0_5_LC_13_7_5  (
            .in0(_gnd_net_),
            .in1(N__7488),
            .in2(N__9183),
            .in3(N__6117),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_5 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_4 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_6_LC_13_7_6 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_6_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_6_LC_13_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNO_0_6_LC_13_7_6  (
            .in0(_gnd_net_),
            .in1(N__7470),
            .in2(N__9190),
            .in3(N__6114),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_6 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_5 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_13_7_7 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_13_7_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_13_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_13_7_7  (
            .in0(_gnd_net_),
            .in1(N__7511),
            .in2(N__9181),
            .in3(N__6111),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_6 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_13_8_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_13_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_13_8_0  (
            .in0(_gnd_net_),
            .in1(N__7451),
            .in2(N__9186),
            .in3(N__6108),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_13_8_0_),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_13_8_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_13_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_13_8_1  (
            .in0(_gnd_net_),
            .in1(N__7161),
            .in2(N__9194),
            .in3(N__6105),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_8 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_LUT4_0_LC_13_8_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_LUT4_0_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_LUT4_0_LC_13_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_LUT4_0_LC_13_8_2  (
            .in0(_gnd_net_),
            .in1(N__7185),
            .in2(N__9187),
            .in3(N__6153),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_9 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_LUT4_0_LC_13_8_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_LUT4_0_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_LUT4_0_LC_13_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_LUT4_0_LC_13_8_3  (
            .in0(_gnd_net_),
            .in1(N__7538),
            .in2(N__9191),
            .in3(N__6150),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_10 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_LUT4_0_LC_13_8_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_LUT4_0_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_LUT4_0_LC_13_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_LUT4_0_LC_13_8_4  (
            .in0(_gnd_net_),
            .in1(N__7426),
            .in2(N__9184),
            .in3(N__6147),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_11 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_LUT4_0_LC_13_8_5 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_LUT4_0_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_LUT4_0_LC_13_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_LUT4_0_LC_13_8_5  (
            .in0(_gnd_net_),
            .in1(N__7259),
            .in2(N__9192),
            .in3(N__6144),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_12 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_LUT4_0_LC_13_8_6 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_LUT4_0_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_LUT4_0_LC_13_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_LUT4_0_LC_13_8_6  (
            .in0(_gnd_net_),
            .in1(N__7232),
            .in2(N__9185),
            .in3(N__6141),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_13 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_LUT4_0_LC_13_8_7 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_LUT4_0_LC_13_8_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_LUT4_0_LC_13_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_LUT4_0_LC_13_8_7  (
            .in0(_gnd_net_),
            .in1(N__7209),
            .in2(N__9193),
            .in3(N__6138),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_14 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_LUT4_0_LC_13_9_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_LUT4_0_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_LUT4_0_LC_13_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_LUT4_0_LC_13_9_0  (
            .in0(_gnd_net_),
            .in1(N__8156),
            .in2(N__9195),
            .in3(N__6135),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_13_9_0_),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_17_LC_13_9_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_17_LC_13_9_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_17_LC_13_9_1 .LUT_INIT=16'b1011000000001011;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_17_LC_13_9_1  (
            .in0(N__10518),
            .in1(N__11013),
            .in2(N__7286),
            .in3(N__6132),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15000),
            .ce(N__14450),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_13_10_0 .C_ON=1'b1;
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_13_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(N__6195),
            .in2(N__9469),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_13_10_0_),
            .carryout(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_1_LC_13_10_1 .C_ON=1'b1;
    defparam \DUT.fifo_tx_inst.rFifoCount_1_LC_13_10_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoCount_1_LC_13_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_1_LC_13_10_1  (
            .in0(_gnd_net_),
            .in1(N__6204),
            .in2(N__9511),
            .in3(N__6210),
            .lcout(\DUT.fifo_tx_inst.rFifoCountZ0Z_1 ),
            .ltout(),
            .carryin(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0 ),
            .carryout(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1 ),
            .clk(N__14997),
            .ce(),
            .sr(N__15219));
    defparam \DUT.fifo_tx_inst.rFifoCount_2_LC_13_10_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_2_LC_13_10_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoCount_2_LC_13_10_2 .LUT_INIT=16'b0110001110011100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_2_LC_13_10_2  (
            .in0(N__6189),
            .in1(N__9325),
            .in2(N__9434),
            .in3(N__6207),
            .lcout(\DUT.fifo_tx_inst.rFifoCountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14997),
            .ce(),
            .sr(N__15219));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNISSQ21_1_LC_13_11_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNISSQ21_1_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNISSQ21_1_LC_13_11_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNISSQ21_1_LC_13_11_0  (
            .in0(N__9496),
            .in1(N__9430),
            .in2(_gnd_net_),
            .in3(N__6187),
            .lcout(\DUT.fifo_tx_inst.rFifoCount_RNISSQ21Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNI0AJL_0_LC_13_11_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNI0AJL_0_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNI0AJL_0_LC_13_11_1 .LUT_INIT=16'b1111000011110001;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNI0AJL_0_LC_13_11_1  (
            .in0(N__9318),
            .in1(N__9495),
            .in2(N__6173),
            .in3(N__9455),
            .lcout(\DUT.fifo_tx_inst.N_108 ),
            .ltout(\DUT.fifo_tx_inst.N_108_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_13_11_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_13_11_2 .LUT_INIT=16'b0000110000111111;
    LogicCell40 \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_13_11_2  (
            .in0(N__9457),
            .in1(N__9429),
            .in2(N__6198),
            .in3(N__12238),
            .lcout(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_2_1_LC_13_11_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_2_1_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_2_1_LC_13_11_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_2_1_LC_13_11_3  (
            .in0(N__9319),
            .in1(N__12311),
            .in2(N__6174),
            .in3(N__12263),
            .lcout(\DUT.fifo_tx_inst.rFifoData_awe3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_0_LC_13_11_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_0_LC_13_11_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoCount_0_LC_13_11_4 .LUT_INIT=16'b1001101010010101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_0_LC_13_11_4  (
            .in0(N__9456),
            .in1(N__6188),
            .in2(N__9435),
            .in3(N__12239),
            .lcout(\DUT.fifo_tx_inst.rFifoCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14995),
            .ce(),
            .sr(N__15218));
    defparam rTxWrite_LC_13_11_5.C_ON=1'b0;
    defparam rTxWrite_LC_13_11_5.SEQ_MODE=4'b1000;
    defparam rTxWrite_LC_13_11_5.LUT_INIT=16'b1100110011111111;
    LogicCell40 rTxWrite_LC_13_11_5 (
            .in0(_gnd_net_),
            .in1(N__14824),
            .in2(_gnd_net_),
            .in3(N__12549),
            .lcout(rTxWriteZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14995),
            .ce(),
            .sr(N__15218));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNI7FOF_2_LC_13_11_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNI7FOF_2_LC_13_11_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNI7FOF_2_LC_13_11_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNI7FOF_2_LC_13_11_6  (
            .in0(_gnd_net_),
            .in1(N__6166),
            .in2(_gnd_net_),
            .in3(N__9317),
            .lcout(\DUT.fifo_tx_inst.N_104 ),
            .ltout(\DUT.fifo_tx_inst.N_104_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_0_1_LC_13_11_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_0_1_LC_13_11_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_0_1_LC_13_11_7 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_0_1_LC_13_11_7  (
            .in0(_gnd_net_),
            .in1(N__12312),
            .in2(N__6156),
            .in3(N__12264),
            .lcout(\DUT.fifo_tx_inst.rFifoData_awe1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_13_12_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_13_12_1 .LUT_INIT=16'b1010111110001101;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_13_12_1  (
            .in0(N__10708),
            .in1(N__10170),
            .in2(N__9210),
            .in3(N__10296),
            .lcout(),
            .ltout(\DUT.uart_inst0.rx_countdown_8_i_o2_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_2_LC_13_12_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_2_LC_13_12_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_2_LC_13_12_2 .LUT_INIT=16'b1100110011001110;
    LogicCell40 \DUT.uart_inst0.rx_countdown_2_LC_13_12_2  (
            .in0(N__7617),
            .in1(N__6231),
            .in2(N__6234),
            .in3(N__8907),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14994),
            .ce(N__14460),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_5_2_LC_13_12_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_5_2_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_5_2_LC_13_12_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_5_2_LC_13_12_3  (
            .in0(N__11568),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11117),
            .lcout(\DUT.uart_inst0.m4_e_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_2_2_LC_13_12_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_2_2_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_2_2_LC_13_12_4 .LUT_INIT=16'b1110000000100000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_2_2_LC_13_12_4  (
            .in0(N__11119),
            .in1(N__10707),
            .in2(N__10851),
            .in3(N__10001),
            .lcout(\DUT.uart_inst0.N_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNIUMLT1_5_LC_13_12_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNIUMLT1_5_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNIUMLT1_5_LC_13_12_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNIUMLT1_5_LC_13_12_5  (
            .in0(N__11489),
            .in1(N__11245),
            .in2(N__11574),
            .in3(N__11118),
            .lcout(),
            .ltout(\DUT.uart_inst0.g0_0_0_a3_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNI7CGS2_1_LC_13_12_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNI7CGS2_1_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNI7CGS2_1_LC_13_12_6 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNI7CGS2_1_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(N__11400),
            .in2(N__6225),
            .in3(N__10101),
            .lcout(\DUT.uart_inst0.g0_0_0_a3_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_3_1_LC_13_12_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_3_1_LC_13_12_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_3_1_LC_13_12_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_3_1_LC_13_12_7  (
            .in0(N__11488),
            .in1(N__11244),
            .in2(N__11573),
            .in3(N__11116),
            .lcout(\DUT.uart_inst0.N_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNIBTN81_0_LC_14_1_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNIBTN81_0_LC_14_1_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNIBTN81_0_LC_14_1_6 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \DUT.uart_inst0.tx_state_RNIBTN81_0_LC_14_1_6  (
            .in0(N__9416),
            .in1(N__8300),
            .in2(_gnd_net_),
            .in3(N__6222),
            .lcout(\DUT.uart_inst0.N_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_14_2_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_14_2_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_14_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_14_2_0  (
            .in0(_gnd_net_),
            .in1(N__8547),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_2_0_),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_1_LC_14_2_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_1_LC_14_2_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_1_LC_14_2_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_1_LC_14_2_1  (
            .in0(_gnd_net_),
            .in1(N__6371),
            .in2(N__9054),
            .in3(N__6357),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_1 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_0 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_1 ),
            .clk(N__15043),
            .ce(),
            .sr(N__8514));
    defparam \DUT.uart_inst0.tx_clk_divider_2_LC_14_2_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_2_LC_14_2_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_2_LC_14_2_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_2_LC_14_2_2  (
            .in0(_gnd_net_),
            .in1(N__6353),
            .in2(N__9058),
            .in3(N__6339),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_2 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_1 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_2 ),
            .clk(N__15043),
            .ce(),
            .sr(N__8514));
    defparam \DUT.uart_inst0.tx_clk_divider_3_LC_14_2_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_3_LC_14_2_3 .SEQ_MODE=4'b1001;
    defparam \DUT.uart_inst0.tx_clk_divider_3_LC_14_2_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_3_LC_14_2_3  (
            .in0(_gnd_net_),
            .in1(N__6336),
            .in2(N__9055),
            .in3(N__6324),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_3 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_2 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_3 ),
            .clk(N__15043),
            .ce(),
            .sr(N__8514));
    defparam \DUT.uart_inst0.tx_clk_divider_4_LC_14_2_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_4_LC_14_2_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_4_LC_14_2_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_4_LC_14_2_4  (
            .in0(_gnd_net_),
            .in1(N__6321),
            .in2(N__9059),
            .in3(N__6309),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_4 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_3 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_4 ),
            .clk(N__15043),
            .ce(),
            .sr(N__8514));
    defparam \DUT.uart_inst0.tx_clk_divider_5_LC_14_2_5 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_5_LC_14_2_5 .SEQ_MODE=4'b1001;
    defparam \DUT.uart_inst0.tx_clk_divider_5_LC_14_2_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_5_LC_14_2_5  (
            .in0(_gnd_net_),
            .in1(N__6306),
            .in2(N__9056),
            .in3(N__6294),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_5 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_4 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_5 ),
            .clk(N__15043),
            .ce(),
            .sr(N__8514));
    defparam \DUT.uart_inst0.tx_clk_divider_6_LC_14_2_6 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_6_LC_14_2_6 .SEQ_MODE=4'b1001;
    defparam \DUT.uart_inst0.tx_clk_divider_6_LC_14_2_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_6_LC_14_2_6  (
            .in0(_gnd_net_),
            .in1(N__6291),
            .in2(N__9060),
            .in3(N__6279),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_6 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_5 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_6 ),
            .clk(N__15043),
            .ce(),
            .sr(N__8514));
    defparam \DUT.uart_inst0.tx_clk_divider_7_LC_14_2_7 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_7_LC_14_2_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_7_LC_14_2_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_7_LC_14_2_7  (
            .in0(_gnd_net_),
            .in1(N__6276),
            .in2(N__9057),
            .in3(N__6264),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_7 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_6 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_7 ),
            .clk(N__15043),
            .ce(),
            .sr(N__8514));
    defparam \DUT.uart_inst0.tx_clk_divider_8_LC_14_3_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_8_LC_14_3_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_8_LC_14_3_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_8_LC_14_3_0  (
            .in0(_gnd_net_),
            .in1(N__6261),
            .in2(N__9126),
            .in3(N__6249),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_8 ),
            .ltout(),
            .carryin(bfn_14_3_0_),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_8 ),
            .clk(N__15036),
            .ce(),
            .sr(N__8509));
    defparam \DUT.uart_inst0.tx_clk_divider_9_LC_14_3_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_9_LC_14_3_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_9_LC_14_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_9_LC_14_3_1  (
            .in0(_gnd_net_),
            .in1(N__6246),
            .in2(N__9128),
            .in3(N__6558),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_9 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_8 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_9 ),
            .clk(N__15036),
            .ce(),
            .sr(N__8509));
    defparam \DUT.uart_inst0.tx_clk_divider_10_LC_14_3_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_10_LC_14_3_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_10_LC_14_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_10_LC_14_3_2  (
            .in0(_gnd_net_),
            .in1(N__6555),
            .in2(N__9124),
            .in3(N__6543),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_10 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_9 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_10 ),
            .clk(N__15036),
            .ce(),
            .sr(N__8509));
    defparam \DUT.uart_inst0.tx_clk_divider_11_LC_14_3_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_11_LC_14_3_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_11_LC_14_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_11_LC_14_3_3  (
            .in0(_gnd_net_),
            .in1(N__6539),
            .in2(N__9127),
            .in3(N__6525),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_11 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_10 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_11 ),
            .clk(N__15036),
            .ce(),
            .sr(N__8509));
    defparam \DUT.uart_inst0.tx_clk_divider_12_LC_14_3_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_12_LC_14_3_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_12_LC_14_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_12_LC_14_3_4  (
            .in0(_gnd_net_),
            .in1(N__6522),
            .in2(N__9125),
            .in3(N__6510),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_12 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_11 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_12 ),
            .clk(N__15036),
            .ce(),
            .sr(N__8509));
    defparam \DUT.uart_inst0.tx_clk_divider_13_LC_14_3_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_13_LC_14_3_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_13_LC_14_3_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_13_LC_14_3_5  (
            .in0(_gnd_net_),
            .in1(N__6503),
            .in2(_gnd_net_),
            .in3(N__6507),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15036),
            .ce(),
            .sr(N__8509));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_1_3_LC_14_4_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_1_3_LC_14_4_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_1_3_LC_14_4_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNO_1_3_LC_14_4_0  (
            .in0(N__6489),
            .in1(N__6393),
            .in2(N__8386),
            .in3(N__6468),
            .lcout(\DUT.uart_inst0.m9_e_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_4_3_LC_14_4_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_4_3_LC_14_4_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_4_3_LC_14_4_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNO_4_3_LC_14_4_1  (
            .in0(N__14547),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6429),
            .lcout(\DUT.uart_inst0.m9_e_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNIMDQK4_0_LC_14_4_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNIMDQK4_0_LC_14_4_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNIMDQK4_0_LC_14_4_2 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \DUT.uart_inst0.tx_state_RNIMDQK4_0_LC_14_4_2  (
            .in0(N__6694),
            .in1(N__7008),
            .in2(N__8301),
            .in3(N__6934),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_state_0_sqmuxa_i_i_a3_c_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNI00K8B_0_LC_14_4_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNI00K8B_0_LC_14_4_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNI00K8B_0_LC_14_4_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_state_RNI00K8B_0_LC_14_4_3  (
            .in0(N__6386),
            .in1(N__7947),
            .in2(N__6375),
            .in3(N__6584),
            .lcout(\DUT.uart_inst0.N_22_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNICODU_0_LC_14_4_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNICODU_0_LC_14_4_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNICODU_0_LC_14_4_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \DUT.uart_inst0.tx_state_RNICODU_0_LC_14_4_4  (
            .in0(_gnd_net_),
            .in1(N__8279),
            .in2(_gnd_net_),
            .in3(N__6908),
            .lcout(\DUT.uart_inst0.N_160 ),
            .ltout(\DUT.uart_inst0.N_160_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNI6Q5N3_1_LC_14_4_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNI6Q5N3_1_LC_14_4_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNI6Q5N3_1_LC_14_4_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \DUT.uart_inst0.tx_state_RNI6Q5N3_1_LC_14_4_5  (
            .in0(N__6933),
            .in1(N__8365),
            .in2(N__6699),
            .in3(N__6693),
            .lcout(\DUT.uart_inst0.N_154 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_2_3_LC_14_4_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_2_3_LC_14_4_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_2_3_LC_14_4_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNO_2_3_LC_14_4_6  (
            .in0(N__9398),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6665),
            .lcout(\DUT.uart_inst0.N_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNIIAMI1_1_LC_14_4_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNIIAMI1_1_LC_14_4_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNIIAMI1_1_LC_14_4_7 .LUT_INIT=16'b1110110011101111;
    LogicCell40 \DUT.uart_inst0.tx_state_RNIIAMI1_1_LC_14_4_7  (
            .in0(N__6909),
            .in1(N__8364),
            .in2(N__8299),
            .in3(N__9399),
            .lcout(\DUT.uart_inst0.N_99 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNI5PJS2_1_LC_14_5_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNI5PJS2_1_LC_14_5_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNI5PJS2_1_LC_14_5_1 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \DUT.uart_inst0.tx_state_RNI5PJS2_1_LC_14_5_1  (
            .in0(N__7959),
            .in1(N__14549),
            .in2(_gnd_net_),
            .in3(N__7012),
            .lcout(\DUT.uart_inst0.N_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_1_LC_14_5_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_1_LC_14_5_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_1_LC_14_5_2 .LUT_INIT=16'b1000000000001000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_0_1_LC_14_5_2  (
            .in0(N__7010),
            .in1(N__7957),
            .in2(N__7083),
            .in3(N__7125),
            .lcout(\DUT.uart_inst0.tx_countdown_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNI8CH01_0_1_LC_14_5_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNI8CH01_0_1_LC_14_5_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNI8CH01_0_1_LC_14_5_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \DUT.uart_inst0.tx_state_RNI8CH01_0_1_LC_14_5_3  (
            .in0(N__7958),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14550),
            .lcout(\DUT.uart_inst0.N_88_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_0_LC_14_5_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_0_LC_14_5_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_state_0_LC_14_5_4 .LUT_INIT=16'b0000000000001110;
    LogicCell40 \DUT.uart_inst0.tx_state_0_LC_14_5_4  (
            .in0(N__8277),
            .in1(N__9397),
            .in2(N__8393),
            .in3(N__6564),
            .lcout(\DUT.tx_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15024),
            .ce(),
            .sr(N__15229));
    defparam \DUT.uart_inst0.tx_state_RNIOJJIA_0_LC_14_5_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNIOJJIA_0_LC_14_5_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNIOJJIA_0_LC_14_5_5 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \DUT.uart_inst0.tx_state_RNIOJJIA_0_LC_14_5_5  (
            .in0(N__6879),
            .in1(N__7028),
            .in2(N__6585),
            .in3(N__7011),
            .lcout(\DUT.uart_inst0.N_218 ),
            .ltout(\DUT.uart_inst0.N_218_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_1_LC_14_5_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_1_LC_14_5_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_state_1_LC_14_5_6 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \DUT.uart_inst0.tx_state_1_LC_14_5_6  (
            .in0(_gnd_net_),
            .in1(N__8382),
            .in2(N__7146),
            .in3(N__7143),
            .lcout(\DUT.tx_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15024),
            .ce(),
            .sr(N__15229));
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_2_LC_14_5_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_2_LC_14_5_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_2_LC_14_5_7 .LUT_INIT=16'b0001111000000000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_0_2_LC_14_5_7  (
            .in0(N__7126),
            .in1(N__7080),
            .in2(N__7331),
            .in3(N__7009),
            .lcout(\DUT.uart_inst0.tx_countdown_7_m1_0_a3_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_14_6_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_14_6_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_14_6_0  (
            .in0(N__6779),
            .in1(N__6852),
            .in2(_gnd_net_),
            .in3(N__7032),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_countdown_RNO_1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_3_LC_14_6_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_3_LC_14_6_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_3_LC_14_6_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \DUT.uart_inst0.tx_countdown_3_LC_14_6_1  (
            .in0(_gnd_net_),
            .in1(N__6945),
            .in2(N__7017),
            .in3(N__7367),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15018),
            .ce(N__14436),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNI9B9Q2_1_LC_14_6_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNI9B9Q2_1_LC_14_6_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNI9B9Q2_1_LC_14_6_2 .LUT_INIT=16'b1111110100000000;
    LogicCell40 \DUT.uart_inst0.tx_state_RNI9B9Q2_1_LC_14_6_2  (
            .in0(N__9408),
            .in1(N__8267),
            .in2(N__8391),
            .in3(N__7013),
            .lcout(\DUT.uart_inst0.N_164 ),
            .ltout(\DUT.uart_inst0.N_164_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_14_6_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_14_6_3 .LUT_INIT=16'b1010000001010000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_14_6_3  (
            .in0(N__6806),
            .in1(_gnd_net_),
            .in2(N__6948),
            .in3(N__6778),
            .lcout(\DUT.uart_inst0.tx_countdown_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNI67HK1_5_LC_14_6_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNI67HK1_5_LC_14_6_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNI67HK1_5_LC_14_6_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNI67HK1_5_LC_14_6_4  (
            .in0(N__6835),
            .in1(N__7317),
            .in2(N__6789),
            .in3(N__6728),
            .lcout(\DUT.uart_inst0.tx_state_ns_i_i_o2_a0_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_2_3_LC_14_6_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_2_3_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_2_3_LC_14_6_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_2_3_LC_14_6_5  (
            .in0(N__8268),
            .in1(N__6915),
            .in2(N__8392),
            .in3(N__6878),
            .lcout(\DUT.uart_inst0.N_163 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNIJKPE2_5_LC_14_6_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNIJKPE2_5_LC_14_6_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNIJKPE2_5_LC_14_6_6 .LUT_INIT=16'b1010101010101001;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNIJKPE2_5_LC_14_6_6  (
            .in0(N__6836),
            .in1(N__6805),
            .in2(N__6790),
            .in3(N__6729),
            .lcout(\DUT.uart_inst0.tx_countdown_30_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_2_LC_14_6_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_2_LC_14_6_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_2_LC_14_6_7 .LUT_INIT=16'b1010101000111111;
    LogicCell40 \DUT.uart_inst0.tx_countdown_2_LC_14_6_7  (
            .in0(N__7318),
            .in1(N__7386),
            .in2(N__7377),
            .in3(N__7368),
            .lcout(\DUT.uart_inst0.N_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15018),
            .ce(N__14436),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNI3ALC_17_LC_14_7_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI3ALC_17_LC_14_7_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI3ALC_17_LC_14_7_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNI3ALC_17_LC_14_7_0  (
            .in0(N__7207),
            .in1(N__7231),
            .in2(N__7287),
            .in3(N__7258),
            .lcout(\DUT.uart_inst0.un2_rx_clk_divider_a_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_13_LC_14_7_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_13_LC_14_7_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_13_LC_14_7_1 .LUT_INIT=16'b1000110000100011;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_13_LC_14_7_1  (
            .in0(N__10504),
            .in1(N__7260),
            .in2(N__11016),
            .in3(N__7266),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15013),
            .ce(N__14443),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_14_LC_14_7_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_14_LC_14_7_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_14_LC_14_7_2 .LUT_INIT=16'b1100001101000001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_14_LC_14_7_2  (
            .in0(N__11012),
            .in1(N__7242),
            .in2(N__7236),
            .in3(N__10505),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15013),
            .ce(N__14443),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_15_LC_14_7_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_15_LC_14_7_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_15_LC_14_7_3 .LUT_INIT=16'b1100010000110001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_15_LC_14_7_3  (
            .in0(N__11005),
            .in1(N__7215),
            .in2(N__10557),
            .in3(N__7208),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15013),
            .ce(N__14443),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_10_LC_14_7_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_10_LC_14_7_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_10_LC_14_7_4 .LUT_INIT=16'b1000010010100101;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_10_LC_14_7_4  (
            .in0(N__7184),
            .in1(N__10502),
            .in2(N__7194),
            .in3(N__11009),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15013),
            .ce(N__14443),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIB99J_10_LC_14_7_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIB99J_10_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIB99J_10_LC_14_7_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIB99J_10_LC_14_7_5  (
            .in0(N__7537),
            .in1(N__7183),
            .in2(N__7428),
            .in3(N__7159),
            .lcout(\DUT.uart_inst0.un2_rx_clk_divider_a_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_9_LC_14_7_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_9_LC_14_7_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_9_LC_14_7_6 .LUT_INIT=16'b1000010010100101;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_9_LC_14_7_6  (
            .in0(N__7160),
            .in1(N__10509),
            .in2(N__7170),
            .in3(N__11010),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15013),
            .ce(N__14443),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_11_LC_14_7_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_11_LC_14_7_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_11_LC_14_7_7 .LUT_INIT=16'b1000001011000011;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_11_LC_14_7_7  (
            .in0(N__10503),
            .in1(N__7539),
            .in2(N__7548),
            .in3(N__11011),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15013),
            .ce(N__14443),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNI6B671_5_LC_14_8_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI6B671_5_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI6B671_5_LC_14_8_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNI6B671_5_LC_14_8_0  (
            .in0(N__7510),
            .in1(N__7469),
            .in2(N__7452),
            .in3(N__7487),
            .lcout(\DUT.uart_inst0.un2_rx_clk_divider_a_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_7_LC_14_8_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_7_LC_14_8_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_7_LC_14_8_1 .LUT_INIT=16'b1100001101000001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_7_LC_14_8_1  (
            .in0(N__10995),
            .in1(N__7521),
            .in2(N__7515),
            .in3(N__10535),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15007),
            .ce(N__14451),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_5_LC_14_8_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_5_LC_14_8_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_5_LC_14_8_2 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_5_LC_14_8_2  (
            .in0(N__7494),
            .in1(N__10996),
            .in2(N__10562),
            .in3(N__10683),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15007),
            .ce(N__14451),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_6_LC_14_8_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_6_LC_14_8_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_6_LC_14_8_3 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_6_LC_14_8_3  (
            .in0(N__10682),
            .in1(N__10531),
            .in2(N__11014),
            .in3(N__7476),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15007),
            .ce(N__14451),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_8_LC_14_8_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_8_LC_14_8_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_8_LC_14_8_4 .LUT_INIT=16'b1010001001010001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_8_LC_14_8_4  (
            .in0(N__7450),
            .in1(N__10997),
            .in2(N__10563),
            .in3(N__7458),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15007),
            .ce(N__14451),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_12_LC_14_8_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_12_LC_14_8_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_12_LC_14_8_5 .LUT_INIT=16'b1000101001000101;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_12_LC_14_8_5  (
            .in0(N__7434),
            .in1(N__10526),
            .in2(N__11015),
            .in3(N__7427),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15007),
            .ce(N__14451),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_16_LC_14_8_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_16_LC_14_8_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_16_LC_14_8_6 .LUT_INIT=16'b1000001011000011;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_16_LC_14_8_6  (
            .in0(N__10527),
            .in1(N__7407),
            .in2(N__8163),
            .in3(N__11004),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15007),
            .ce(N__14451),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_LC_14_8_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_LC_14_8_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_3_LC_14_8_7 .LUT_INIT=16'b0000000011011101;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_LC_14_8_7  (
            .in0(N__10994),
            .in1(N__10536),
            .in2(_gnd_net_),
            .in3(N__7575),
            .lcout(\DUT.uart_inst0.rx_countdownZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15007),
            .ce(N__14451),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_6_2_LC_14_9_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_6_2_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_6_2_LC_14_9_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_6_2_LC_14_9_0  (
            .in0(_gnd_net_),
            .in1(N__10276),
            .in2(_gnd_net_),
            .in3(N__10157),
            .lcout(),
            .ltout(\DUT.uart_inst0.m7_e_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_3_2_LC_14_9_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_3_2_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_3_2_LC_14_9_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_3_2_LC_14_9_1  (
            .in0(N__9909),
            .in1(N__9984),
            .in2(N__7590),
            .in3(N__10218),
            .lcout(),
            .ltout(\DUT.uart_inst0.m7_e_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_2_LC_14_9_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_2_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_2_LC_14_9_2 .LUT_INIT=16'b0011111111011101;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_2_LC_14_9_2  (
            .in0(N__7554),
            .in1(N__10677),
            .in2(N__7587),
            .in3(N__10099),
            .lcout(),
            .ltout(\DUT.uart_inst0.m9_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_2_LC_14_9_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_2_LC_14_9_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_2_LC_14_9_3 .LUT_INIT=16'b1000000010001010;
    LogicCell40 \DUT.uart_inst0.recv_state_2_LC_14_9_3  (
            .in0(N__10812),
            .in1(N__8799),
            .in2(N__7584),
            .in3(N__7581),
            .lcout(DUT_uart_inst0_recv_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15003),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_1_2_LC_14_9_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_1_2_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_1_2_LC_14_9_4 .LUT_INIT=16'b1010001011110011;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_1_2_LC_14_9_4  (
            .in0(N__8619),
            .in1(N__8874),
            .in2(N__10482),
            .in3(N__8798),
            .lcout(\DUT.uart_inst0.N_11_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_3_1_LC_14_9_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_3_1_LC_14_9_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_3_1_LC_14_9_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_3_1_LC_14_9_5  (
            .in0(N__10275),
            .in1(N__9983),
            .in2(N__10168),
            .in3(N__10217),
            .lcout(\DUT.uart_inst0.g1_i_a4_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_3_LC_14_9_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_3_LC_14_9_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_3_LC_14_9_6 .LUT_INIT=16'b0000000100001101;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_0_3_LC_14_9_6  (
            .in0(N__11220),
            .in1(N__10676),
            .in2(N__10890),
            .in3(N__10158),
            .lcout(\DUT.uart_inst0.N_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_2_2_LC_14_9_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_2_2_LC_14_9_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_2_2_LC_14_9_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_2_2_LC_14_9_7  (
            .in0(N__11498),
            .in1(N__11219),
            .in2(N__7569),
            .in3(N__11399),
            .lcout(\DUT.uart_inst0.m4_e_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_1_LC_14_10_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_1_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_1_LC_14_10_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_0_1_LC_14_10_0  (
            .in0(N__7623),
            .in1(N__10695),
            .in2(_gnd_net_),
            .in3(N__7653),
            .lcout(\DUT.uart_inst0.N_13_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNI9JOT_0_LC_14_10_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNI9JOT_0_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNI9JOT_0_LC_14_10_1 .LUT_INIT=16'b0011110000001111;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNI9JOT_0_LC_14_10_1  (
            .in0(_gnd_net_),
            .in1(N__8637),
            .in2(N__8688),
            .in3(N__8783),
            .lcout(\DUT.uart_inst0.m5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_4_1_LC_14_10_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_4_1_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_4_1_LC_14_10_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_4_1_LC_14_10_2  (
            .in0(N__10271),
            .in1(N__10142),
            .in2(N__9995),
            .in3(N__10216),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_21_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_2_1_LC_14_10_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_2_1_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_2_1_LC_14_10_3 .LUT_INIT=16'b0000010111110101;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_2_1_LC_14_10_3  (
            .in0(N__8677),
            .in1(_gnd_net_),
            .in2(N__7656),
            .in3(N__7641),
            .lcout(\DUT.uart_inst0.N_21_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNIO2V22_1_LC_14_10_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNIO2V22_1_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNIO2V22_1_LC_14_10_4 .LUT_INIT=16'b0000000001110011;
    LogicCell40 \DUT.uart_inst0.recv_state_RNIO2V22_1_LC_14_10_4  (
            .in0(N__8784),
            .in1(N__8863),
            .in2(N__10567),
            .in3(N__7647),
            .lcout(\DUT.uart_inst0.N_6 ),
            .ltout(\DUT.uart_inst0.N_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_1_LC_14_10_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_1_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_1_LC_14_10_5 .LUT_INIT=16'b0000111101010101;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_1_1_LC_14_10_5  (
            .in0(N__8676),
            .in1(_gnd_net_),
            .in2(N__7635),
            .in3(N__7632),
            .lcout(\DUT.uart_inst0.N_18_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_0_LC_14_10_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_0_LC_14_10_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_bits_remaining_0_LC_14_10_6 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_0_LC_14_10_6  (
            .in0(N__8638),
            .in1(N__8865),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.uart_inst0.rx_bits_remainingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15001),
            .ce(N__8826),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_14_10_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_14_10_7 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_14_10_7  (
            .in0(N__8864),
            .in1(N__10547),
            .in2(_gnd_net_),
            .in3(N__8785),
            .lcout(\DUT.uart_inst0.N_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_1_1_LC_14_11_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_1_1_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_1_1_LC_14_11_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_1_1_LC_14_11_0  (
            .in0(N__11040),
            .in1(N__10093),
            .in2(N__7605),
            .in3(N__9926),
            .lcout(),
            .ltout(\DUT.uart_inst0.g1_i_a4_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_1_LC_14_11_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_1_LC_14_11_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_1_LC_14_11_1 .LUT_INIT=16'b0000110001000100;
    LogicCell40 \DUT.uart_inst0.recv_state_1_LC_14_11_1  (
            .in0(N__9819),
            .in1(N__8577),
            .in2(N__7593),
            .in3(N__10702),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14998),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNIS6O94_0_LC_14_11_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNIS6O94_0_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNIS6O94_0_LC_14_11_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNIS6O94_0_LC_14_11_2  (
            .in0(N__7677),
            .in1(N__10291),
            .in2(_gnd_net_),
            .in3(N__10229),
            .lcout(),
            .ltout(\DUT.uart_inst0.g0_0_0_a3_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNIL139C_1_LC_14_11_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNIL139C_1_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNIL139C_1_LC_14_11_3 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNIL139C_1_LC_14_11_3  (
            .in0(N__7686),
            .in1(N__7713),
            .in2(N__7680),
            .in3(N__10701),
            .lcout(\DUT.uart_inst0.recv_state_RNIL139CZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_3_6_LC_14_11_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_3_6_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_3_6_LC_14_11_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_3_6_LC_14_11_4  (
            .in0(N__10164),
            .in1(N__9925),
            .in2(N__10002),
            .in3(N__10290),
            .lcout(\DUT.uart_inst0.m13_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNI69LM2_0_LC_14_11_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNI69LM2_0_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNI69LM2_0_LC_14_11_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNI69LM2_0_LC_14_11_5  (
            .in0(N__9997),
            .in1(N__9913),
            .in2(N__10100),
            .in3(N__10163),
            .lcout(\DUT.uart_inst0.g0_0_0_a3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI4PUO_1_LC_14_11_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI4PUO_1_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI4PUO_1_LC_14_11_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_RNI4PUO_1_LC_14_11_6  (
            .in0(N__14561),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12659),
            .lcout(\DUT.fifo_tx_inst.un1_i11_i ),
            .ltout(\DUT.fifo_tx_inst.un1_i11_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_1_LC_14_11_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_1_LC_14_11_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rWritePtr_1_LC_14_11_7 .LUT_INIT=16'b0000110000000110;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_1_LC_14_11_7  (
            .in0(N__12315),
            .in1(N__12271),
            .in2(N__7671),
            .in3(N__12240),
            .lcout(\DUT.fifo_tx_inst.rWritePtrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14998),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_0_LC_14_12_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_0_LC_14_12_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rWritePtr_0_LC_14_12_0 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_0_LC_14_12_0  (
            .in0(N__12369),
            .in1(N__12179),
            .in2(_gnd_net_),
            .in3(N__7664),
            .lcout(\DUT.fifo_rx_inst.rWritePtrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14996),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_1_LC_14_12_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_1_LC_14_12_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rWritePtr_1_LC_14_12_1 .LUT_INIT=16'b0001010101000000;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_1_LC_14_12_1  (
            .in0(N__7665),
            .in1(N__12370),
            .in2(N__12183),
            .in3(N__12329),
            .lcout(\DUT.fifo_rx_inst.rWritePtrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14996),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI96D91_2_LC_14_12_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI96D91_2_LC_14_12_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI96D91_2_LC_14_12_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNI96D91_2_LC_14_12_2  (
            .in0(N__12328),
            .in1(N__12592),
            .in2(N__12374),
            .in3(N__13902),
            .lcout(\DUT.fifo_rx_inst.N_57 ),
            .ltout(\DUT.fifo_rx_inst.N_57_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI5KNB1_2_LC_14_12_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI5KNB1_2_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI5KNB1_2_LC_14_12_3 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNI5KNB1_2_LC_14_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7668),
            .in3(N__14562),
            .lcout(\DUT.fifo_rx_inst.un1_i11_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_2_6_LC_14_12_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_2_6_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_2_6_LC_14_12_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_2_6_LC_14_12_4  (
            .in0(N__10230),
            .in1(N__10791),
            .in2(N__10568),
            .in3(N__11337),
            .lcout(),
            .ltout(\DUT.uart_inst0.m13_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_6_LC_14_12_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_6_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_6_LC_14_12_5 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_6_LC_14_12_5  (
            .in0(N__10578),
            .in1(N__10097),
            .in2(N__7725),
            .in3(N__7722),
            .lcout(),
            .ltout(\DUT.uart_inst0.P19_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_6_LC_14_12_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_6_LC_14_12_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_6_LC_14_12_6 .LUT_INIT=16'b0011000010010000;
    LogicCell40 \DUT.uart_inst0.recv_state_6_LC_14_12_6  (
            .in0(N__10098),
            .in1(N__10710),
            .in2(N__7716),
            .in3(N__9927),
            .lcout(\DUT.wRcvd ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14996),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNIBTG71_1_LC_14_12_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNIBTG71_1_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNIBTG71_1_LC_14_12_7 .LUT_INIT=16'b1111010000000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNIBTG71_1_LC_14_12_7  (
            .in0(N__10548),
            .in1(N__8869),
            .in2(N__8808),
            .in3(N__14563),
            .lcout(\DUT.uart_inst0.g0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ioFifoData_iobuf_RNO_0_LC_15_2_0.C_ON=1'b0;
    defparam ioFifoData_iobuf_RNO_0_LC_15_2_0.SEQ_MODE=4'b0000;
    defparam ioFifoData_iobuf_RNO_0_LC_15_2_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 ioFifoData_iobuf_RNO_0_LC_15_2_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13836),
            .lcout(N_1257_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.oTxFull_0_LC_15_3_0 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.oTxFull_0_LC_15_3_0 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.oTxFull_0_LC_15_3_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_inst.ftdi_input_inst.oTxFull_0_LC_15_3_0  (
            .in0(N__7845),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7898),
            .lcout(fifo_inst_ftdi_input_inst_oTxFull_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_1_LC_15_3_1 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_1_LC_15_3_1 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_1_LC_15_3_1 .LUT_INIT=16'b0001001100100000;
    LogicCell40 \fifo_inst.ftdi_input_inst.rPacketCount_latch_1_LC_15_3_1  (
            .in0(N__7925),
            .in1(N__15285),
            .in2(N__7880),
            .in3(N__7846),
            .lcout(G_111),
            .ltout(G_111_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.SUM_2_LC_15_3_2 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.SUM_2_LC_15_3_2 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.SUM_2_LC_15_3_2 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \fifo_inst.ftdi_input_inst.SUM_2_LC_15_3_2  (
            .in0(N__7827),
            .in1(_gnd_net_),
            .in2(N__7692),
            .in3(N__7868),
            .lcout(),
            .ltout(\fifo_inst.ftdi_input_inst.SUMZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_2_LC_15_3_3 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_2_LC_15_3_3 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_2_LC_15_3_3 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \fifo_inst.ftdi_input_inst.rPacketCount_latch_2_LC_15_3_3  (
            .in0(N__7926),
            .in1(N__7828),
            .in2(N__7689),
            .in3(N__15286),
            .lcout(G_112),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_3_LC_15_3_4 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_3_LC_15_3_4 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_3_LC_15_3_4 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \fifo_inst.ftdi_input_inst.rPacketCount_latch_3_LC_15_3_4  (
            .in0(N__7924),
            .in1(N__7908),
            .in2(N__15291),
            .in3(N__7900),
            .lcout(G_109),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_0_LC_15_3_5 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_0_LC_15_3_5 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_0_LC_15_3_5 .LUT_INIT=16'b0000001100110000;
    LogicCell40 \fifo_inst.ftdi_input_inst.rPacketCount_latch_0_LC_15_3_5  (
            .in0(_gnd_net_),
            .in1(N__15284),
            .in2(N__7879),
            .in3(N__7923),
            .lcout(G_110),
            .ltout(G_110_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.wTxEn_1_LC_15_3_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.wTxEn_1_LC_15_3_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.wTxEn_1_LC_15_3_6 .LUT_INIT=16'b1100100011001100;
    LogicCell40 \DUT.fifo_tx_inst.wTxEn_1_LC_15_3_6  (
            .in0(N__7826),
            .in1(N__14546),
            .in2(N__7935),
            .in3(N__7932),
            .lcout(G_114),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.rPacketCount15_LC_15_3_7 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.rPacketCount15_LC_15_3_7 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.rPacketCount15_LC_15_3_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_inst.ftdi_input_inst.rPacketCount15_LC_15_3_7  (
            .in0(N__7899),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9570),
            .lcout(G_108),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.SUM_3_LC_15_4_1 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.SUM_3_LC_15_4_1 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.SUM_3_LC_15_4_1 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \fifo_inst.ftdi_input_inst.SUM_3_LC_15_4_1  (
            .in0(N__7829),
            .in1(N__7847),
            .in2(N__7881),
            .in3(N__7901),
            .lcout(\fifo_inst.ftdi_input_inst.SUMZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.un2_oPacketAvail_i_LC_15_4_2 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.un2_oPacketAvail_i_LC_15_4_2 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.un2_oPacketAvail_i_LC_15_4_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \fifo_inst.ftdi_input_inst.un2_oPacketAvail_i_LC_15_4_2  (
            .in0(N__7902),
            .in1(N__7878),
            .in2(N__7851),
            .in3(N__7830),
            .lcout(\fifo_inst.ftdi_input_inst.un2_oPacketAvail_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_7_LC_15_4_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_7_LC_15_4_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_7_LC_15_4_3 .LUT_INIT=16'b0000000000101010;
    LogicCell40 \DUT.uart_inst0.tx_data_7_LC_15_4_3  (
            .in0(N__8940),
            .in1(N__9609),
            .in2(N__9624),
            .in3(N__8278),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15037),
            .ce(N__7970),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_0_LC_15_5_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_0_LC_15_5_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_0_LC_15_5_0 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \DUT.uart_inst0.tx_data_0_LC_15_5_0  (
            .in0(N__8260),
            .in1(N__9273),
            .in2(N__8037),
            .in3(N__9588),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15030),
            .ce(N__7971),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_RNO_2_LC_15_5_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_RNO_2_LC_15_5_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_out_RNO_2_LC_15_5_1 .LUT_INIT=16'b1000000011000000;
    LogicCell40 \DUT.uart_inst0.tx_out_RNO_2_LC_15_5_1  (
            .in0(N__7790),
            .in1(N__8369),
            .in2(N__7778),
            .in3(N__8259),
            .lcout(\DUT.uart_inst0.N_116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_1_LC_15_5_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_1_LC_15_5_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_1_LC_15_5_2 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \DUT.uart_inst0.tx_data_1_LC_15_5_2  (
            .in0(N__8261),
            .in1(N__9249),
            .in2(N__8028),
            .in3(N__9589),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15030),
            .ce(N__7971),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_2_LC_15_5_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_2_LC_15_5_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_2_LC_15_5_3 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \DUT.uart_inst0.tx_data_2_LC_15_5_3  (
            .in0(N__9590),
            .in1(N__11760),
            .in2(N__8019),
            .in3(N__8264),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15030),
            .ce(N__7971),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_3_LC_15_5_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_3_LC_15_5_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_3_LC_15_5_4 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \DUT.uart_inst0.tx_data_3_LC_15_5_4  (
            .in0(N__8262),
            .in1(N__11589),
            .in2(N__8007),
            .in3(N__9591),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15030),
            .ce(N__7971),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_4_LC_15_5_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_4_LC_15_5_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_4_LC_15_5_5 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \DUT.uart_inst0.tx_data_4_LC_15_5_5  (
            .in0(N__9592),
            .in1(N__9240),
            .in2(N__7998),
            .in3(N__8265),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15030),
            .ce(N__7971),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_5_LC_15_5_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_5_LC_15_5_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_5_LC_15_5_6 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \DUT.uart_inst0.tx_data_5_LC_15_5_6  (
            .in0(N__8263),
            .in1(N__9543),
            .in2(N__7980),
            .in3(N__9593),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15030),
            .ce(N__7971),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_6_LC_15_5_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_6_LC_15_5_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_6_LC_15_5_7 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \DUT.uart_inst0.tx_data_6_LC_15_5_7  (
            .in0(N__9594),
            .in1(N__9519),
            .in2(N__7989),
            .in3(N__8266),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15030),
            .ce(N__7971),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNICU6U_1_LC_15_6_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNICU6U_1_LC_15_6_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNICU6U_1_LC_15_6_0 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \DUT.uart_inst0.tx_state_RNICU6U_1_LC_15_6_0  (
            .in0(N__8361),
            .in1(N__9372),
            .in2(_gnd_net_),
            .in3(N__8250),
            .lcout(\DUT.uart_inst0.N_102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.rWrState_latch_1_LC_15_6_2 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.rWrState_latch_1_LC_15_6_2 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.rWrState_latch_1_LC_15_6_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \fifo_inst.ftdi_input_inst.rWrState_latch_1_LC_15_6_2  (
            .in0(N__9754),
            .in1(N__14552),
            .in2(_gnd_net_),
            .in3(N__9730),
            .lcout(G_113),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNI8CH01_1_LC_15_6_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNI8CH01_1_LC_15_6_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNI8CH01_1_LC_15_6_4 .LUT_INIT=16'b1010111110111111;
    LogicCell40 \DUT.uart_inst0.tx_state_RNI8CH01_1_LC_15_6_4  (
            .in0(N__8362),
            .in1(N__9373),
            .in2(N__14575),
            .in3(N__8251),
            .lcout(\DUT.uart_inst0.tx_state_0_sqmuxa_i_i_a3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIN9O8_0_LC_15_6_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIN9O8_0_LC_15_6_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIN9O8_0_LC_15_6_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNIN9O8_0_LC_15_6_5  (
            .in0(N__9513),
            .in1(N__9477),
            .in2(_gnd_net_),
            .in3(N__9333),
            .lcout(),
            .ltout(\DUT.N_114_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.rTransmit_LC_15_6_6 .C_ON=1'b0;
    defparam \DUT.rTransmit_LC_15_6_6 .SEQ_MODE=4'b1000;
    defparam \DUT.rTransmit_LC_15_6_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \DUT.rTransmit_LC_15_6_6  (
            .in0(N__8363),
            .in1(N__14551),
            .in2(N__8310),
            .in3(N__8252),
            .lcout(\DUT.rTransmitZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15025),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_0_LC_15_7_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_0_LC_15_7_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_0_LC_15_7_0 .LUT_INIT=16'b1111111110110011;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_0_LC_15_7_0  (
            .in0(N__10953),
            .in1(N__14557),
            .in2(N__10558),
            .in3(N__12608),
            .lcout(\DUT.uart_inst0.G_19_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIMQ571_1_LC_15_7_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIMQ571_1_LC_15_7_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIMQ571_1_LC_15_7_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIMQ571_1_LC_15_7_1  (
            .in0(N__8048),
            .in1(N__8074),
            .in2(N__8462),
            .in3(N__8101),
            .lcout(),
            .ltout(\DUT.uart_inst0.un2_rx_clk_divider_a_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIJI4K1_16_LC_15_7_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIJI4K1_16_LC_15_7_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIJI4K1_16_LC_15_7_2 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIJI4K1_16_LC_15_7_2  (
            .in0(_gnd_net_),
            .in1(N__8155),
            .in2(N__8139),
            .in3(N__8128),
            .lcout(\DUT.uart_inst0.un2_rx_clk_divider_a_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_0_LC_15_7_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_0_LC_15_7_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_0_LC_15_7_3 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_0_LC_15_7_3  (
            .in0(N__8129),
            .in1(N__10513),
            .in2(_gnd_net_),
            .in3(N__10959),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15019),
            .ce(N__14452),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_LC_15_7_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_1_LC_15_7_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_LC_15_7_4 .LUT_INIT=16'b1000101001000101;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_LC_15_7_4  (
            .in0(N__8102),
            .in1(N__10519),
            .in2(N__10993),
            .in3(N__8115),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15019),
            .ce(N__14452),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_2_LC_15_7_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_2_LC_15_7_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_2_LC_15_7_5 .LUT_INIT=16'b1010001001010001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_2_LC_15_7_5  (
            .in0(N__8088),
            .in1(N__10955),
            .in2(N__10560),
            .in3(N__8075),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15019),
            .ce(N__14452),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_3_LC_15_7_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_3_LC_15_7_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_3_LC_15_7_6 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_3_LC_15_7_6  (
            .in0(N__10954),
            .in1(N__8061),
            .in2(N__10559),
            .in3(N__10686),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15019),
            .ce(N__14452),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_4_LC_15_7_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_4_LC_15_7_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_4_LC_15_7_7 .LUT_INIT=16'b1001000010011001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_4_LC_15_7_7  (
            .in0(N__8458),
            .in1(N__8475),
            .in2(N__10561),
            .in3(N__10960),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15019),
            .ce(N__14452),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNINK4E1_2_LC_15_8_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNINK4E1_2_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNINK4E1_2_LC_15_8_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNINK4E1_2_LC_15_8_0  (
            .in0(N__8787),
            .in1(N__11455),
            .in2(N__14576),
            .in3(N__11218),
            .lcout(),
            .ltout(\DUT.uart_inst0.m6_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNI3V794_0_LC_15_8_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNI3V794_0_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNI3V794_0_LC_15_8_1 .LUT_INIT=16'b0001010110111111;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNI3V794_0_LC_15_8_1  (
            .in0(N__10057),
            .in1(N__9771),
            .in2(N__8442),
            .in3(N__9903),
            .lcout(\DUT.uart_inst0.G_30_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \top_pll_inst.top_pll_inst_RNIIIF42_LC_15_8_2 .C_ON=1'b0;
    defparam \top_pll_inst.top_pll_inst_RNIIIF42_LC_15_8_2 .SEQ_MODE=4'b0000;
    defparam \top_pll_inst.top_pll_inst_RNIIIF42_LC_15_8_2 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \top_pll_inst.top_pll_inst_RNIIIF42_LC_15_8_2  (
            .in0(N__8788),
            .in1(N__10824),
            .in2(N__9921),
            .in3(N__9982),
            .lcout(),
            .ltout(\top_pll_inst.m12_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \top_pll_inst.top_pll_inst_RNI0MK94_LC_15_8_3 .C_ON=1'b0;
    defparam \top_pll_inst.top_pll_inst_RNI0MK94_LC_15_8_3 .SEQ_MODE=4'b0000;
    defparam \top_pll_inst.top_pll_inst_RNI0MK94_LC_15_8_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \top_pll_inst.top_pll_inst_RNI0MK94_LC_15_8_3  (
            .in0(N__10159),
            .in1(N__10277),
            .in2(N__8439),
            .in3(N__10219),
            .lcout(),
            .ltout(P18_mux_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNIEGJTC_0_LC_15_8_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNIEGJTC_0_LC_15_8_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNIEGJTC_0_LC_15_8_4 .LUT_INIT=16'b1000000000110001;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNIEGJTC_0_LC_15_8_4  (
            .in0(N__10065),
            .in1(N__8436),
            .in2(N__8430),
            .in3(N__10675),
            .lcout(\DUT.uart_inst0.rx_bits_remaining_2_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNI7H9R3_10_LC_15_8_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI7H9R3_10_LC_15_8_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI7H9R3_10_LC_15_8_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNI7H9R3_10_LC_15_8_5  (
            .in0(N__8427),
            .in1(N__8418),
            .in2(N__8412),
            .in3(N__8403),
            .lcout(\DUT.uart_inst0.un2_rx_clk_divider_0 ),
            .ltout(\DUT.uart_inst0.un2_rx_clk_divider_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNI15HA8_0_LC_15_8_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNI15HA8_0_LC_15_8_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNI15HA8_0_LC_15_8_6 .LUT_INIT=16'b1111001101111011;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNI15HA8_0_LC_15_8_6  (
            .in0(N__10064),
            .in1(N__9792),
            .in2(N__8397),
            .in3(N__9919),
            .lcout(\DUT.uart_inst0.rx_countdown_8_i_o2_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_4_3_LC_15_9_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.recv_state_RNO_4_3_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_4_3_LC_15_9_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_4_3_LC_15_9_0  (
            .in0(N__11149),
            .in1(N__10049),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.uart_inst0.m6_e_2 ),
            .ltout(),
            .carryin(bfn_15_9_0_),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_s1_c_RNIKPDT_LC_15_9_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_s1_c_RNIKPDT_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_s1_c_RNIKPDT_LC_15_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_0_s1_c_RNIKPDT_LC_15_9_1  (
            .in0(_gnd_net_),
            .in1(N__9113),
            .in2(N__11393),
            .in3(N__8562),
            .lcout(DUT_uart_inst0_rx_countdown_3_s1_1),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_countdown_3_cry_0_s1 ),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNIMVNN_LC_15_9_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNIMVNN_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNIMVNN_LC_15_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNIMVNN_LC_15_9_2  (
            .in0(_gnd_net_),
            .in1(N__9177),
            .in2(N__11156),
            .in3(N__8559),
            .lcout(DUT_uart_inst0_rx_countdown_3_s1_2),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_countdown_3_cry_1_s1 ),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_2_s1_c_RNIO52I_LC_15_9_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_2_s1_c_RNIO52I_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_2_s1_c_RNIO52I_LC_15_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_2_s1_c_RNIO52I_LC_15_9_3  (
            .in0(_gnd_net_),
            .in1(N__9114),
            .in2(N__11224),
            .in3(N__8556),
            .lcout(DUT_uart_inst0_rx_countdown_3_s1_3),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_countdown_3_cry_2_s1 ),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_s1_c_RNIQBCS_LC_15_9_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_s1_c_RNIQBCS_LC_15_9_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_s1_c_RNIQBCS_LC_15_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_3_s1_c_RNIQBCS_LC_15_9_4  (
            .in0(_gnd_net_),
            .in1(N__9178),
            .in2(N__11467),
            .in3(N__8553),
            .lcout(DUT_uart_inst0_rx_countdown_3_s1_4),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_countdown_3_cry_3_s1 ),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_4_s1_c_RNISHMM_LC_15_9_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_4_s1_c_RNISHMM_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_4_s1_c_RNISHMM_LC_15_9_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_4_s1_c_RNISHMM_LC_15_9_5  (
            .in0(_gnd_net_),
            .in1(N__11544),
            .in2(_gnd_net_),
            .in3(N__8550),
            .lcout(DUT_uart_inst0_rx_countdown_3_s1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_0_LC_15_9_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_0_LC_15_9_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_0_LC_15_9_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_0_LC_15_9_6  (
            .in0(N__9115),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8536),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15008),
            .ce(),
            .sr(N__8513));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIP8561_0_LC_15_10_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIP8561_0_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIP8561_0_LC_15_10_0 .LUT_INIT=16'b0001111000001111;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNIP8561_0_LC_15_10_0  (
            .in0(N__8678),
            .in1(N__8639),
            .in2(N__8739),
            .in3(N__8786),
            .lcout(\DUT.uart_inst0.m6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_2_LC_15_10_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_2_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_2_LC_15_10_1 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_1_2_LC_15_10_1  (
            .in0(N__9225),
            .in1(N__8729),
            .in2(_gnd_net_),
            .in3(N__8921),
            .lcout(\DUT.uart_inst0.N_19_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_4_2_LC_15_10_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_4_2_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_4_2_LC_15_10_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_4_2_LC_15_10_2  (
            .in0(N__10292),
            .in1(N__10228),
            .in2(N__10169),
            .in3(N__9985),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_2_2_LC_15_10_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_2_2_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_2_2_LC_15_10_3 .LUT_INIT=16'b0000001111110011;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_2_2_LC_15_10_3  (
            .in0(_gnd_net_),
            .in1(N__8730),
            .in2(N__8607),
            .in3(N__8922),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_21_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_2_LC_15_10_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_2_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_2_LC_15_10_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_0_2_LC_15_10_4  (
            .in0(N__10699),
            .in1(_gnd_net_),
            .in2(N__8604),
            .in3(N__8601),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_2_LC_15_10_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_2_LC_15_10_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_bits_remaining_2_LC_15_10_5 .LUT_INIT=16'b1100110001001110;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_2_LC_15_10_5  (
            .in0(N__10814),
            .in1(N__8731),
            .in2(N__8595),
            .in3(N__10314),
            .lcout(\DUT.uart_inst0.rx_bits_remainingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15004),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNI40IN5_1_LC_15_10_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNI40IN5_1_LC_15_10_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNI40IN5_1_LC_15_10_6 .LUT_INIT=16'b1010111111111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNI40IN5_1_LC_15_10_6  (
            .in0(N__9908),
            .in1(N__11392),
            .in2(N__10709),
            .in3(N__10081),
            .lcout(\DUT.uart_inst0.rx_countdown_8_i_o2_2_0_2 ),
            .ltout(\DUT.uart_inst0.rx_countdown_8_i_o2_2_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_1_LC_15_10_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_1_LC_15_10_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_bits_remaining_1_LC_15_10_7 .LUT_INIT=16'b1111011100000010;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_1_LC_15_10_7  (
            .in0(N__10813),
            .in1(N__8592),
            .in2(N__8586),
            .in3(N__8679),
            .lcout(\DUT.uart_inst0.rx_bits_remainingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15004),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_5_LC_15_11_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_5_LC_15_11_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_5_LC_15_11_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \DUT.uart_inst0.recv_state_5_LC_15_11_0  (
            .in0(N__8568),
            .in1(N__8905),
            .in2(N__10823),
            .in3(N__8913),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15002),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_0_LC_15_11_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_0_LC_15_11_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rWritePtr_0_LC_15_11_1 .LUT_INIT=16'b0000000010011001;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_0_LC_15_11_1  (
            .in0(N__12314),
            .in1(N__12243),
            .in2(_gnd_net_),
            .in3(N__8583),
            .lcout(\DUT.fifo_tx_inst.rWritePtrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15002),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_1_LC_15_11_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_1_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_1_LC_15_11_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_1_LC_15_11_2  (
            .in0(N__8867),
            .in1(N__14564),
            .in2(_gnd_net_),
            .in3(N__11035),
            .lcout(\DUT.uart_inst0.g0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_5_LC_15_11_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_5_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_5_LC_15_11_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_5_LC_15_11_3  (
            .in0(N__11332),
            .in1(N__10555),
            .in2(_gnd_net_),
            .in3(N__8868),
            .lcout(\DUT.uart_inst0.N_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNI8OBB2_1_LC_15_11_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNI8OBB2_1_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNI8OBB2_1_LC_15_11_4 .LUT_INIT=16'b0001000100110001;
    LogicCell40 \DUT.uart_inst0.recv_state_RNI8OBB2_1_LC_15_11_4  (
            .in0(N__8866),
            .in1(N__8928),
            .in2(N__10569),
            .in3(N__8800),
            .lcout(\DUT.uart_inst0.N_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNI4AOF7_3_LC_15_11_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNI4AOF7_3_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNI4AOF7_3_LC_15_11_5 .LUT_INIT=16'b0011001111110101;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNI4AOF7_3_LC_15_11_5  (
            .in0(N__9216),
            .in1(N__10302),
            .in2(N__11265),
            .in3(N__10700),
            .lcout(\DUT.uart_inst0.recv_state_srsts_1_5 ),
            .ltout(\DUT.uart_inst0.recv_state_srsts_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_4_LC_15_11_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_4_LC_15_11_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_4_LC_15_11_6 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \DUT.uart_inst0.recv_state_4_LC_15_11_6  (
            .in0(N__10879),
            .in1(N__8906),
            .in2(N__8883),
            .in3(N__8880),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15002),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_4_LC_15_11_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_4_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_4_LC_15_11_7 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_4_LC_15_11_7  (
            .in0(N__14565),
            .in1(N__11175),
            .in2(_gnd_net_),
            .in3(N__10878),
            .lcout(\DUT.uart_inst0.recv_state_srsts_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_3_LC_15_12_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_3_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_3_LC_15_12_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_0_3_LC_15_12_0  (
            .in0(_gnd_net_),
            .in1(N__8693),
            .in2(_gnd_net_),
            .in3(N__8649),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_43_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_3_LC_15_12_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_3_LC_15_12_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_bits_remaining_3_LC_15_12_1 .LUT_INIT=16'b1110111011101011;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_3_LC_15_12_1  (
            .in0(N__8873),
            .in1(N__8709),
            .in2(N__8829),
            .in3(N__8742),
            .lcout(\DUT.uart_inst0.rx_bits_remainingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__14999),
            .ce(N__8825),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIV9PG_3_LC_15_12_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIV9PG_3_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIV9PG_3_LC_15_12_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNIV9PG_3_LC_15_12_2  (
            .in0(_gnd_net_),
            .in1(N__8707),
            .in2(_gnd_net_),
            .in3(N__8647),
            .lcout(),
            .ltout(\DUT.uart_inst0.m3_e_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIAVHE1_2_LC_15_12_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIAVHE1_2_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIAVHE1_2_LC_15_12_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNIAVHE1_2_LC_15_12_3  (
            .in0(N__8692),
            .in1(N__8741),
            .in2(N__8811),
            .in3(N__8801),
            .lcout(\DUT.uart_inst0.N_15_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_4_2_LC_15_12_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_4_2_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_4_2_LC_15_12_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_4_2_LC_15_12_4  (
            .in0(N__8740),
            .in1(N__8708),
            .in2(N__8694),
            .in3(N__8648),
            .lcout(\DUT.uart_inst0.recv_state_RNO_4Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_3_2_LC_15_12_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_3_2_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_3_2_LC_15_12_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_3_2_LC_15_12_5  (
            .in0(N__11490),
            .in1(N__11261),
            .in2(N__11572),
            .in3(N__11139),
            .lcout(\DUT.uart_inst0.N_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNIEQQU_2_LC_15_12_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNIEQQU_2_LC_15_12_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNIEQQU_2_LC_15_12_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNIEQQU_2_LC_15_12_6  (
            .in0(N__11140),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11491),
            .lcout(\DUT.uart_inst0.G_8_i_a3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_3_2_LC_15_12_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_3_2_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_3_2_LC_15_12_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_3_2_LC_15_12_7  (
            .in0(N__11492),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11262),
            .lcout(\DUT.uart_inst0.rx_countdown_8_i_o2_1_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_16_2_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_16_2_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_16_2_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_16_2_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_16_3_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_16_3_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_16_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_16_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12903),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15049),
            .ce(N__11853),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_16_3_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_16_3_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_16_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_16_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13116),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15049),
            .ce(N__11853),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_16_4_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_16_4_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_16_4_0 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_16_4_0  (
            .in0(N__11744),
            .in1(N__11781),
            .in2(N__11678),
            .in3(N__8934),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_16_4_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_16_4_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_16_4_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_16_4_1  (
            .in0(N__12690),
            .in1(N__11865),
            .in2(N__8943),
            .in3(N__11674),
            .lcout(\DUT.rFifoDatarx_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_16_4_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_16_4_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_16_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_16_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12963),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15044),
            .ce(N__11834),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_16_4_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_16_4_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_16_4_3 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_16_4_3  (
            .in0(N__9264),
            .in1(N__11666),
            .in2(N__11073),
            .in3(N__11743),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_16_4_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_16_4_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_16_4_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_16_4_4  (
            .in0(N__11673),
            .in1(N__12474),
            .in2(N__9276),
            .in3(N__11925),
            .lcout(\DUT.rFifoDatarx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_16_4_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_16_4_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_16_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_16_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13011),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15044),
            .ce(N__11834),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_16_4_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_16_4_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_16_4_6 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_16_4_6  (
            .in0(N__11745),
            .in1(N__11064),
            .in2(N__11679),
            .in3(N__9258),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_16_4_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_16_4_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_16_4_7 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_16_4_7  (
            .in0(N__12462),
            .in1(N__11913),
            .in2(N__9252),
            .in3(N__11675),
            .lcout(\DUT.rFifoDatarx_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_16_5_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_16_5_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_16_5_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_16_5_0  (
            .in0(N__9234),
            .in1(N__11657),
            .in2(N__11058),
            .in3(N__11740),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_16_5_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_16_5_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_16_5_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_16_5_1  (
            .in0(N__11662),
            .in1(N__12723),
            .in2(N__9243),
            .in3(N__11886),
            .lcout(\DUT.rFifoDatarx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_16_5_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_16_5_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_16_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_16_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13292),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15038),
            .ce(N__11848),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_16_5_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_16_5_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_16_5_3 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_16_5_3  (
            .in0(N__11739),
            .in1(N__11799),
            .in2(N__11677),
            .in3(N__9537),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_16_5_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_16_5_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_16_5_4 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_16_5_4  (
            .in0(N__12711),
            .in1(N__11880),
            .in2(N__9228),
            .in3(N__11664),
            .lcout(\DUT.rFifoDatarx_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_16_5_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_16_5_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_16_5_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_16_5_5  (
            .in0(N__13058),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15038),
            .ce(N__11848),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_16_5_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_16_5_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_16_5_6 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_16_5_6  (
            .in0(N__9531),
            .in1(N__11658),
            .in2(N__11790),
            .in3(N__11741),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_16_5_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_16_5_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_16_5_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_16_5_7  (
            .in0(N__11663),
            .in1(N__12699),
            .in2(N__9522),
            .in3(N__11874),
            .lcout(\DUT.rFifoDatarx_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIME2J_0_LC_16_6_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIME2J_0_LC_16_6_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIME2J_0_LC_16_6_0 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNIME2J_0_LC_16_6_0  (
            .in0(N__9512),
            .in1(N__9476),
            .in2(N__9412),
            .in3(N__9332),
            .lcout(\DUT.fifo_tx_inst.rReadPtr11 ),
            .ltout(\DUT.fifo_tx_inst.rReadPtr11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rReadPtr_RNILV421_0_LC_16_6_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rReadPtr_RNILV421_0_LC_16_6_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rReadPtr_RNILV421_0_LC_16_6_1 .LUT_INIT=16'b1101010101010101;
    LogicCell40 \DUT.fifo_tx_inst.rReadPtr_RNILV421_0_LC_16_6_1  (
            .in0(N__14556),
            .in1(N__11636),
            .in2(N__9297),
            .in3(N__11728),
            .lcout(\DUT.fifo_tx_inst.un1_i11_2_i ),
            .ltout(\DUT.fifo_tx_inst.un1_i11_2_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rReadPtr_1_LC_16_6_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rReadPtr_1_LC_16_6_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rReadPtr_1_LC_16_6_2 .LUT_INIT=16'b0000011000001010;
    LogicCell40 \DUT.fifo_tx_inst.rReadPtr_1_LC_16_6_2  (
            .in0(N__11637),
            .in1(N__11742),
            .in2(N__9294),
            .in3(N__9291),
            .lcout(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15031),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rReadPtr_0_LC_16_6_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rReadPtr_0_LC_16_6_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rReadPtr_0_LC_16_6_3 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \DUT.fifo_tx_inst.rReadPtr_0_LC_16_6_3  (
            .in0(N__9290),
            .in1(N__9282),
            .in2(_gnd_net_),
            .in3(N__11729),
            .lcout(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15031),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_16_6_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_16_6_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_16_6_4 .LUT_INIT=16'b0010111101111111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_16_6_4  (
            .in0(N__11726),
            .in1(N__11936),
            .in2(N__11665),
            .in3(N__11948),
            .lcout(\DUT.rFifoDataror_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_RNI86BE_LC_16_6_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_RNI86BE_LC_16_6_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_RNI86BE_LC_16_6_5 .LUT_INIT=16'b1100111111011101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_0_RNI86BE_LC_16_6_5  (
            .in0(N__12012),
            .in1(N__11635),
            .in2(N__11964),
            .in3(N__11727),
            .lcout(\DUT.rFifoDataror_1 ),
            .ltout(\DUT.rFifoDataror_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_RNIKCMS_LC_16_6_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_RNIKCMS_LC_16_6_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_RNIKCMS_LC_16_6_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_0_RNIKCMS_LC_16_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9612),
            .in3(N__9605),
            .lcout(\DUT.rFifoDataror_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.rRamWrEn_latch_LC_16_6_7 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.rRamWrEn_latch_LC_16_6_7 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.rRamWrEn_latch_LC_16_6_7 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \fifo_inst.ftdi_input_inst.rRamWrEn_latch_LC_16_6_7  (
            .in0(N__9731),
            .in1(N__15282),
            .in2(N__9765),
            .in3(N__9556),
            .lcout(G_115),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_0_LC_16_7_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_0_LC_16_7_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_0_LC_16_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_0_LC_16_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13569),
            .lcout(\DUT.wRxByte_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15026),
            .ce(N__9783),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_1_LC_16_7_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_1_LC_16_7_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_1_LC_16_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_1_LC_16_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15146),
            .lcout(\DUT.wRxByte_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15026),
            .ce(N__9783),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_2_LC_16_7_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_2_LC_16_7_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_2_LC_16_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_2_LC_16_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13515),
            .lcout(\DUT.wRxByte_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15026),
            .ce(N__9783),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_3_LC_16_7_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_3_LC_16_7_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_3_LC_16_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_3_LC_16_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13467),
            .lcout(\DUT.wRxByte_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15026),
            .ce(N__9783),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_4_LC_16_7_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_4_LC_16_7_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_4_LC_16_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_4_LC_16_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15081),
            .lcout(\DUT.wRxByte_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15026),
            .ce(N__9783),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_5_LC_16_7_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_5_LC_16_7_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_5_LC_16_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_5_LC_16_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13415),
            .lcout(\DUT.wRxByte_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15026),
            .ce(N__9783),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_6_LC_16_7_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_6_LC_16_7_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_6_LC_16_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_6_LC_16_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14066),
            .lcout(\DUT.wRxByte_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15026),
            .ce(N__9783),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_7_LC_16_7_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_7_LC_16_7_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_7_LC_16_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_7_LC_16_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10517),
            .lcout(\DUT.wRxByte_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15026),
            .ce(N__9783),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNIK68E1_1_LC_16_8_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNIK68E1_1_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNIK68E1_1_LC_16_8_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNIK68E1_1_LC_16_8_0  (
            .in0(N__11545),
            .in1(N__11157),
            .in2(_gnd_net_),
            .in3(N__11377),
            .lcout(\DUT.uart_inst0.m6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.un1_rWrState_1_LC_16_8_1 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.un1_rWrState_1_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.un1_rWrState_1_LC_16_8_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \fifo_inst.ftdi_input_inst.un1_rWrState_1_LC_16_8_1  (
            .in0(N__9764),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9735),
            .lcout(\fifo_inst.ftdi_input_inst.un1_rWrStateZ0Z_1 ),
            .ltout(\fifo_inst.ftdi_input_inst.un1_rWrStateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_2_LC_16_8_2 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_2_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_2_LC_16_8_2 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_2_LC_16_8_2  (
            .in0(N__15281),
            .in1(N__9690),
            .in2(N__9714),
            .in3(N__9704),
            .lcout(G_118),
            .ltout(G_118_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.SUM_0_2_LC_16_8_3 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.SUM_0_2_LC_16_8_3 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.SUM_0_2_LC_16_8_3 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \fifo_inst.ftdi_input_inst.SUM_0_2_LC_16_8_3  (
            .in0(N__9640),
            .in1(_gnd_net_),
            .in2(N__9693),
            .in3(N__9676),
            .lcout(G_119),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_0_LC_16_8_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_0_LC_16_8_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_0_LC_16_8_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_0_LC_16_8_4  (
            .in0(N__9839),
            .in1(N__10685),
            .in2(_gnd_net_),
            .in3(N__10071),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15020),
            .ce(N__14456),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_4_LC_16_8_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_4_LC_16_8_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_4_LC_16_8_5 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_4_LC_16_8_5  (
            .in0(N__10684),
            .in1(N__9840),
            .in2(N__11487),
            .in3(N__10289),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15020),
            .ce(N__14456),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_0_LC_16_8_6 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_0_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_0_LC_16_8_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_0_LC_16_8_6  (
            .in0(N__15279),
            .in1(N__9659),
            .in2(_gnd_net_),
            .in3(N__9677),
            .lcout(G_116),
            .ltout(G_116_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_1_LC_16_8_7 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_1_LC_16_8_7 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_1_LC_16_8_7 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_1_LC_16_8_7  (
            .in0(N__9660),
            .in1(N__9641),
            .in2(N__9651),
            .in3(N__15280),
            .lcout(G_117),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_2_1_LC_16_9_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_2_1_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_2_1_LC_16_9_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_2_1_LC_16_9_0  (
            .in0(N__11547),
            .in1(N__11039),
            .in2(N__9807),
            .in3(N__11153),
            .lcout(\DUT.uart_inst0.g1_i_a4_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_4_1_LC_16_9_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_4_1_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_4_1_LC_16_9_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_4_1_LC_16_9_1  (
            .in0(N__10050),
            .in1(N__11256),
            .in2(N__11497),
            .in3(N__11379),
            .lcout(\DUT.uart_inst0.g1_i_a4_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_1_LC_16_9_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_1_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_1_LC_16_9_2 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_0_1_LC_16_9_2  (
            .in0(N__11380),
            .in1(N__10889),
            .in2(N__9920),
            .in3(N__10678),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_78_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_1_LC_16_9_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_1_LC_16_9_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_1_LC_16_9_3 .LUT_INIT=16'b1111010111110000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_1_LC_16_9_3  (
            .in0(N__10424),
            .in1(_gnd_net_),
            .in2(N__9798),
            .in3(N__10952),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15014),
            .ce(N__14461),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNIEQQU_1_LC_16_9_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNIEQQU_1_LC_16_9_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNIEQQU_1_LC_16_9_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNIEQQU_1_LC_16_9_5  (
            .in0(_gnd_net_),
            .in1(N__11546),
            .in2(_gnd_net_),
            .in3(N__11378),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_10_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNI2GC23_0_LC_16_9_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNI2GC23_0_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNI2GC23_0_LC_16_9_6 .LUT_INIT=16'b0011000001110100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNI2GC23_0_LC_16_9_6  (
            .in0(N__9899),
            .in1(N__10051),
            .in2(N__9795),
            .in3(N__10214),
            .lcout(\DUT.uart_inst0.P6_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_5_LC_16_9_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_5_LC_16_9_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_5_LC_16_9_7 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_5_LC_16_9_7  (
            .in0(N__10215),
            .in1(N__9838),
            .in2(N__10706),
            .in3(N__11548),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15014),
            .ce(N__14461),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_3_0_LC_16_10_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_3_0_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_3_0_LC_16_10_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_3_0_LC_16_10_0  (
            .in0(N__10221),
            .in1(N__11174),
            .in2(_gnd_net_),
            .in3(N__9981),
            .lcout(),
            .ltout(\DUT.uart_inst0.G_19_0_a5_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_1_0_LC_16_10_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_1_0_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_1_0_LC_16_10_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_1_0_LC_16_10_1  (
            .in0(N__10153),
            .in1(N__10694),
            .in2(N__9786),
            .in3(N__10274),
            .lcout(),
            .ltout(\DUT.uart_inst0.G_19_0_a5_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_0_LC_16_10_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_0_LC_16_10_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_0_LC_16_10_2 .LUT_INIT=16'b1010101011111110;
    LogicCell40 \DUT.uart_inst0.recv_state_0_LC_16_10_2  (
            .in0(N__10329),
            .in1(N__9846),
            .in2(N__10317),
            .in3(N__10313),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15009),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rReadPtr_0_LC_16_10_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rReadPtr_0_LC_16_10_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rReadPtr_0_LC_16_10_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \DUT.fifo_rx_inst.rReadPtr_0_LC_16_10_3  (
            .in0(N__11048),
            .in1(N__13817),
            .in2(_gnd_net_),
            .in3(N__12573),
            .lcout(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15009),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNI8H662_LC_16_10_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNI8H662_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNI8H662_LC_16_10_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNI8H662_LC_16_10_4  (
            .in0(N__10272),
            .in1(N__9977),
            .in2(_gnd_net_),
            .in3(N__10151),
            .lcout(\DUT.uart_inst0.G_8_i_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_2_3_LC_16_10_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_2_3_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_2_3_LC_16_10_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_2_3_LC_16_10_5  (
            .in0(_gnd_net_),
            .in1(N__10273),
            .in2(_gnd_net_),
            .in3(N__10220),
            .lcout(\DUT.uart_inst0.m10_e_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rReadPtr_1_LC_16_10_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rReadPtr_1_LC_16_10_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rReadPtr_1_LC_16_10_6 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \DUT.fifo_rx_inst.rReadPtr_1_LC_16_10_6  (
            .in0(N__12572),
            .in1(N__13733),
            .in2(N__13821),
            .in3(N__11049),
            .lcout(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15009),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_3_3_LC_16_10_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_3_3_LC_16_10_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_3_3_LC_16_10_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_3_3_LC_16_10_7  (
            .in0(N__10152),
            .in1(N__10080),
            .in2(N__9996),
            .in3(N__9907),
            .lcout(\DUT.uart_inst0.m10_e_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_2_0_LC_16_11_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_2_0_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_2_0_LC_16_11_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_2_0_LC_16_11_0  (
            .in0(N__10692),
            .in1(N__11564),
            .in2(N__11085),
            .in3(N__11480),
            .lcout(\DUT.uart_inst0.G_19_0_a5_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNIHH651_5_LC_16_11_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNIHH651_5_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNIHH651_5_LC_16_11_1 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \DUT.uart_inst0.recv_state_RNIHH651_5_LC_16_11_1  (
            .in0(N__10927),
            .in1(N__10877),
            .in2(_gnd_net_),
            .in3(N__10565),
            .lcout(\DUT.uart_inst0.N_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_1_1_LC_16_11_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_1_1_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_1_1_LC_16_11_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_1_1_LC_16_11_2  (
            .in0(N__12301),
            .in1(N__12272),
            .in2(_gnd_net_),
            .in3(N__12241),
            .lcout(\DUT.fifo_tx_inst.rFifoData_awe0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rReadPtr_RNI4NC92_0_LC_16_11_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rReadPtr_RNI4NC92_0_LC_16_11_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rReadPtr_RNI4NC92_0_LC_16_11_3 .LUT_INIT=16'b1000000011111111;
    LogicCell40 \DUT.fifo_rx_inst.rReadPtr_RNI4NC92_0_LC_16_11_3  (
            .in0(N__13736),
            .in1(N__13813),
            .in2(N__12566),
            .in3(N__14566),
            .lcout(\DUT.fifo_rx_inst.N_77_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNI237O_0_LC_16_11_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNI237O_0_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNI237O_0_LC_16_11_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNI237O_0_LC_16_11_4  (
            .in0(N__10564),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10925),
            .lcout(\DUT.uart_inst0.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_4_2_LC_16_11_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_4_2_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_4_2_LC_16_11_5 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_4_2_LC_16_11_5  (
            .in0(N__10926),
            .in1(N__10876),
            .in2(_gnd_net_),
            .in3(N__10566),
            .lcout(\DUT.uart_inst0.rx_countdown_8_i_a2_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_3_LC_16_11_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_3_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_3_LC_16_11_6 .LUT_INIT=16'b0010011100001111;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_3_LC_16_11_6  (
            .in0(N__10836),
            .in1(N__11285),
            .in2(N__11336),
            .in3(N__10830),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_20_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_3_LC_16_11_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_3_LC_16_11_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_3_LC_16_11_7 .LUT_INIT=16'b0000110001000100;
    LogicCell40 \DUT.uart_inst0.recv_state_3_LC_16_11_7  (
            .in0(N__11271),
            .in1(N__10821),
            .in2(N__10713),
            .in3(N__10693),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15005),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_4_6_LC_16_12_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_4_6_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_4_6_LC_16_12_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_4_6_LC_16_12_0  (
            .in0(N__11321),
            .in1(N__11493),
            .in2(N__10338),
            .in3(N__11264),
            .lcout(),
            .ltout(\DUT.uart_inst0.m7_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_1_6_LC_16_12_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_1_6_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_1_6_LC_16_12_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_1_6_LC_16_12_1  (
            .in0(N__11562),
            .in1(N__11155),
            .in2(N__10581),
            .in3(N__11397),
            .lcout(\DUT.uart_inst0.N_28_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_5_6_LC_16_12_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_5_6_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_5_6_LC_16_12_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_5_6_LC_16_12_3  (
            .in0(N__10556),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14572),
            .lcout(\DUT.uart_inst0.m2_e_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.oRxFlag_RNIHCKH1_LC_16_12_4 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.oRxFlag_RNIHCKH1_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_output_inst.oRxFlag_RNIHCKH1_LC_16_12_4 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \fifo_inst.ftdi_output_inst.oRxFlag_RNIHCKH1_LC_16_12_4  (
            .in0(N__15278),
            .in1(N__14812),
            .in2(_gnd_net_),
            .in3(N__12539),
            .lcout(rTxByte_1_sqmuxa_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_5_3_LC_16_12_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_5_3_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_5_3_LC_16_12_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_5_3_LC_16_12_5  (
            .in0(N__11563),
            .in1(N__11257),
            .in2(N__11499),
            .in3(N__11398),
            .lcout(),
            .ltout(\DUT.uart_inst0.m6_e_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_1_3_LC_16_12_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_1_3_LC_16_12_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_1_3_LC_16_12_6 .LUT_INIT=16'b0001010111010101;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_1_3_LC_16_12_6  (
            .in0(N__11322),
            .in1(N__11301),
            .in2(N__11289),
            .in3(N__11286),
            .lcout(\DUT.uart_inst0.N_18_mux_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_4_0_LC_16_12_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_4_0_LC_16_12_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_4_0_LC_16_12_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_4_0_LC_16_12_7  (
            .in0(N__11263),
            .in1(N__11173),
            .in2(_gnd_net_),
            .in3(N__11154),
            .lcout(\DUT.uart_inst0.G_19_0_a5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_17_4_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_17_4_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_17_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_17_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13007),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15050),
            .ce(N__11997),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_17_4_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_17_4_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_17_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_17_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12902),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15050),
            .ce(N__11997),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_17_4_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_17_4_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_17_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_17_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12843),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15050),
            .ce(N__11997),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_17_4_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_17_4_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_17_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_17_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13371),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15050),
            .ce(N__11997),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_17_4_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_17_4_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_17_4_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_17_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13293),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15050),
            .ce(N__11997),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_17_4_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_17_4_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_17_4_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_17_4_5  (
            .in0(N__13059),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15050),
            .ce(N__11997),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_17_4_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_17_4_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_17_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_17_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13115),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15050),
            .ce(N__11997),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_17_4_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_17_4_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_17_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_17_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12959),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15050),
            .ce(N__11997),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_17_5_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_17_5_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_17_5_0 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_17_5_0  (
            .in0(N__11751),
            .in1(N__11654),
            .in2(N__11775),
            .in3(N__11731),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_17_5_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_17_5_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_17_5_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_17_5_1  (
            .in0(N__11656),
            .in1(N__12738),
            .in2(N__11763),
            .in3(N__11901),
            .lcout(\DUT.rFifoDatarx_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_17_5_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_17_5_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_17_5_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_17_5_2  (
            .in0(N__12839),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15045),
            .ce(N__11852),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_17_5_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_17_5_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_17_5_3 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_17_5_3  (
            .in0(N__11730),
            .in1(N__11688),
            .in2(N__11676),
            .in3(N__11580),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_17_5_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_17_5_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_17_5_4 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_17_5_4  (
            .in0(N__12732),
            .in1(N__11892),
            .in2(N__11682),
            .in3(N__11655),
            .lcout(\DUT.rFifoDatarx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_17_5_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_17_5_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_17_5_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_17_5_5  (
            .in0(N__13367),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15045),
            .ce(N__11852),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_17_6_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_17_6_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_17_6_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_17_6_0  (
            .in0(N__13000),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15039),
            .ce(N__12207),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_17_6_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_17_6_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_17_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_17_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12895),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15039),
            .ce(N__12207),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_17_6_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_17_6_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_17_6_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_17_6_2  (
            .in0(_gnd_net_),
            .in1(N__12838),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15039),
            .ce(N__12207),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_17_6_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_17_6_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_17_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_17_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13366),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15039),
            .ce(N__12207),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_17_6_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_17_6_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_17_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_17_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13285),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15039),
            .ce(N__12207),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_17_6_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_17_6_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_17_6_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_17_6_5  (
            .in0(N__13051),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15039),
            .ce(N__12207),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_17_6_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_17_6_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_17_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_17_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13108),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15039),
            .ce(N__12207),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_17_6_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_17_6_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_17_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_17_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12958),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15039),
            .ce(N__12207),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_3_LC_17_7_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_3_LC_17_7_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_3_LC_17_7_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_3_LC_17_7_0  (
            .in0(_gnd_net_),
            .in1(N__12083),
            .in2(_gnd_net_),
            .in3(N__12026),
            .lcout(\DUT.fifo_rx_inst.rFifoDataro_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15032),
            .ce(),
            .sr(N__15231));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_LC_17_7_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_LC_17_7_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_LC_17_7_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_0_LC_17_7_1  (
            .in0(_gnd_net_),
            .in1(N__12011),
            .in2(_gnd_net_),
            .in3(N__11838),
            .lcout(\DUT.fifo_tx_inst.rFifoDataro_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15032),
            .ce(),
            .sr(N__15231));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_1_LC_17_7_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_1_LC_17_7_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_1_LC_17_7_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_1_LC_17_7_2  (
            .in0(_gnd_net_),
            .in1(N__11963),
            .in2(_gnd_net_),
            .in3(N__11993),
            .lcout(\DUT.fifo_tx_inst.rFifoDataro_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15032),
            .ce(),
            .sr(N__15231));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_LC_17_7_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_LC_17_7_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_LC_17_7_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_2_LC_17_7_3  (
            .in0(_gnd_net_),
            .in1(N__12203),
            .in2(_gnd_net_),
            .in3(N__11949),
            .lcout(\DUT.fifo_tx_inst.rFifoDataro_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15032),
            .ce(),
            .sr(N__15231));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_3_LC_17_7_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_3_LC_17_7_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_3_LC_17_7_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_3_LC_17_7_4  (
            .in0(_gnd_net_),
            .in1(N__11937),
            .in2(_gnd_net_),
            .in3(N__12671),
            .lcout(\DUT.fifo_tx_inst.rFifoDataro_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15032),
            .ce(),
            .sr(N__15231));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_17_8_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_17_8_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_17_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_17_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13612),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15027),
            .ce(N__12084),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_17_8_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_17_8_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_17_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_17_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13570),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15027),
            .ce(N__12084),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_17_8_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_17_8_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_17_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_17_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15147),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15027),
            .ce(N__12084),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_17_8_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_17_8_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_17_8_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_17_8_3  (
            .in0(N__13516),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15027),
            .ce(N__12084),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_17_8_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_17_8_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_17_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_17_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13468),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15027),
            .ce(N__12084),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_17_8_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_17_8_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_17_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_17_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15082),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15027),
            .ce(N__12084),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_17_8_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_17_8_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_17_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_17_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13416),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15027),
            .ce(N__12084),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_17_8_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_17_8_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_17_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_17_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14067),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15027),
            .ce(N__12084),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_17_9_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_17_9_0 .LUT_INIT=16'b0100011001010111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_17_9_0  (
            .in0(N__13808),
            .in1(N__13700),
            .in2(N__14100),
            .in3(N__12048),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIT6K22_6_LC_17_9_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIT6K22_6_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIT6K22_6_LC_17_9_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIT6K22_6_LC_17_9_1  (
            .in0(N__12057),
            .in1(N__13155),
            .in2(N__12051),
            .in3(N__13709),
            .lcout(\DUT.fifo_rx_inst.rFifoDatarx_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_17_9_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_17_9_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_17_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_17_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13426),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15021),
            .ce(N__14859),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_17_9_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_17_9_3 .LUT_INIT=16'b0000010111110011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_17_9_3  (
            .in0(N__14040),
            .in1(N__12033),
            .in2(N__13734),
            .in3(N__13809),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI1BK22_7_LC_17_9_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI1BK22_7_LC_17_9_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI1BK22_7_LC_17_9_4 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI1BK22_7_LC_17_9_4  (
            .in0(N__12042),
            .in1(N__13149),
            .in2(N__12036),
            .in3(N__13704),
            .lcout(\DUT.fifo_rx_inst.rFifoDatarx_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_17_9_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_17_9_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_17_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_17_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14086),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15021),
            .ce(N__14859),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_17_9_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_17_9_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_17_9_6 .LUT_INIT=16'b0010010101110101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_17_9_6  (
            .in0(N__13807),
            .in1(N__12027),
            .in2(N__13735),
            .in3(N__12417),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoDataror_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNI5NR43_LC_17_9_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNI5NR43_LC_17_9_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNI5NR43_LC_17_9_7 .LUT_INIT=16'b1111000000110101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_0_RNI5NR43_LC_17_9_7  (
            .in0(N__12434),
            .in1(N__12450),
            .in2(N__12138),
            .in3(N__13708),
            .lcout(\DUT.fifo_rx_inst.rFifoDataror_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_17_10_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_17_10_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_17_10_0 .LUT_INIT=16'b0000010111110011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_17_10_0  (
            .in0(N__13494),
            .in1(N__12123),
            .in2(N__13739),
            .in3(N__13810),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIHQJ22_3_LC_17_10_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIHQJ22_3_LC_17_10_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIHQJ22_3_LC_17_10_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIHQJ22_3_LC_17_10_1  (
            .in0(N__12135),
            .in1(N__12759),
            .in2(N__12126),
            .in3(N__13731),
            .lcout(\DUT.fifo_rx_inst.rFifoDatarx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_17_10_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_17_10_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_17_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_17_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13536),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15015),
            .ce(N__14866),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_17_10_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_17_10_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_17_10_3 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_17_10_3  (
            .in0(N__13811),
            .in1(N__13446),
            .in2(N__12105),
            .in3(N__13729),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNILUJ22_4_LC_17_10_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNILUJ22_4_LC_17_10_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNILUJ22_4_LC_17_10_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNILUJ22_4_LC_17_10_4  (
            .in0(N__13730),
            .in1(N__12117),
            .in2(N__12108),
            .in3(N__12747),
            .lcout(\DUT.fifo_rx_inst.rFifoDatarx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_17_10_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_17_10_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_17_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_17_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13480),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15015),
            .ce(N__14866),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_17_10_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_17_10_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_17_10_6 .LUT_INIT=16'b0000010111110011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_17_10_6  (
            .in0(N__13440),
            .in1(N__15063),
            .in2(N__13740),
            .in3(N__13812),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIP2K22_5_LC_17_10_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIP2K22_5_LC_17_10_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIP2K22_5_LC_17_10_7 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIP2K22_5_LC_17_10_7  (
            .in0(N__12096),
            .in1(N__13167),
            .in2(N__12087),
            .in3(N__13732),
            .lcout(\DUT.fifo_rx_inst.rFifoDatarx_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_LC_17_11_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_LC_17_11_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_LC_17_11_0 .LUT_INIT=16'b1100110111001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_0_LC_17_11_0  (
            .in0(N__12349),
            .in1(N__12449),
            .in2(N__12401),
            .in3(N__12167),
            .lcout(\DUT.fifo_rx_inst.rFifoDataro_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15010),
            .ce(),
            .sr(N__15224));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_1_LC_17_11_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_1_LC_17_11_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_1_LC_17_11_1 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_1_LC_17_11_1  (
            .in0(N__12168),
            .in1(N__12396),
            .in2(N__12435),
            .in3(N__12350),
            .lcout(\DUT.fifo_rx_inst.rFifoDataro_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15010),
            .ce(),
            .sr(N__15224));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_LC_17_11_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_LC_17_11_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_LC_17_11_2 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_2_LC_17_11_2  (
            .in0(N__12351),
            .in1(N__12169),
            .in2(N__12402),
            .in3(N__12416),
            .lcout(\DUT.fifo_rx_inst.rFifoDataro_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15010),
            .ce(),
            .sr(N__15224));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_17_11_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_17_11_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_17_11_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_17_11_3  (
            .in0(N__12164),
            .in1(N__12388),
            .in2(_gnd_net_),
            .in3(N__12346),
            .lcout(\DUT.fifo_rx_inst.rFifoData_awe1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_17_11_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_17_11_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_17_11_4 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_17_11_4  (
            .in0(N__12348),
            .in1(_gnd_net_),
            .in2(N__12400),
            .in3(N__12166),
            .lcout(\DUT.fifo_rx_inst.rFifoData_awe2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_17_11_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_17_11_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_17_11_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_17_11_5  (
            .in0(N__12165),
            .in1(N__12389),
            .in2(_gnd_net_),
            .in3(N__12347),
            .lcout(\DUT.fifo_rx_inst.rFifoData_awe0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_1_LC_17_11_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_1_LC_17_11_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_1_LC_17_11_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_1_LC_17_11_7  (
            .in0(N__12313),
            .in1(N__12276),
            .in2(_gnd_net_),
            .in3(N__12242),
            .lcout(\DUT.fifo_tx_inst.rFifoData_awe2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_17_12_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_17_12_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_17_12_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_17_12_0  (
            .in0(_gnd_net_),
            .in1(N__12604),
            .in2(_gnd_net_),
            .in3(N__13895),
            .lcout(\DUT.fifo_rx_inst.rWritePtr16 ),
            .ltout(\DUT.fifo_rx_inst.rWritePtr16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_17_12_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_17_12_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_17_12_1 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_17_12_1  (
            .in0(N__13925),
            .in1(N__14011),
            .in2(N__12186),
            .in3(N__13947),
            .lcout(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_0_LC_17_12_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_0_LC_17_12_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoCount_0_LC_17_12_2 .LUT_INIT=16'b0101101000111100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_0_LC_17_12_2  (
            .in0(N__13949),
            .in1(N__12170),
            .in2(N__14015),
            .in3(N__13928),
            .lcout(\DUT.fifo_rx_inst.rFifoCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15006),
            .ce(),
            .sr(N__15223));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI110Q1_1_LC_17_12_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI110Q1_1_LC_17_12_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI110Q1_1_LC_17_12_3 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNI110Q1_1_LC_17_12_3  (
            .in0(N__13894),
            .in1(N__13968),
            .in2(N__12609),
            .in3(N__14005),
            .lcout(\DUT.fifo_rx_inst.N_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI9EGD1_1_LC_17_12_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI9EGD1_1_LC_17_12_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI9EGD1_1_LC_17_12_4 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNI9EGD1_1_LC_17_12_4  (
            .in0(N__14006),
            .in1(N__13924),
            .in2(N__13976),
            .in3(N__13896),
            .lcout(\DUT.fifo_rx_inst.N_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIPTFQ1_1_LC_17_12_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIPTFQ1_1_LC_17_12_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIPTFQ1_1_LC_17_12_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNIPTFQ1_1_LC_17_12_5  (
            .in0(N__13926),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13948),
            .lcout(\DUT.fifo_rx_inst.rFifoCount_RNIPTFQ1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_1_LC_17_12_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_1_LC_17_12_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_1_LC_17_12_6 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_1_LC_17_12_6  (
            .in0(N__14007),
            .in1(_gnd_net_),
            .in2(N__13977),
            .in3(N__13897),
            .lcout(N_69_mux),
            .ltout(N_69_mux_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rRxRead_LC_17_12_7.C_ON=1'b0;
    defparam rRxRead_LC_17_12_7.SEQ_MODE=4'b1000;
    defparam rRxRead_LC_17_12_7.LUT_INIT=16'b1010101000001111;
    LogicCell40 rRxRead_LC_17_12_7 (
            .in0(N__13927),
            .in1(_gnd_net_),
            .in2(N__12528),
            .in3(N__14813),
            .lcout(rRxReadZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15006),
            .ce(),
            .sr(N__15223));
    defparam ioFifoData_iobuf_RNO_1_LC_18_1_4.C_ON=1'b0;
    defparam ioFifoData_iobuf_RNO_1_LC_18_1_4.SEQ_MODE=4'b0000;
    defparam ioFifoData_iobuf_RNO_1_LC_18_1_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 ioFifoData_iobuf_RNO_1_LC_18_1_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13851),
            .lcout(N_1258_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.oTx_n_RNIPDL9_LC_18_3_2 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.oTx_n_RNIPDL9_LC_18_3_2 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_output_inst.oTx_n_RNIPDL9_LC_18_3_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \fifo_inst.ftdi_output_inst.oTx_n_RNIPDL9_LC_18_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14215),
            .lcout(P1A4_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_18_5_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_18_5_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_18_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_18_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12999),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15051),
            .ce(N__12678),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_18_5_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_18_5_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_18_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_18_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12894),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15051),
            .ce(N__12678),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_18_5_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_18_5_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_18_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_18_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12837),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15051),
            .ce(N__12678),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_18_5_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_18_5_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_18_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_18_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13365),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15051),
            .ce(N__12678),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_18_5_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_18_5_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_18_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_18_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13275),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15051),
            .ce(N__12678),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_18_5_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_18_5_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_18_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_18_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13050),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15051),
            .ce(N__12678),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_18_5_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_18_5_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_18_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_18_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13104),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15051),
            .ce(N__12678),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_18_5_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_18_5_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_18_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_18_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12948),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15051),
            .ce(N__12678),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_3_LC_18_6_4 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_3_LC_18_6_4 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_3_LC_18_6_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \fifo_inst.ftdi_output_inst.rRxData_esr_3_LC_18_6_4  (
            .in0(N__12648),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(wRxFifoData_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15046),
            .ce(N__14267),
            .sr(N__15240));
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_1_LC_18_7_1 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_1_LC_18_7_1 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_1_LC_18_7_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \fifo_inst.ftdi_output_inst.rRxData_esr_1_LC_18_7_1  (
            .in0(N__12633),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(wRxFifoData_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15040),
            .ce(N__14268),
            .sr(N__15236));
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_5_LC_18_7_2 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_5_LC_18_7_2 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_5_LC_18_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rRxData_esr_5_LC_18_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12618),
            .lcout(wRxFifoData_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15040),
            .ce(N__14268),
            .sr(N__15236));
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_2_LC_18_7_3 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_2_LC_18_7_3 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_2_LC_18_7_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \fifo_inst.ftdi_output_inst.rRxData_esr_2_LC_18_7_3  (
            .in0(N__12810),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(wRxFifoData_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15040),
            .ce(N__14268),
            .sr(N__15236));
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_0_LC_18_7_4 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_0_LC_18_7_4 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_0_LC_18_7_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \fifo_inst.ftdi_output_inst.rRxData_esr_0_LC_18_7_4  (
            .in0(N__12798),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(wRxFifoData_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15040),
            .ce(N__14268),
            .sr(N__15236));
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_6_LC_18_7_6 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_6_LC_18_7_6 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_6_LC_18_7_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \fifo_inst.ftdi_output_inst.rRxData_esr_6_LC_18_7_6  (
            .in0(_gnd_net_),
            .in1(N__12786),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(wRxFifoData_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15040),
            .ce(N__14268),
            .sr(N__15236));
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_4_LC_18_7_7 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_4_LC_18_7_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_4_LC_18_7_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \fifo_inst.ftdi_output_inst.rRxData_esr_4_LC_18_7_7  (
            .in0(N__12771),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(wRxFifoData_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15040),
            .ce(N__14268),
            .sr(N__15236));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_18_8_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_18_8_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_18_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_18_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13630),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15033),
            .ce(N__13143),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_18_8_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_18_8_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_18_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_18_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13588),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15033),
            .ce(N__13143),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_18_8_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_18_8_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_18_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_18_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15166),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15033),
            .ce(N__13143),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_18_8_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_18_8_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_18_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_18_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13534),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15033),
            .ce(N__13143),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_18_8_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_18_8_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_18_8_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_18_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13487),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15033),
            .ce(N__13143),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_18_8_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_18_8_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_18_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_18_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15106),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15033),
            .ce(N__13143),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_18_8_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_18_8_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_18_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_18_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13433),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15033),
            .ce(N__13143),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_18_8_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_18_8_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_18_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_18_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14087),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15033),
            .ce(N__13143),
            .sr(_gnd_net_));
    defparam rTxByte_esr_6_LC_18_9_0.C_ON=1'b0;
    defparam rTxByte_esr_6_LC_18_9_0.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_6_LC_18_9_0.LUT_INIT=16'b1100000011001010;
    LogicCell40 rTxByte_esr_6_LC_18_9_0 (
            .in0(N__13131),
            .in1(N__13125),
            .in2(N__14826),
            .in3(N__13337),
            .lcout(rTxByteZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15028),
            .ce(N__13257),
            .sr(N__15230));
    defparam rTxByte_esr_5_LC_18_9_1.C_ON=1'b0;
    defparam rTxByte_esr_5_LC_18_9_1.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_5_LC_18_9_1.LUT_INIT=16'b1101000111000000;
    LogicCell40 rTxByte_esr_5_LC_18_9_1 (
            .in0(N__13336),
            .in1(N__14819),
            .in2(N__13077),
            .in3(N__13065),
            .lcout(rTxByteZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15028),
            .ce(N__13257),
            .sr(N__15230));
    defparam rTxByte_esr_0_LC_18_9_2.C_ON=1'b0;
    defparam rTxByte_esr_0_LC_18_9_2.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_0_LC_18_9_2.LUT_INIT=16'b1010000011100100;
    LogicCell40 rTxByte_esr_0_LC_18_9_2 (
            .in0(N__14814),
            .in1(N__13221),
            .in2(N__13023),
            .in3(N__13331),
            .lcout(rTxByteZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15028),
            .ce(N__13257),
            .sr(N__15230));
    defparam rTxByte_esr_7_LC_18_9_3.C_ON=1'b0;
    defparam rTxByte_esr_7_LC_18_9_3.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_7_LC_18_9_3.LUT_INIT=16'b1101000111000000;
    LogicCell40 rTxByte_esr_7_LC_18_9_3 (
            .in0(N__13338),
            .in1(N__14823),
            .in2(N__14286),
            .in3(N__12969),
            .lcout(rTxByteZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15028),
            .ce(N__13257),
            .sr(N__15230));
    defparam rTxByte_esr_1_LC_18_9_4.C_ON=1'b0;
    defparam rTxByte_esr_1_LC_18_9_4.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_1_LC_18_9_4.LUT_INIT=16'b1010000011100100;
    LogicCell40 rTxByte_esr_1_LC_18_9_4 (
            .in0(N__14815),
            .in1(N__13185),
            .in2(N__12915),
            .in3(N__13332),
            .lcout(rTxByteZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15028),
            .ce(N__13257),
            .sr(N__15230));
    defparam rTxByte_esr_2_LC_18_9_5.C_ON=1'b0;
    defparam rTxByte_esr_2_LC_18_9_5.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_2_LC_18_9_5.LUT_INIT=16'b1101000111000000;
    LogicCell40 rTxByte_esr_2_LC_18_9_5 (
            .in0(N__13333),
            .in1(N__14816),
            .in2(N__12855),
            .in3(N__13638),
            .lcout(rTxByteZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15028),
            .ce(N__13257),
            .sr(N__15230));
    defparam rTxByte_esr_3_LC_18_9_6.C_ON=1'b0;
    defparam rTxByte_esr_3_LC_18_9_6.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_3_LC_18_9_6.LUT_INIT=16'b1010000011100100;
    LogicCell40 rTxByte_esr_3_LC_18_9_6 (
            .in0(N__14817),
            .in1(N__13389),
            .in2(N__13383),
            .in3(N__13334),
            .lcout(rTxByteZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15028),
            .ce(N__13257),
            .sr(N__15230));
    defparam rTxByte_esr_4_LC_18_9_7.C_ON=1'b0;
    defparam rTxByte_esr_4_LC_18_9_7.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_4_LC_18_9_7.LUT_INIT=16'b1101000111000000;
    LogicCell40 rTxByte_esr_4_LC_18_9_7 (
            .in0(N__13335),
            .in1(N__14818),
            .in2(N__13311),
            .in3(N__13299),
            .lcout(rTxByteZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15028),
            .ce(N__13257),
            .sr(N__15230));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_18_10_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_18_10_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_18_10_0 .LUT_INIT=16'b0000010111110011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_18_10_0  (
            .in0(N__13596),
            .in1(N__13215),
            .in2(N__13737),
            .in3(N__13815),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI5EJ22_0_LC_18_10_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI5EJ22_0_LC_18_10_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI5EJ22_0_LC_18_10_1 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI5EJ22_0_LC_18_10_1  (
            .in0(N__13245),
            .in1(N__13236),
            .in2(N__13224),
            .in3(N__13721),
            .lcout(\DUT.fifo_rx_inst.rFifoDatarx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_18_10_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_18_10_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_18_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_18_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13631),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15022),
            .ce(N__14867),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_18_10_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_18_10_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_18_10_3 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_18_10_3  (
            .in0(N__13814),
            .in1(N__13548),
            .in2(N__13179),
            .in3(N__13716),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI9IJ22_1_LC_18_10_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI9IJ22_1_LC_18_10_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI9IJ22_1_LC_18_10_4 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI9IJ22_1_LC_18_10_4  (
            .in0(N__13720),
            .in1(N__13209),
            .in2(N__13197),
            .in3(N__13194),
            .lcout(\DUT.fifo_rx_inst.rFifoDatarx_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_18_10_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_18_10_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_18_10_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_18_10_5  (
            .in0(N__13589),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15022),
            .ce(N__14867),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_18_10_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_18_10_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_18_10_6 .LUT_INIT=16'b0000010111110011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_18_10_6  (
            .in0(N__13542),
            .in1(N__15120),
            .in2(N__13738),
            .in3(N__13816),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIDMJ22_2_LC_18_10_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIDMJ22_2_LC_18_10_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIDMJ22_2_LC_18_10_7 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIDMJ22_2_LC_18_10_7  (
            .in0(N__13764),
            .in1(N__13752),
            .in2(N__13743),
            .in3(N__13722),
            .lcout(\DUT.fifo_rx_inst.rFifoDatarx_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_18_11_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_18_11_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_18_11_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_18_11_0  (
            .in0(N__13632),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15016),
            .ce(N__14028),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_18_11_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_18_11_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_18_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_18_11_1  (
            .in0(N__13590),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15016),
            .ce(N__14028),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_18_11_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_18_11_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_18_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_18_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15167),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15016),
            .ce(N__14028),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_18_11_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_18_11_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_18_11_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_18_11_3  (
            .in0(N__13535),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15016),
            .ce(N__14028),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_18_11_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_18_11_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_18_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_18_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13488),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15016),
            .ce(N__14028),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_18_11_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_18_11_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_18_11_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_18_11_5  (
            .in0(N__15111),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15016),
            .ce(N__14028),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_18_11_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_18_11_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_18_11_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_18_11_6  (
            .in0(_gnd_net_),
            .in1(N__13434),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15016),
            .ce(N__14028),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_18_11_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_18_11_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_18_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_18_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14088),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15016),
            .ce(N__14028),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_LC_18_12_0 .C_ON=1'b1;
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_LC_18_12_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_LC_18_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_LC_18_12_0  (
            .in0(_gnd_net_),
            .in1(N__14022),
            .in2(N__14016),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_12_0_),
            .carryout(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_1_LC_18_12_1 .C_ON=1'b1;
    defparam \DUT.fifo_rx_inst.rFifoCount_1_LC_18_12_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoCount_1_LC_18_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_1_LC_18_12_1  (
            .in0(_gnd_net_),
            .in1(N__13975),
            .in2(N__13986),
            .in3(N__13953),
            .lcout(\DUT.fifo_rx_inst.rFifoCountZ0Z_1 ),
            .ltout(),
            .carryin(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0 ),
            .carryout(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1 ),
            .clk(N__15011),
            .ce(),
            .sr(N__15225));
    defparam \DUT.fifo_rx_inst.rFifoCount_2_LC_18_12_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_2_LC_18_12_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoCount_2_LC_18_12_2 .LUT_INIT=16'b1001010101101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_2_LC_18_12_2  (
            .in0(N__13901),
            .in1(N__13950),
            .in2(N__13932),
            .in3(N__13905),
            .lcout(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15011),
            .ce(),
            .sr(N__15225));
    defparam ioFifoData_iobuf_RNO_4_LC_20_3_6.C_ON=1'b0;
    defparam ioFifoData_iobuf_RNO_4_LC_20_3_6.SEQ_MODE=4'b0000;
    defparam ioFifoData_iobuf_RNO_4_LC_20_3_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 ioFifoData_iobuf_RNO_4_LC_20_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13860),
            .lcout(N_1261_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.oTx_n_rep4_ess_LC_20_6_1 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.oTx_n_rep4_ess_LC_20_6_1 .SEQ_MODE=4'b1001;
    defparam \fifo_inst.ftdi_output_inst.oTx_n_rep4_ess_LC_20_6_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \fifo_inst.ftdi_output_inst.oTx_n_rep4_ess_LC_20_6_1  (
            .in0(N__15358),
            .in1(_gnd_net_),
            .in2(N__15422),
            .in3(_gnd_net_),
            .lcout(oTx_n_rep4_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15053),
            .ce(N__15302),
            .sr(N__15248));
    defparam \fifo_inst.ftdi_output_inst.oTx_n_rep1_ess_LC_20_6_3 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.oTx_n_rep1_ess_LC_20_6_3 .SEQ_MODE=4'b1001;
    defparam \fifo_inst.ftdi_output_inst.oTx_n_rep1_ess_LC_20_6_3 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \fifo_inst.ftdi_output_inst.oTx_n_rep1_ess_LC_20_6_3  (
            .in0(N__15357),
            .in1(_gnd_net_),
            .in2(N__15421),
            .in3(_gnd_net_),
            .lcout(oTx_n_rep1_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15053),
            .ce(N__15302),
            .sr(N__15248));
    defparam \fifo_inst.ftdi_output_inst.oTx_n_rep0_ess_LC_20_6_4 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.oTx_n_rep0_ess_LC_20_6_4 .SEQ_MODE=4'b1001;
    defparam \fifo_inst.ftdi_output_inst.oTx_n_rep0_ess_LC_20_6_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.oTx_n_rep0_ess_LC_20_6_4  (
            .in0(_gnd_net_),
            .in1(N__15410),
            .in2(_gnd_net_),
            .in3(N__15356),
            .lcout(oTx_n_rep0_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15053),
            .ce(N__15302),
            .sr(N__15248));
    defparam \fifo_inst.ftdi_output_inst.oRamRdAddr_0_LC_20_7_0 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.oRamRdAddr_0_LC_20_7_0 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.oRamRdAddr_0_LC_20_7_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.oRamRdAddr_0_LC_20_7_0  (
            .in0(N__15341),
            .in1(N__14567),
            .in2(N__15408),
            .in3(N__14172),
            .lcout(\fifo_inst.wRamRdAddr_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15052),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIFFVH_4_LC_20_7_1 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIFFVH_4_LC_20_7_1 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIFFVH_4_LC_20_7_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_RNIFFVH_4_LC_20_7_1  (
            .in0(_gnd_net_),
            .in1(N__15387),
            .in2(_gnd_net_),
            .in3(N__15339),
            .lcout(\fifo_inst.ftdi_output_inst.N_77_0 ),
            .ltout(\fifo_inst.ftdi_output_inst.N_77_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIUEQM_3_LC_20_7_2 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIUEQM_3_LC_20_7_2 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIUEQM_3_LC_20_7_2 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_RNIUEQM_3_LC_20_7_2  (
            .in0(_gnd_net_),
            .in1(N__15290),
            .in2(N__14235),
            .in3(N__14113),
            .lcout(\fifo_inst.ftdi_output_inst.N_88_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.oTx_n_LC_20_7_3 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.oTx_n_LC_20_7_3 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.oTx_n_LC_20_7_3 .LUT_INIT=16'b1111111101001111;
    LogicCell40 \fifo_inst.ftdi_output_inst.oTx_n_LC_20_7_3  (
            .in0(N__14114),
            .in1(N__14197),
            .in2(N__14577),
            .in3(N__14336),
            .lcout(P1A4_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15052),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIBT9K_4_LC_20_7_5 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIBT9K_4_LC_20_7_5 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIBT9K_4_LC_20_7_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_RNIBT9K_4_LC_20_7_5  (
            .in0(N__14571),
            .in1(N__15388),
            .in2(_gnd_net_),
            .in3(N__15340),
            .lcout(\fifo_inst.ftdi_output_inst.oPacketRead_1_sqmuxa_1 ),
            .ltout(\fifo_inst.ftdi_output_inst.oPacketRead_1_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.oRamRdAddr_1_LC_20_7_6 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.oRamRdAddr_1_LC_20_7_6 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.oRamRdAddr_1_LC_20_7_6 .LUT_INIT=16'b0011110011001100;
    LogicCell40 \fifo_inst.ftdi_output_inst.oRamRdAddr_1_LC_20_7_6  (
            .in0(_gnd_net_),
            .in1(N__14149),
            .in2(N__14181),
            .in3(N__14173),
            .lcout(\fifo_inst.wRamRdAddr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15052),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.oRamRdAddr_2_LC_20_7_7 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.oRamRdAddr_2_LC_20_7_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.oRamRdAddr_2_LC_20_7_7 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \fifo_inst.ftdi_output_inst.oRamRdAddr_2_LC_20_7_7  (
            .in0(N__14174),
            .in1(N__14126),
            .in2(N__14156),
            .in3(N__14136),
            .lcout(\fifo_inst.wRamRdAddr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15052),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_3_LC_20_8_0 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_3_LC_20_8_0 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_3_LC_20_8_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_3_LC_20_8_0  (
            .in0(N__14324),
            .in1(N__14648),
            .in2(N__14679),
            .in3(N__14603),
            .lcout(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15048),
            .ce(),
            .sr(N__15241));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_4_LC_20_8_1 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_4_LC_20_8_1 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_4_LC_20_8_1 .LUT_INIT=16'b1111111100001010;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_4_LC_20_8_1  (
            .in0(N__15343),
            .in1(_gnd_net_),
            .in2(N__15409),
            .in3(N__14115),
            .lcout(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15048),
            .ce(),
            .sr(N__15241));
    defparam \fifo_inst.ftdi_output_inst.rWrDelay_LC_20_8_2 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rWrDelay_LC_20_8_2 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rWrDelay_LC_20_8_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \fifo_inst.ftdi_output_inst.rWrDelay_LC_20_8_2  (
            .in0(_gnd_net_),
            .in1(N__15392),
            .in2(_gnd_net_),
            .in3(N__15342),
            .lcout(\fifo_inst.ftdi_output_inst.rWrDelayZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15048),
            .ce(),
            .sr(N__15241));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_1_LC_20_8_3 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_1_LC_20_8_3 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_1_LC_20_8_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_1_LC_20_8_3  (
            .in0(N__14647),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14323),
            .lcout(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15048),
            .ce(),
            .sr(N__15241));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_2_LC_20_8_5 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_2_LC_20_8_5 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_2_LC_20_8_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_2_LC_20_8_5  (
            .in0(N__14694),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15048),
            .ce(),
            .sr(N__15241));
    defparam \fifo_inst.ftdi_output_inst.oRxFlag_LC_20_8_6 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.oRxFlag_LC_20_8_6 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.oRxFlag_LC_20_8_6 .LUT_INIT=16'b1111111101000100;
    LogicCell40 \fifo_inst.ftdi_output_inst.oRxFlag_LC_20_8_6  (
            .in0(N__14357),
            .in1(N__14773),
            .in2(_gnd_net_),
            .in3(N__14693),
            .lcout(P1A2_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15048),
            .ce(),
            .sr(N__15241));
    defparam \fifo_inst.ftdi_output_inst.oRx_n_LC_20_8_7 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.oRx_n_LC_20_8_7 .SEQ_MODE=4'b1001;
    defparam \fifo_inst.ftdi_output_inst.oRx_n_LC_20_8_7 .LUT_INIT=16'b1110110011101110;
    LogicCell40 \fifo_inst.ftdi_output_inst.oRx_n_LC_20_8_7  (
            .in0(N__14710),
            .in1(N__14356),
            .in2(N__14649),
            .in3(N__14325),
            .lcout(P1A3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15048),
            .ce(),
            .sr(N__15241));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIDTQ4_1_LC_20_9_1 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIDTQ4_1_LC_20_9_1 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIDTQ4_1_LC_20_9_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_RNIDTQ4_1_LC_20_9_1  (
            .in0(_gnd_net_),
            .in1(N__15283),
            .in2(_gnd_net_),
            .in3(N__14692),
            .lcout(\fifo_inst.ftdi_output_inst.rFifoState_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNO_0_0_LC_20_9_2 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNO_0_0_LC_20_9_2 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNO_0_0_LC_20_9_2 .LUT_INIT=16'b1000110000000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_RNO_0_0_LC_20_9_2  (
            .in0(N__14669),
            .in1(N__14636),
            .in2(N__14607),
            .in3(N__14322),
            .lcout(),
            .ltout(\fifo_inst.ftdi_output_inst.N_87_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_0_LC_20_9_3 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_0_LC_20_9_3 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_0_LC_20_9_3 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_0_LC_20_9_3  (
            .in0(N__14573),
            .in1(N__14358),
            .in2(N__14343),
            .in3(N__14340),
            .lcout(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15041),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_7_LC_20_10_1 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_7_LC_20_10_1 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_7_LC_20_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rRxData_esr_7_LC_20_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14307),
            .lcout(wRxFifoData_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15034),
            .ce(N__14266),
            .sr(N__15232));
    defparam ioFifoData_iobuf_RNO_3_LC_21_1_2.C_ON=1'b0;
    defparam ioFifoData_iobuf_RNO_3_LC_21_1_2.SEQ_MODE=4'b0000;
    defparam ioFifoData_iobuf_RNO_3_LC_21_1_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 ioFifoData_iobuf_RNO_3_LC_21_1_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15432),
            .lcout(N_1260_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ioFifoData_iobuf_RNO_2_LC_21_4_0.C_ON=1'b0;
    defparam ioFifoData_iobuf_RNO_2_LC_21_4_0.SEQ_MODE=4'b0000;
    defparam ioFifoData_iobuf_RNO_2_LC_21_4_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 ioFifoData_iobuf_RNO_2_LC_21_4_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15312),
            .lcout(N_1259_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.oTx_n_rep3_ess_LC_21_6_1 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.oTx_n_rep3_ess_LC_21_6_1 .SEQ_MODE=4'b1001;
    defparam \fifo_inst.ftdi_output_inst.oTx_n_rep3_ess_LC_21_6_1 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \fifo_inst.ftdi_output_inst.oTx_n_rep3_ess_LC_21_6_1  (
            .in0(N__15360),
            .in1(_gnd_net_),
            .in2(N__15423),
            .in3(_gnd_net_),
            .lcout(oTx_n_rep3_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15054),
            .ce(N__15303),
            .sr(N__15249));
    defparam \fifo_inst.ftdi_output_inst.oTx_n_rep2_ess_LC_21_6_2 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.oTx_n_rep2_ess_LC_21_6_2 .SEQ_MODE=4'b1001;
    defparam \fifo_inst.ftdi_output_inst.oTx_n_rep2_ess_LC_21_6_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.oTx_n_rep2_ess_LC_21_6_2  (
            .in0(_gnd_net_),
            .in1(N__15417),
            .in2(_gnd_net_),
            .in3(N__15359),
            .lcout(oTx_n_rep2_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15054),
            .ce(N__15303),
            .sr(N__15249));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_21_10_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_21_10_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_21_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_21_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15171),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15042),
            .ce(N__14868),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_21_10_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_21_10_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_21_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_21_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15110),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__15042),
            .ce(N__14868),
            .sr(_gnd_net_));
endmodule // top
