// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Mar 29 2020 11:31:56

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    ioFifoData,
    P1A9,
    P1A1,
    P1A8,
    oRx_n,
    P1A7,
    P1A3,
    iTxE_n,
    iRxF_n,
    iClk,
    P1A2,
    BTN_N,
    BTN1,
    oTx_n,
    P1A4);

    inout [7:0] ioFifoData;
    output P1A9;
    input P1A1;
    output P1A8;
    output oRx_n;
    output P1A7;
    output P1A3;
    input iTxE_n;
    input iRxF_n;
    input iClk;
    output P1A2;
    input BTN_N;
    input BTN1;
    output oTx_n;
    output P1A4;

    wire N__13366;
    wire N__13352;
    wire N__13351;
    wire N__13350;
    wire N__13343;
    wire N__13342;
    wire N__13341;
    wire N__13334;
    wire N__13333;
    wire N__13332;
    wire N__13325;
    wire N__13324;
    wire N__13323;
    wire N__13316;
    wire N__13315;
    wire N__13314;
    wire N__13307;
    wire N__13306;
    wire N__13305;
    wire N__13298;
    wire N__13297;
    wire N__13296;
    wire N__13289;
    wire N__13288;
    wire N__13287;
    wire N__13280;
    wire N__13279;
    wire N__13278;
    wire N__13271;
    wire N__13270;
    wire N__13269;
    wire N__13262;
    wire N__13261;
    wire N__13260;
    wire N__13253;
    wire N__13252;
    wire N__13251;
    wire N__13244;
    wire N__13243;
    wire N__13242;
    wire N__13235;
    wire N__13234;
    wire N__13233;
    wire N__13226;
    wire N__13225;
    wire N__13224;
    wire N__13217;
    wire N__13216;
    wire N__13215;
    wire N__13208;
    wire N__13207;
    wire N__13206;
    wire N__13199;
    wire N__13198;
    wire N__13197;
    wire N__13190;
    wire N__13189;
    wire N__13188;
    wire N__13181;
    wire N__13180;
    wire N__13179;
    wire N__13162;
    wire N__13159;
    wire N__13158;
    wire N__13155;
    wire N__13152;
    wire N__13147;
    wire N__13144;
    wire N__13143;
    wire N__13140;
    wire N__13137;
    wire N__13132;
    wire N__13129;
    wire N__13128;
    wire N__13125;
    wire N__13122;
    wire N__13119;
    wire N__13116;
    wire N__13111;
    wire N__13108;
    wire N__13107;
    wire N__13104;
    wire N__13101;
    wire N__13096;
    wire N__13093;
    wire N__13090;
    wire N__13089;
    wire N__13086;
    wire N__13083;
    wire N__13078;
    wire N__13077;
    wire N__13076;
    wire N__13075;
    wire N__13074;
    wire N__13073;
    wire N__13072;
    wire N__13071;
    wire N__13068;
    wire N__13065;
    wire N__13062;
    wire N__13059;
    wire N__13056;
    wire N__13055;
    wire N__13052;
    wire N__13049;
    wire N__13046;
    wire N__13045;
    wire N__13044;
    wire N__13043;
    wire N__13042;
    wire N__13041;
    wire N__13034;
    wire N__13023;
    wire N__13020;
    wire N__13017;
    wire N__13016;
    wire N__13013;
    wire N__13012;
    wire N__13009;
    wire N__13008;
    wire N__13005;
    wire N__13004;
    wire N__13003;
    wire N__13002;
    wire N__12999;
    wire N__12998;
    wire N__12997;
    wire N__12996;
    wire N__12993;
    wire N__12988;
    wire N__12973;
    wire N__12972;
    wire N__12969;
    wire N__12966;
    wire N__12965;
    wire N__12962;
    wire N__12961;
    wire N__12960;
    wire N__12957;
    wire N__12954;
    wire N__12953;
    wire N__12950;
    wire N__12949;
    wire N__12946;
    wire N__12945;
    wire N__12944;
    wire N__12939;
    wire N__12936;
    wire N__12923;
    wire N__12920;
    wire N__12917;
    wire N__12912;
    wire N__12901;
    wire N__12898;
    wire N__12893;
    wire N__12890;
    wire N__12883;
    wire N__12880;
    wire N__12877;
    wire N__12874;
    wire N__12871;
    wire N__12866;
    wire N__12863;
    wire N__12858;
    wire N__12855;
    wire N__12850;
    wire N__12849;
    wire N__12848;
    wire N__12845;
    wire N__12842;
    wire N__12839;
    wire N__12832;
    wire N__12831;
    wire N__12830;
    wire N__12829;
    wire N__12828;
    wire N__12827;
    wire N__12826;
    wire N__12825;
    wire N__12824;
    wire N__12823;
    wire N__12822;
    wire N__12821;
    wire N__12820;
    wire N__12819;
    wire N__12818;
    wire N__12817;
    wire N__12816;
    wire N__12815;
    wire N__12814;
    wire N__12813;
    wire N__12812;
    wire N__12811;
    wire N__12810;
    wire N__12809;
    wire N__12808;
    wire N__12807;
    wire N__12806;
    wire N__12805;
    wire N__12804;
    wire N__12803;
    wire N__12802;
    wire N__12801;
    wire N__12800;
    wire N__12799;
    wire N__12798;
    wire N__12797;
    wire N__12796;
    wire N__12795;
    wire N__12794;
    wire N__12793;
    wire N__12792;
    wire N__12791;
    wire N__12790;
    wire N__12789;
    wire N__12788;
    wire N__12787;
    wire N__12786;
    wire N__12785;
    wire N__12784;
    wire N__12783;
    wire N__12782;
    wire N__12781;
    wire N__12780;
    wire N__12779;
    wire N__12778;
    wire N__12777;
    wire N__12776;
    wire N__12775;
    wire N__12774;
    wire N__12773;
    wire N__12772;
    wire N__12771;
    wire N__12770;
    wire N__12769;
    wire N__12640;
    wire N__12637;
    wire N__12636;
    wire N__12633;
    wire N__12630;
    wire N__12627;
    wire N__12624;
    wire N__12621;
    wire N__12618;
    wire N__12613;
    wire N__12612;
    wire N__12609;
    wire N__12606;
    wire N__12601;
    wire N__12598;
    wire N__12595;
    wire N__12594;
    wire N__12591;
    wire N__12588;
    wire N__12583;
    wire N__12580;
    wire N__12579;
    wire N__12576;
    wire N__12573;
    wire N__12570;
    wire N__12565;
    wire N__12562;
    wire N__12559;
    wire N__12558;
    wire N__12555;
    wire N__12552;
    wire N__12547;
    wire N__12544;
    wire N__12543;
    wire N__12540;
    wire N__12537;
    wire N__12532;
    wire N__12529;
    wire N__12526;
    wire N__12525;
    wire N__12522;
    wire N__12519;
    wire N__12514;
    wire N__12511;
    wire N__12510;
    wire N__12507;
    wire N__12504;
    wire N__12501;
    wire N__12496;
    wire N__12493;
    wire N__12492;
    wire N__12489;
    wire N__12486;
    wire N__12481;
    wire N__12478;
    wire N__12475;
    wire N__12472;
    wire N__12469;
    wire N__12466;
    wire N__12463;
    wire N__12460;
    wire N__12457;
    wire N__12454;
    wire N__12451;
    wire N__12448;
    wire N__12445;
    wire N__12442;
    wire N__12441;
    wire N__12440;
    wire N__12439;
    wire N__12438;
    wire N__12437;
    wire N__12434;
    wire N__12433;
    wire N__12432;
    wire N__12429;
    wire N__12428;
    wire N__12425;
    wire N__12424;
    wire N__12423;
    wire N__12422;
    wire N__12421;
    wire N__12418;
    wire N__12415;
    wire N__12410;
    wire N__12407;
    wire N__12404;
    wire N__12401;
    wire N__12398;
    wire N__12395;
    wire N__12392;
    wire N__12389;
    wire N__12386;
    wire N__12383;
    wire N__12380;
    wire N__12377;
    wire N__12376;
    wire N__12375;
    wire N__12372;
    wire N__12369;
    wire N__12366;
    wire N__12363;
    wire N__12360;
    wire N__12357;
    wire N__12354;
    wire N__12353;
    wire N__12350;
    wire N__12347;
    wire N__12346;
    wire N__12345;
    wire N__12344;
    wire N__12341;
    wire N__12340;
    wire N__12301;
    wire N__12298;
    wire N__12295;
    wire N__12292;
    wire N__12289;
    wire N__12286;
    wire N__12283;
    wire N__12282;
    wire N__12281;
    wire N__12278;
    wire N__12275;
    wire N__12272;
    wire N__12269;
    wire N__12266;
    wire N__12263;
    wire N__12260;
    wire N__12257;
    wire N__12250;
    wire N__12249;
    wire N__12248;
    wire N__12247;
    wire N__12246;
    wire N__12245;
    wire N__12244;
    wire N__12243;
    wire N__12240;
    wire N__12237;
    wire N__12234;
    wire N__12231;
    wire N__12230;
    wire N__12225;
    wire N__12224;
    wire N__12223;
    wire N__12218;
    wire N__12215;
    wire N__12212;
    wire N__12205;
    wire N__12202;
    wire N__12197;
    wire N__12196;
    wire N__12193;
    wire N__12190;
    wire N__12187;
    wire N__12180;
    wire N__12177;
    wire N__12174;
    wire N__12163;
    wire N__12162;
    wire N__12159;
    wire N__12158;
    wire N__12157;
    wire N__12154;
    wire N__12147;
    wire N__12142;
    wire N__12139;
    wire N__12136;
    wire N__12135;
    wire N__12134;
    wire N__12133;
    wire N__12132;
    wire N__12127;
    wire N__12124;
    wire N__12119;
    wire N__12112;
    wire N__12109;
    wire N__12106;
    wire N__12103;
    wire N__12100;
    wire N__12097;
    wire N__12094;
    wire N__12091;
    wire N__12088;
    wire N__12085;
    wire N__12084;
    wire N__12083;
    wire N__12082;
    wire N__12081;
    wire N__12080;
    wire N__12079;
    wire N__12078;
    wire N__12075;
    wire N__12070;
    wire N__12063;
    wire N__12058;
    wire N__12049;
    wire N__12048;
    wire N__12047;
    wire N__12046;
    wire N__12045;
    wire N__12044;
    wire N__12043;
    wire N__12042;
    wire N__12039;
    wire N__12034;
    wire N__12029;
    wire N__12024;
    wire N__12019;
    wire N__12010;
    wire N__12009;
    wire N__12008;
    wire N__12007;
    wire N__12006;
    wire N__12003;
    wire N__12000;
    wire N__11995;
    wire N__11990;
    wire N__11983;
    wire N__11980;
    wire N__11979;
    wire N__11978;
    wire N__11977;
    wire N__11976;
    wire N__11975;
    wire N__11972;
    wire N__11965;
    wire N__11960;
    wire N__11953;
    wire N__11950;
    wire N__11947;
    wire N__11944;
    wire N__11943;
    wire N__11942;
    wire N__11935;
    wire N__11932;
    wire N__11929;
    wire N__11926;
    wire N__11925;
    wire N__11922;
    wire N__11921;
    wire N__11920;
    wire N__11919;
    wire N__11918;
    wire N__11917;
    wire N__11914;
    wire N__11911;
    wire N__11902;
    wire N__11899;
    wire N__11890;
    wire N__11887;
    wire N__11884;
    wire N__11883;
    wire N__11882;
    wire N__11879;
    wire N__11876;
    wire N__11875;
    wire N__11874;
    wire N__11873;
    wire N__11870;
    wire N__11867;
    wire N__11862;
    wire N__11857;
    wire N__11848;
    wire N__11845;
    wire N__11842;
    wire N__11839;
    wire N__11836;
    wire N__11833;
    wire N__11832;
    wire N__11829;
    wire N__11826;
    wire N__11821;
    wire N__11820;
    wire N__11819;
    wire N__11818;
    wire N__11815;
    wire N__11812;
    wire N__11809;
    wire N__11808;
    wire N__11805;
    wire N__11804;
    wire N__11803;
    wire N__11802;
    wire N__11801;
    wire N__11798;
    wire N__11795;
    wire N__11792;
    wire N__11789;
    wire N__11784;
    wire N__11779;
    wire N__11776;
    wire N__11773;
    wire N__11764;
    wire N__11755;
    wire N__11754;
    wire N__11753;
    wire N__11750;
    wire N__11749;
    wire N__11748;
    wire N__11747;
    wire N__11746;
    wire N__11743;
    wire N__11740;
    wire N__11737;
    wire N__11730;
    wire N__11727;
    wire N__11724;
    wire N__11719;
    wire N__11716;
    wire N__11713;
    wire N__11712;
    wire N__11711;
    wire N__11708;
    wire N__11705;
    wire N__11702;
    wire N__11699;
    wire N__11696;
    wire N__11693;
    wire N__11680;
    wire N__11679;
    wire N__11678;
    wire N__11677;
    wire N__11676;
    wire N__11675;
    wire N__11674;
    wire N__11671;
    wire N__11670;
    wire N__11667;
    wire N__11666;
    wire N__11665;
    wire N__11662;
    wire N__11661;
    wire N__11660;
    wire N__11659;
    wire N__11658;
    wire N__11657;
    wire N__11656;
    wire N__11653;
    wire N__11652;
    wire N__11651;
    wire N__11648;
    wire N__11641;
    wire N__11636;
    wire N__11625;
    wire N__11614;
    wire N__11607;
    wire N__11604;
    wire N__11603;
    wire N__11602;
    wire N__11595;
    wire N__11592;
    wire N__11589;
    wire N__11584;
    wire N__11581;
    wire N__11576;
    wire N__11569;
    wire N__11566;
    wire N__11563;
    wire N__11562;
    wire N__11561;
    wire N__11554;
    wire N__11551;
    wire N__11548;
    wire N__11545;
    wire N__11542;
    wire N__11541;
    wire N__11540;
    wire N__11539;
    wire N__11538;
    wire N__11537;
    wire N__11536;
    wire N__11535;
    wire N__11534;
    wire N__11531;
    wire N__11524;
    wire N__11523;
    wire N__11522;
    wire N__11517;
    wire N__11512;
    wire N__11511;
    wire N__11508;
    wire N__11507;
    wire N__11504;
    wire N__11501;
    wire N__11496;
    wire N__11491;
    wire N__11488;
    wire N__11483;
    wire N__11480;
    wire N__11475;
    wire N__11472;
    wire N__11461;
    wire N__11460;
    wire N__11459;
    wire N__11456;
    wire N__11453;
    wire N__11450;
    wire N__11443;
    wire N__11442;
    wire N__11441;
    wire N__11438;
    wire N__11437;
    wire N__11436;
    wire N__11435;
    wire N__11434;
    wire N__11433;
    wire N__11432;
    wire N__11429;
    wire N__11428;
    wire N__11427;
    wire N__11424;
    wire N__11423;
    wire N__11422;
    wire N__11419;
    wire N__11412;
    wire N__11409;
    wire N__11408;
    wire N__11407;
    wire N__11406;
    wire N__11399;
    wire N__11396;
    wire N__11395;
    wire N__11394;
    wire N__11393;
    wire N__11392;
    wire N__11391;
    wire N__11388;
    wire N__11385;
    wire N__11380;
    wire N__11375;
    wire N__11372;
    wire N__11371;
    wire N__11370;
    wire N__11363;
    wire N__11360;
    wire N__11357;
    wire N__11350;
    wire N__11345;
    wire N__11342;
    wire N__11339;
    wire N__11336;
    wire N__11331;
    wire N__11328;
    wire N__11325;
    wire N__11318;
    wire N__11313;
    wire N__11296;
    wire N__11293;
    wire N__11290;
    wire N__11287;
    wire N__11284;
    wire N__11281;
    wire N__11278;
    wire N__11275;
    wire N__11272;
    wire N__11269;
    wire N__11266;
    wire N__11263;
    wire N__11260;
    wire N__11257;
    wire N__11254;
    wire N__11251;
    wire N__11250;
    wire N__11249;
    wire N__11248;
    wire N__11245;
    wire N__11242;
    wire N__11241;
    wire N__11240;
    wire N__11239;
    wire N__11236;
    wire N__11235;
    wire N__11232;
    wire N__11227;
    wire N__11224;
    wire N__11215;
    wire N__11212;
    wire N__11209;
    wire N__11206;
    wire N__11201;
    wire N__11198;
    wire N__11195;
    wire N__11188;
    wire N__11185;
    wire N__11182;
    wire N__11181;
    wire N__11178;
    wire N__11175;
    wire N__11172;
    wire N__11171;
    wire N__11170;
    wire N__11167;
    wire N__11164;
    wire N__11159;
    wire N__11156;
    wire N__11149;
    wire N__11148;
    wire N__11147;
    wire N__11146;
    wire N__11143;
    wire N__11138;
    wire N__11135;
    wire N__11134;
    wire N__11131;
    wire N__11130;
    wire N__11129;
    wire N__11126;
    wire N__11125;
    wire N__11124;
    wire N__11123;
    wire N__11120;
    wire N__11119;
    wire N__11118;
    wire N__11117;
    wire N__11116;
    wire N__11115;
    wire N__11114;
    wire N__11113;
    wire N__11112;
    wire N__11111;
    wire N__11074;
    wire N__11071;
    wire N__11068;
    wire N__11065;
    wire N__11062;
    wire N__11059;
    wire N__11056;
    wire N__11055;
    wire N__11054;
    wire N__11051;
    wire N__11048;
    wire N__11045;
    wire N__11044;
    wire N__11043;
    wire N__11042;
    wire N__11041;
    wire N__11040;
    wire N__11039;
    wire N__11038;
    wire N__11031;
    wire N__11028;
    wire N__11019;
    wire N__11016;
    wire N__11013;
    wire N__11010;
    wire N__11007;
    wire N__11000;
    wire N__10997;
    wire N__10994;
    wire N__10991;
    wire N__10986;
    wire N__10983;
    wire N__10980;
    wire N__10975;
    wire N__10974;
    wire N__10973;
    wire N__10972;
    wire N__10971;
    wire N__10970;
    wire N__10969;
    wire N__10966;
    wire N__10957;
    wire N__10956;
    wire N__10953;
    wire N__10950;
    wire N__10947;
    wire N__10946;
    wire N__10943;
    wire N__10940;
    wire N__10939;
    wire N__10934;
    wire N__10931;
    wire N__10928;
    wire N__10923;
    wire N__10920;
    wire N__10917;
    wire N__10906;
    wire N__10903;
    wire N__10900;
    wire N__10897;
    wire N__10894;
    wire N__10891;
    wire N__10888;
    wire N__10887;
    wire N__10884;
    wire N__10883;
    wire N__10880;
    wire N__10875;
    wire N__10870;
    wire N__10867;
    wire N__10864;
    wire N__10861;
    wire N__10860;
    wire N__10859;
    wire N__10856;
    wire N__10853;
    wire N__10852;
    wire N__10849;
    wire N__10846;
    wire N__10843;
    wire N__10840;
    wire N__10837;
    wire N__10828;
    wire N__10827;
    wire N__10822;
    wire N__10819;
    wire N__10816;
    wire N__10813;
    wire N__10810;
    wire N__10807;
    wire N__10804;
    wire N__10801;
    wire N__10798;
    wire N__10795;
    wire N__10792;
    wire N__10791;
    wire N__10790;
    wire N__10787;
    wire N__10784;
    wire N__10781;
    wire N__10774;
    wire N__10771;
    wire N__10770;
    wire N__10769;
    wire N__10768;
    wire N__10767;
    wire N__10764;
    wire N__10759;
    wire N__10754;
    wire N__10747;
    wire N__10744;
    wire N__10741;
    wire N__10738;
    wire N__10735;
    wire N__10732;
    wire N__10729;
    wire N__10726;
    wire N__10725;
    wire N__10722;
    wire N__10721;
    wire N__10718;
    wire N__10715;
    wire N__10712;
    wire N__10705;
    wire N__10702;
    wire N__10699;
    wire N__10696;
    wire N__10695;
    wire N__10694;
    wire N__10687;
    wire N__10684;
    wire N__10683;
    wire N__10682;
    wire N__10679;
    wire N__10676;
    wire N__10675;
    wire N__10666;
    wire N__10663;
    wire N__10662;
    wire N__10661;
    wire N__10660;
    wire N__10659;
    wire N__10648;
    wire N__10645;
    wire N__10642;
    wire N__10641;
    wire N__10640;
    wire N__10639;
    wire N__10638;
    wire N__10635;
    wire N__10634;
    wire N__10633;
    wire N__10630;
    wire N__10627;
    wire N__10626;
    wire N__10625;
    wire N__10622;
    wire N__10619;
    wire N__10616;
    wire N__10613;
    wire N__10610;
    wire N__10607;
    wire N__10604;
    wire N__10601;
    wire N__10598;
    wire N__10595;
    wire N__10592;
    wire N__10585;
    wire N__10582;
    wire N__10579;
    wire N__10576;
    wire N__10573;
    wire N__10570;
    wire N__10567;
    wire N__10564;
    wire N__10559;
    wire N__10556;
    wire N__10553;
    wire N__10546;
    wire N__10543;
    wire N__10540;
    wire N__10537;
    wire N__10532;
    wire N__10529;
    wire N__10526;
    wire N__10523;
    wire N__10520;
    wire N__10517;
    wire N__10514;
    wire N__10509;
    wire N__10504;
    wire N__10501;
    wire N__10498;
    wire N__10497;
    wire N__10496;
    wire N__10495;
    wire N__10486;
    wire N__10483;
    wire N__10480;
    wire N__10477;
    wire N__10474;
    wire N__10471;
    wire N__10470;
    wire N__10467;
    wire N__10464;
    wire N__10461;
    wire N__10456;
    wire N__10453;
    wire N__10452;
    wire N__10451;
    wire N__10450;
    wire N__10447;
    wire N__10444;
    wire N__10439;
    wire N__10432;
    wire N__10429;
    wire N__10428;
    wire N__10425;
    wire N__10422;
    wire N__10417;
    wire N__10414;
    wire N__10413;
    wire N__10412;
    wire N__10409;
    wire N__10408;
    wire N__10405;
    wire N__10404;
    wire N__10403;
    wire N__10400;
    wire N__10397;
    wire N__10392;
    wire N__10389;
    wire N__10386;
    wire N__10377;
    wire N__10372;
    wire N__10369;
    wire N__10368;
    wire N__10367;
    wire N__10364;
    wire N__10359;
    wire N__10356;
    wire N__10351;
    wire N__10348;
    wire N__10347;
    wire N__10344;
    wire N__10343;
    wire N__10342;
    wire N__10341;
    wire N__10340;
    wire N__10337;
    wire N__10336;
    wire N__10335;
    wire N__10334;
    wire N__10333;
    wire N__10330;
    wire N__10323;
    wire N__10322;
    wire N__10321;
    wire N__10316;
    wire N__10309;
    wire N__10306;
    wire N__10303;
    wire N__10302;
    wire N__10301;
    wire N__10298;
    wire N__10295;
    wire N__10292;
    wire N__10285;
    wire N__10282;
    wire N__10279;
    wire N__10276;
    wire N__10273;
    wire N__10270;
    wire N__10265;
    wire N__10252;
    wire N__10251;
    wire N__10248;
    wire N__10245;
    wire N__10242;
    wire N__10239;
    wire N__10234;
    wire N__10233;
    wire N__10230;
    wire N__10227;
    wire N__10222;
    wire N__10219;
    wire N__10218;
    wire N__10217;
    wire N__10214;
    wire N__10211;
    wire N__10208;
    wire N__10201;
    wire N__10198;
    wire N__10195;
    wire N__10192;
    wire N__10189;
    wire N__10186;
    wire N__10183;
    wire N__10182;
    wire N__10179;
    wire N__10176;
    wire N__10175;
    wire N__10172;
    wire N__10169;
    wire N__10166;
    wire N__10159;
    wire N__10158;
    wire N__10155;
    wire N__10152;
    wire N__10151;
    wire N__10148;
    wire N__10145;
    wire N__10142;
    wire N__10141;
    wire N__10134;
    wire N__10131;
    wire N__10126;
    wire N__10123;
    wire N__10120;
    wire N__10117;
    wire N__10116;
    wire N__10113;
    wire N__10112;
    wire N__10109;
    wire N__10106;
    wire N__10103;
    wire N__10102;
    wire N__10095;
    wire N__10092;
    wire N__10087;
    wire N__10084;
    wire N__10081;
    wire N__10080;
    wire N__10079;
    wire N__10078;
    wire N__10075;
    wire N__10072;
    wire N__10071;
    wire N__10068;
    wire N__10065;
    wire N__10062;
    wire N__10061;
    wire N__10058;
    wire N__10055;
    wire N__10052;
    wire N__10049;
    wire N__10046;
    wire N__10043;
    wire N__10038;
    wire N__10033;
    wire N__10028;
    wire N__10027;
    wire N__10024;
    wire N__10019;
    wire N__10016;
    wire N__10009;
    wire N__10006;
    wire N__10003;
    wire N__10002;
    wire N__10001;
    wire N__9998;
    wire N__9995;
    wire N__9994;
    wire N__9993;
    wire N__9990;
    wire N__9987;
    wire N__9980;
    wire N__9973;
    wire N__9970;
    wire N__9967;
    wire N__9964;
    wire N__9963;
    wire N__9962;
    wire N__9961;
    wire N__9958;
    wire N__9953;
    wire N__9950;
    wire N__9943;
    wire N__9940;
    wire N__9939;
    wire N__9938;
    wire N__9935;
    wire N__9932;
    wire N__9929;
    wire N__9922;
    wire N__9919;
    wire N__9916;
    wire N__9915;
    wire N__9914;
    wire N__9911;
    wire N__9910;
    wire N__9907;
    wire N__9906;
    wire N__9903;
    wire N__9900;
    wire N__9897;
    wire N__9892;
    wire N__9883;
    wire N__9882;
    wire N__9881;
    wire N__9878;
    wire N__9871;
    wire N__9870;
    wire N__9869;
    wire N__9866;
    wire N__9863;
    wire N__9862;
    wire N__9861;
    wire N__9860;
    wire N__9857;
    wire N__9856;
    wire N__9855;
    wire N__9852;
    wire N__9849;
    wire N__9844;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9824;
    wire N__9821;
    wire N__9818;
    wire N__9813;
    wire N__9810;
    wire N__9807;
    wire N__9802;
    wire N__9801;
    wire N__9800;
    wire N__9797;
    wire N__9794;
    wire N__9791;
    wire N__9784;
    wire N__9781;
    wire N__9778;
    wire N__9775;
    wire N__9772;
    wire N__9771;
    wire N__9770;
    wire N__9765;
    wire N__9762;
    wire N__9761;
    wire N__9760;
    wire N__9759;
    wire N__9756;
    wire N__9753;
    wire N__9748;
    wire N__9747;
    wire N__9746;
    wire N__9743;
    wire N__9738;
    wire N__9735;
    wire N__9730;
    wire N__9721;
    wire N__9720;
    wire N__9717;
    wire N__9716;
    wire N__9715;
    wire N__9714;
    wire N__9713;
    wire N__9712;
    wire N__9711;
    wire N__9708;
    wire N__9707;
    wire N__9706;
    wire N__9705;
    wire N__9702;
    wire N__9697;
    wire N__9694;
    wire N__9689;
    wire N__9682;
    wire N__9677;
    wire N__9664;
    wire N__9661;
    wire N__9658;
    wire N__9655;
    wire N__9652;
    wire N__9651;
    wire N__9650;
    wire N__9647;
    wire N__9644;
    wire N__9641;
    wire N__9640;
    wire N__9639;
    wire N__9634;
    wire N__9631;
    wire N__9630;
    wire N__9629;
    wire N__9628;
    wire N__9627;
    wire N__9626;
    wire N__9625;
    wire N__9620;
    wire N__9617;
    wire N__9614;
    wire N__9607;
    wire N__9602;
    wire N__9599;
    wire N__9586;
    wire N__9583;
    wire N__9580;
    wire N__9577;
    wire N__9576;
    wire N__9575;
    wire N__9572;
    wire N__9571;
    wire N__9568;
    wire N__9565;
    wire N__9562;
    wire N__9561;
    wire N__9560;
    wire N__9559;
    wire N__9558;
    wire N__9557;
    wire N__9556;
    wire N__9553;
    wire N__9552;
    wire N__9551;
    wire N__9548;
    wire N__9543;
    wire N__9536;
    wire N__9531;
    wire N__9526;
    wire N__9523;
    wire N__9520;
    wire N__9505;
    wire N__9504;
    wire N__9503;
    wire N__9500;
    wire N__9499;
    wire N__9498;
    wire N__9497;
    wire N__9494;
    wire N__9491;
    wire N__9488;
    wire N__9487;
    wire N__9486;
    wire N__9483;
    wire N__9480;
    wire N__9479;
    wire N__9476;
    wire N__9471;
    wire N__9468;
    wire N__9465;
    wire N__9462;
    wire N__9459;
    wire N__9452;
    wire N__9439;
    wire N__9436;
    wire N__9435;
    wire N__9432;
    wire N__9431;
    wire N__9430;
    wire N__9429;
    wire N__9428;
    wire N__9425;
    wire N__9422;
    wire N__9421;
    wire N__9420;
    wire N__9419;
    wire N__9418;
    wire N__9417;
    wire N__9416;
    wire N__9413;
    wire N__9410;
    wire N__9405;
    wire N__9400;
    wire N__9397;
    wire N__9388;
    wire N__9385;
    wire N__9380;
    wire N__9367;
    wire N__9364;
    wire N__9363;
    wire N__9362;
    wire N__9355;
    wire N__9354;
    wire N__9353;
    wire N__9352;
    wire N__9351;
    wire N__9350;
    wire N__9349;
    wire N__9348;
    wire N__9347;
    wire N__9346;
    wire N__9343;
    wire N__9332;
    wire N__9327;
    wire N__9324;
    wire N__9321;
    wire N__9320;
    wire N__9319;
    wire N__9318;
    wire N__9317;
    wire N__9316;
    wire N__9315;
    wire N__9314;
    wire N__9313;
    wire N__9312;
    wire N__9311;
    wire N__9310;
    wire N__9309;
    wire N__9308;
    wire N__9305;
    wire N__9300;
    wire N__9287;
    wire N__9284;
    wire N__9281;
    wire N__9278;
    wire N__9271;
    wire N__9264;
    wire N__9259;
    wire N__9254;
    wire N__9241;
    wire N__9238;
    wire N__9237;
    wire N__9236;
    wire N__9235;
    wire N__9234;
    wire N__9231;
    wire N__9224;
    wire N__9223;
    wire N__9222;
    wire N__9221;
    wire N__9220;
    wire N__9219;
    wire N__9216;
    wire N__9213;
    wire N__9210;
    wire N__9205;
    wire N__9198;
    wire N__9187;
    wire N__9184;
    wire N__9181;
    wire N__9178;
    wire N__9175;
    wire N__9172;
    wire N__9169;
    wire N__9166;
    wire N__9163;
    wire N__9160;
    wire N__9157;
    wire N__9154;
    wire N__9153;
    wire N__9150;
    wire N__9149;
    wire N__9148;
    wire N__9139;
    wire N__9138;
    wire N__9137;
    wire N__9136;
    wire N__9135;
    wire N__9132;
    wire N__9123;
    wire N__9118;
    wire N__9115;
    wire N__9112;
    wire N__9109;
    wire N__9106;
    wire N__9103;
    wire N__9102;
    wire N__9099;
    wire N__9096;
    wire N__9093;
    wire N__9090;
    wire N__9085;
    wire N__9082;
    wire N__9081;
    wire N__9078;
    wire N__9075;
    wire N__9072;
    wire N__9069;
    wire N__9064;
    wire N__9061;
    wire N__9060;
    wire N__9057;
    wire N__9054;
    wire N__9053;
    wire N__9050;
    wire N__9047;
    wire N__9046;
    wire N__9043;
    wire N__9040;
    wire N__9037;
    wire N__9034;
    wire N__9031;
    wire N__9028;
    wire N__9025;
    wire N__9022;
    wire N__9019;
    wire N__9016;
    wire N__9007;
    wire N__9004;
    wire N__9001;
    wire N__8998;
    wire N__8995;
    wire N__8992;
    wire N__8989;
    wire N__8986;
    wire N__8985;
    wire N__8984;
    wire N__8983;
    wire N__8982;
    wire N__8981;
    wire N__8978;
    wire N__8969;
    wire N__8966;
    wire N__8959;
    wire N__8956;
    wire N__8953;
    wire N__8950;
    wire N__8947;
    wire N__8944;
    wire N__8941;
    wire N__8938;
    wire N__8935;
    wire N__8932;
    wire N__8929;
    wire N__8926;
    wire N__8923;
    wire N__8920;
    wire N__8917;
    wire N__8914;
    wire N__8911;
    wire N__8908;
    wire N__8905;
    wire N__8902;
    wire N__8899;
    wire N__8896;
    wire N__8893;
    wire N__8890;
    wire N__8887;
    wire N__8884;
    wire N__8881;
    wire N__8878;
    wire N__8875;
    wire N__8872;
    wire N__8869;
    wire N__8866;
    wire N__8863;
    wire N__8860;
    wire N__8857;
    wire N__8854;
    wire N__8851;
    wire N__8848;
    wire N__8845;
    wire N__8842;
    wire N__8839;
    wire N__8836;
    wire N__8833;
    wire N__8830;
    wire N__8827;
    wire N__8824;
    wire N__8821;
    wire N__8818;
    wire N__8815;
    wire N__8812;
    wire N__8809;
    wire N__8806;
    wire N__8803;
    wire N__8800;
    wire N__8797;
    wire N__8794;
    wire N__8791;
    wire N__8788;
    wire N__8785;
    wire N__8782;
    wire N__8779;
    wire N__8776;
    wire N__8773;
    wire N__8770;
    wire N__8767;
    wire N__8764;
    wire N__8761;
    wire N__8758;
    wire N__8755;
    wire N__8752;
    wire N__8749;
    wire N__8746;
    wire N__8743;
    wire N__8740;
    wire N__8737;
    wire N__8734;
    wire N__8731;
    wire N__8728;
    wire N__8725;
    wire N__8722;
    wire N__8719;
    wire N__8716;
    wire N__8713;
    wire N__8710;
    wire N__8707;
    wire N__8706;
    wire N__8703;
    wire N__8702;
    wire N__8701;
    wire N__8698;
    wire N__8695;
    wire N__8692;
    wire N__8689;
    wire N__8686;
    wire N__8683;
    wire N__8674;
    wire N__8673;
    wire N__8672;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8662;
    wire N__8661;
    wire N__8660;
    wire N__8655;
    wire N__8652;
    wire N__8645;
    wire N__8642;
    wire N__8635;
    wire N__8632;
    wire N__8631;
    wire N__8628;
    wire N__8625;
    wire N__8622;
    wire N__8617;
    wire N__8614;
    wire N__8613;
    wire N__8610;
    wire N__8609;
    wire N__8606;
    wire N__8605;
    wire N__8604;
    wire N__8601;
    wire N__8598;
    wire N__8591;
    wire N__8586;
    wire N__8581;
    wire N__8578;
    wire N__8575;
    wire N__8572;
    wire N__8569;
    wire N__8568;
    wire N__8565;
    wire N__8562;
    wire N__8557;
    wire N__8556;
    wire N__8555;
    wire N__8554;
    wire N__8553;
    wire N__8552;
    wire N__8551;
    wire N__8548;
    wire N__8543;
    wire N__8540;
    wire N__8533;
    wire N__8524;
    wire N__8521;
    wire N__8518;
    wire N__8515;
    wire N__8514;
    wire N__8511;
    wire N__8510;
    wire N__8507;
    wire N__8506;
    wire N__8503;
    wire N__8500;
    wire N__8497;
    wire N__8494;
    wire N__8491;
    wire N__8488;
    wire N__8483;
    wire N__8482;
    wire N__8479;
    wire N__8476;
    wire N__8473;
    wire N__8470;
    wire N__8461;
    wire N__8460;
    wire N__8459;
    wire N__8456;
    wire N__8453;
    wire N__8450;
    wire N__8449;
    wire N__8446;
    wire N__8441;
    wire N__8438;
    wire N__8431;
    wire N__8430;
    wire N__8427;
    wire N__8424;
    wire N__8419;
    wire N__8418;
    wire N__8415;
    wire N__8412;
    wire N__8409;
    wire N__8406;
    wire N__8403;
    wire N__8400;
    wire N__8395;
    wire N__8392;
    wire N__8389;
    wire N__8386;
    wire N__8383;
    wire N__8380;
    wire N__8377;
    wire N__8374;
    wire N__8371;
    wire N__8368;
    wire N__8365;
    wire N__8362;
    wire N__8361;
    wire N__8358;
    wire N__8355;
    wire N__8350;
    wire N__8347;
    wire N__8344;
    wire N__8343;
    wire N__8340;
    wire N__8337;
    wire N__8332;
    wire N__8329;
    wire N__8326;
    wire N__8325;
    wire N__8322;
    wire N__8319;
    wire N__8314;
    wire N__8311;
    wire N__8308;
    wire N__8305;
    wire N__8302;
    wire N__8299;
    wire N__8296;
    wire N__8293;
    wire N__8290;
    wire N__8287;
    wire N__8284;
    wire N__8281;
    wire N__8280;
    wire N__8279;
    wire N__8276;
    wire N__8273;
    wire N__8270;
    wire N__8265;
    wire N__8260;
    wire N__8257;
    wire N__8256;
    wire N__8253;
    wire N__8250;
    wire N__8247;
    wire N__8244;
    wire N__8241;
    wire N__8236;
    wire N__8235;
    wire N__8234;
    wire N__8231;
    wire N__8226;
    wire N__8221;
    wire N__8220;
    wire N__8217;
    wire N__8214;
    wire N__8211;
    wire N__8208;
    wire N__8205;
    wire N__8202;
    wire N__8197;
    wire N__8196;
    wire N__8195;
    wire N__8192;
    wire N__8187;
    wire N__8182;
    wire N__8181;
    wire N__8176;
    wire N__8173;
    wire N__8170;
    wire N__8167;
    wire N__8166;
    wire N__8163;
    wire N__8160;
    wire N__8155;
    wire N__8152;
    wire N__8149;
    wire N__8146;
    wire N__8145;
    wire N__8140;
    wire N__8137;
    wire N__8134;
    wire N__8131;
    wire N__8130;
    wire N__8125;
    wire N__8122;
    wire N__8119;
    wire N__8116;
    wire N__8115;
    wire N__8114;
    wire N__8111;
    wire N__8108;
    wire N__8103;
    wire N__8100;
    wire N__8095;
    wire N__8092;
    wire N__8091;
    wire N__8088;
    wire N__8085;
    wire N__8080;
    wire N__8079;
    wire N__8074;
    wire N__8071;
    wire N__8068;
    wire N__8065;
    wire N__8062;
    wire N__8059;
    wire N__8056;
    wire N__8053;
    wire N__8050;
    wire N__8047;
    wire N__8046;
    wire N__8043;
    wire N__8040;
    wire N__8039;
    wire N__8036;
    wire N__8033;
    wire N__8032;
    wire N__8031;
    wire N__8030;
    wire N__8029;
    wire N__8028;
    wire N__8027;
    wire N__8026;
    wire N__8023;
    wire N__8022;
    wire N__8017;
    wire N__8012;
    wire N__8005;
    wire N__8002;
    wire N__7995;
    wire N__7984;
    wire N__7981;
    wire N__7978;
    wire N__7975;
    wire N__7972;
    wire N__7969;
    wire N__7968;
    wire N__7965;
    wire N__7962;
    wire N__7957;
    wire N__7954;
    wire N__7951;
    wire N__7948;
    wire N__7945;
    wire N__7942;
    wire N__7941;
    wire N__7938;
    wire N__7935;
    wire N__7930;
    wire N__7929;
    wire N__7926;
    wire N__7923;
    wire N__7920;
    wire N__7915;
    wire N__7914;
    wire N__7913;
    wire N__7908;
    wire N__7905;
    wire N__7900;
    wire N__7897;
    wire N__7896;
    wire N__7895;
    wire N__7890;
    wire N__7887;
    wire N__7882;
    wire N__7881;
    wire N__7876;
    wire N__7873;
    wire N__7870;
    wire N__7869;
    wire N__7866;
    wire N__7863;
    wire N__7860;
    wire N__7857;
    wire N__7854;
    wire N__7851;
    wire N__7848;
    wire N__7847;
    wire N__7844;
    wire N__7841;
    wire N__7838;
    wire N__7831;
    wire N__7830;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7819;
    wire N__7814;
    wire N__7811;
    wire N__7808;
    wire N__7805;
    wire N__7802;
    wire N__7799;
    wire N__7796;
    wire N__7791;
    wire N__7788;
    wire N__7785;
    wire N__7784;
    wire N__7781;
    wire N__7778;
    wire N__7775;
    wire N__7768;
    wire N__7767;
    wire N__7762;
    wire N__7759;
    wire N__7756;
    wire N__7753;
    wire N__7750;
    wire N__7747;
    wire N__7744;
    wire N__7741;
    wire N__7738;
    wire N__7735;
    wire N__7732;
    wire N__7729;
    wire N__7728;
    wire N__7725;
    wire N__7722;
    wire N__7717;
    wire N__7716;
    wire N__7713;
    wire N__7710;
    wire N__7705;
    wire N__7704;
    wire N__7701;
    wire N__7698;
    wire N__7695;
    wire N__7690;
    wire N__7687;
    wire N__7684;
    wire N__7681;
    wire N__7678;
    wire N__7675;
    wire N__7672;
    wire N__7669;
    wire N__7666;
    wire N__7663;
    wire N__7660;
    wire N__7657;
    wire N__7654;
    wire N__7653;
    wire N__7652;
    wire N__7649;
    wire N__7648;
    wire N__7647;
    wire N__7646;
    wire N__7643;
    wire N__7640;
    wire N__7631;
    wire N__7628;
    wire N__7621;
    wire N__7618;
    wire N__7617;
    wire N__7616;
    wire N__7613;
    wire N__7612;
    wire N__7611;
    wire N__7608;
    wire N__7605;
    wire N__7598;
    wire N__7591;
    wire N__7590;
    wire N__7587;
    wire N__7584;
    wire N__7583;
    wire N__7582;
    wire N__7579;
    wire N__7576;
    wire N__7573;
    wire N__7570;
    wire N__7563;
    wire N__7560;
    wire N__7555;
    wire N__7552;
    wire N__7549;
    wire N__7546;
    wire N__7543;
    wire N__7540;
    wire N__7537;
    wire N__7534;
    wire N__7531;
    wire N__7528;
    wire N__7527;
    wire N__7526;
    wire N__7523;
    wire N__7520;
    wire N__7517;
    wire N__7516;
    wire N__7513;
    wire N__7510;
    wire N__7507;
    wire N__7504;
    wire N__7495;
    wire N__7492;
    wire N__7489;
    wire N__7486;
    wire N__7483;
    wire N__7480;
    wire N__7477;
    wire N__7474;
    wire N__7471;
    wire N__7468;
    wire N__7465;
    wire N__7462;
    wire N__7459;
    wire N__7456;
    wire N__7455;
    wire N__7452;
    wire N__7449;
    wire N__7448;
    wire N__7445;
    wire N__7442;
    wire N__7439;
    wire N__7438;
    wire N__7433;
    wire N__7430;
    wire N__7427;
    wire N__7420;
    wire N__7417;
    wire N__7414;
    wire N__7413;
    wire N__7412;
    wire N__7409;
    wire N__7406;
    wire N__7403;
    wire N__7400;
    wire N__7397;
    wire N__7394;
    wire N__7393;
    wire N__7390;
    wire N__7387;
    wire N__7384;
    wire N__7381;
    wire N__7372;
    wire N__7371;
    wire N__7370;
    wire N__7367;
    wire N__7364;
    wire N__7361;
    wire N__7360;
    wire N__7357;
    wire N__7354;
    wire N__7351;
    wire N__7348;
    wire N__7339;
    wire N__7336;
    wire N__7333;
    wire N__7330;
    wire N__7329;
    wire N__7326;
    wire N__7323;
    wire N__7322;
    wire N__7319;
    wire N__7316;
    wire N__7313;
    wire N__7312;
    wire N__7309;
    wire N__7304;
    wire N__7301;
    wire N__7294;
    wire N__7291;
    wire N__7290;
    wire N__7289;
    wire N__7286;
    wire N__7283;
    wire N__7280;
    wire N__7279;
    wire N__7276;
    wire N__7273;
    wire N__7270;
    wire N__7267;
    wire N__7258;
    wire N__7255;
    wire N__7252;
    wire N__7249;
    wire N__7246;
    wire N__7245;
    wire N__7242;
    wire N__7241;
    wire N__7238;
    wire N__7237;
    wire N__7234;
    wire N__7231;
    wire N__7228;
    wire N__7225;
    wire N__7220;
    wire N__7215;
    wire N__7214;
    wire N__7211;
    wire N__7208;
    wire N__7205;
    wire N__7198;
    wire N__7195;
    wire N__7194;
    wire N__7193;
    wire N__7192;
    wire N__7189;
    wire N__7186;
    wire N__7183;
    wire N__7180;
    wire N__7173;
    wire N__7170;
    wire N__7167;
    wire N__7164;
    wire N__7159;
    wire N__7158;
    wire N__7155;
    wire N__7152;
    wire N__7151;
    wire N__7150;
    wire N__7145;
    wire N__7142;
    wire N__7139;
    wire N__7134;
    wire N__7131;
    wire N__7130;
    wire N__7127;
    wire N__7124;
    wire N__7121;
    wire N__7114;
    wire N__7113;
    wire N__7110;
    wire N__7107;
    wire N__7106;
    wire N__7105;
    wire N__7100;
    wire N__7097;
    wire N__7094;
    wire N__7089;
    wire N__7086;
    wire N__7085;
    wire N__7082;
    wire N__7079;
    wire N__7076;
    wire N__7069;
    wire N__7068;
    wire N__7065;
    wire N__7062;
    wire N__7061;
    wire N__7058;
    wire N__7055;
    wire N__7052;
    wire N__7051;
    wire N__7044;
    wire N__7041;
    wire N__7040;
    wire N__7037;
    wire N__7034;
    wire N__7031;
    wire N__7024;
    wire N__7023;
    wire N__7022;
    wire N__7019;
    wire N__7016;
    wire N__7013;
    wire N__7012;
    wire N__7007;
    wire N__7004;
    wire N__7001;
    wire N__7000;
    wire N__6997;
    wire N__6992;
    wire N__6989;
    wire N__6982;
    wire N__6979;
    wire N__6976;
    wire N__6973;
    wire N__6972;
    wire N__6967;
    wire N__6964;
    wire N__6961;
    wire N__6958;
    wire N__6955;
    wire N__6952;
    wire N__6949;
    wire N__6946;
    wire N__6943;
    wire N__6940;
    wire N__6937;
    wire N__6936;
    wire N__6933;
    wire N__6930;
    wire N__6925;
    wire N__6922;
    wire N__6919;
    wire N__6916;
    wire N__6913;
    wire N__6910;
    wire N__6907;
    wire N__6904;
    wire N__6901;
    wire N__6900;
    wire N__6897;
    wire N__6894;
    wire N__6889;
    wire N__6886;
    wire N__6883;
    wire N__6880;
    wire N__6877;
    wire N__6876;
    wire N__6875;
    wire N__6868;
    wire N__6865;
    wire N__6862;
    wire N__6859;
    wire N__6856;
    wire N__6855;
    wire N__6854;
    wire N__6851;
    wire N__6848;
    wire N__6845;
    wire N__6840;
    wire N__6835;
    wire N__6832;
    wire N__6829;
    wire N__6826;
    wire N__6823;
    wire N__6820;
    wire N__6817;
    wire N__6814;
    wire N__6811;
    wire N__6810;
    wire N__6807;
    wire N__6806;
    wire N__6803;
    wire N__6802;
    wire N__6797;
    wire N__6794;
    wire N__6791;
    wire N__6784;
    wire N__6783;
    wire N__6782;
    wire N__6779;
    wire N__6778;
    wire N__6777;
    wire N__6776;
    wire N__6773;
    wire N__6770;
    wire N__6767;
    wire N__6764;
    wire N__6757;
    wire N__6748;
    wire N__6745;
    wire N__6744;
    wire N__6743;
    wire N__6742;
    wire N__6741;
    wire N__6738;
    wire N__6735;
    wire N__6728;
    wire N__6721;
    wire N__6718;
    wire N__6715;
    wire N__6712;
    wire N__6709;
    wire N__6706;
    wire N__6703;
    wire N__6700;
    wire N__6697;
    wire N__6694;
    wire N__6691;
    wire N__6690;
    wire N__6689;
    wire N__6686;
    wire N__6683;
    wire N__6682;
    wire N__6679;
    wire N__6674;
    wire N__6671;
    wire N__6668;
    wire N__6665;
    wire N__6660;
    wire N__6655;
    wire N__6652;
    wire N__6649;
    wire N__6646;
    wire N__6643;
    wire N__6640;
    wire N__6639;
    wire N__6636;
    wire N__6633;
    wire N__6630;
    wire N__6625;
    wire N__6622;
    wire N__6619;
    wire N__6618;
    wire N__6617;
    wire N__6614;
    wire N__6613;
    wire N__6610;
    wire N__6607;
    wire N__6604;
    wire N__6601;
    wire N__6598;
    wire N__6595;
    wire N__6594;
    wire N__6591;
    wire N__6588;
    wire N__6583;
    wire N__6580;
    wire N__6571;
    wire N__6570;
    wire N__6567;
    wire N__6564;
    wire N__6559;
    wire N__6556;
    wire N__6553;
    wire N__6552;
    wire N__6549;
    wire N__6546;
    wire N__6541;
    wire N__6538;
    wire N__6535;
    wire N__6532;
    wire N__6529;
    wire N__6526;
    wire N__6523;
    wire N__6520;
    wire N__6517;
    wire N__6514;
    wire N__6511;
    wire N__6508;
    wire N__6505;
    wire N__6502;
    wire N__6501;
    wire N__6500;
    wire N__6497;
    wire N__6494;
    wire N__6491;
    wire N__6484;
    wire N__6483;
    wire N__6480;
    wire N__6477;
    wire N__6472;
    wire N__6469;
    wire N__6468;
    wire N__6465;
    wire N__6462;
    wire N__6459;
    wire N__6454;
    wire N__6451;
    wire N__6450;
    wire N__6447;
    wire N__6444;
    wire N__6441;
    wire N__6438;
    wire N__6433;
    wire N__6430;
    wire N__6427;
    wire N__6424;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire N__6412;
    wire N__6409;
    wire N__6406;
    wire N__6403;
    wire N__6400;
    wire N__6397;
    wire N__6394;
    wire N__6391;
    wire N__6388;
    wire N__6387;
    wire N__6382;
    wire N__6379;
    wire N__6376;
    wire N__6375;
    wire N__6372;
    wire N__6369;
    wire N__6368;
    wire N__6367;
    wire N__6362;
    wire N__6361;
    wire N__6360;
    wire N__6359;
    wire N__6358;
    wire N__6357;
    wire N__6354;
    wire N__6351;
    wire N__6348;
    wire N__6337;
    wire N__6328;
    wire N__6327;
    wire N__6326;
    wire N__6325;
    wire N__6324;
    wire N__6321;
    wire N__6318;
    wire N__6317;
    wire N__6316;
    wire N__6313;
    wire N__6308;
    wire N__6299;
    wire N__6292;
    wire N__6289;
    wire N__6286;
    wire N__6283;
    wire N__6280;
    wire N__6277;
    wire N__6274;
    wire N__6271;
    wire N__6268;
    wire N__6267;
    wire N__6264;
    wire N__6261;
    wire N__6258;
    wire N__6253;
    wire N__6250;
    wire N__6247;
    wire N__6244;
    wire N__6241;
    wire N__6238;
    wire N__6235;
    wire N__6232;
    wire N__6229;
    wire N__6226;
    wire N__6223;
    wire N__6220;
    wire N__6217;
    wire N__6214;
    wire N__6211;
    wire N__6208;
    wire N__6205;
    wire N__6202;
    wire N__6199;
    wire N__6196;
    wire N__6193;
    wire N__6190;
    wire N__6187;
    wire N__6184;
    wire N__6181;
    wire N__6178;
    wire N__6175;
    wire N__6172;
    wire N__6169;
    wire N__6166;
    wire N__6163;
    wire N__6160;
    wire N__6157;
    wire N__6154;
    wire N__6151;
    wire N__6150;
    wire N__6147;
    wire N__6144;
    wire N__6139;
    wire N__6136;
    wire N__6133;
    wire N__6130;
    wire N__6127;
    wire N__6124;
    wire N__6121;
    wire N__6118;
    wire N__6115;
    wire N__6114;
    wire N__6113;
    wire N__6110;
    wire N__6107;
    wire N__6104;
    wire N__6103;
    wire N__6102;
    wire N__6097;
    wire N__6094;
    wire N__6091;
    wire N__6088;
    wire N__6085;
    wire N__6078;
    wire N__6073;
    wire N__6070;
    wire N__6067;
    wire N__6064;
    wire N__6061;
    wire N__6058;
    wire N__6055;
    wire N__6052;
    wire N__6049;
    wire N__6046;
    wire N__6043;
    wire N__6040;
    wire N__6037;
    wire N__6034;
    wire N__6031;
    wire N__6028;
    wire N__6025;
    wire N__6022;
    wire N__6019;
    wire N__6016;
    wire N__6015;
    wire N__6014;
    wire N__6013;
    wire N__6012;
    wire N__6011;
    wire N__6010;
    wire N__6009;
    wire N__6002;
    wire N__5991;
    wire N__5986;
    wire N__5983;
    wire N__5980;
    wire N__5977;
    wire N__5974;
    wire N__5971;
    wire N__5968;
    wire N__5965;
    wire N__5962;
    wire N__5959;
    wire N__5956;
    wire N__5955;
    wire N__5954;
    wire N__5953;
    wire N__5950;
    wire N__5949;
    wire N__5948;
    wire N__5947;
    wire N__5946;
    wire N__5945;
    wire N__5944;
    wire N__5943;
    wire N__5942;
    wire N__5941;
    wire N__5938;
    wire N__5933;
    wire N__5930;
    wire N__5925;
    wire N__5920;
    wire N__5915;
    wire N__5908;
    wire N__5903;
    wire N__5900;
    wire N__5887;
    wire N__5886;
    wire N__5885;
    wire N__5882;
    wire N__5881;
    wire N__5880;
    wire N__5879;
    wire N__5878;
    wire N__5877;
    wire N__5876;
    wire N__5875;
    wire N__5874;
    wire N__5871;
    wire N__5870;
    wire N__5869;
    wire N__5866;
    wire N__5865;
    wire N__5862;
    wire N__5861;
    wire N__5858;
    wire N__5855;
    wire N__5854;
    wire N__5853;
    wire N__5852;
    wire N__5851;
    wire N__5848;
    wire N__5847;
    wire N__5844;
    wire N__5841;
    wire N__5838;
    wire N__5831;
    wire N__5822;
    wire N__5819;
    wire N__5814;
    wire N__5811;
    wire N__5800;
    wire N__5793;
    wire N__5790;
    wire N__5787;
    wire N__5784;
    wire N__5767;
    wire N__5764;
    wire N__5761;
    wire N__5758;
    wire N__5755;
    wire N__5752;
    wire N__5749;
    wire N__5746;
    wire N__5743;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5731;
    wire N__5728;
    wire N__5725;
    wire N__5722;
    wire N__5719;
    wire N__5718;
    wire N__5715;
    wire N__5712;
    wire N__5709;
    wire N__5706;
    wire N__5701;
    wire N__5698;
    wire N__5695;
    wire N__5692;
    wire N__5689;
    wire N__5686;
    wire N__5683;
    wire N__5680;
    wire N__5677;
    wire N__5674;
    wire N__5671;
    wire N__5670;
    wire N__5665;
    wire N__5664;
    wire N__5663;
    wire N__5662;
    wire N__5661;
    wire N__5658;
    wire N__5653;
    wire N__5650;
    wire N__5647;
    wire N__5642;
    wire N__5635;
    wire N__5634;
    wire N__5629;
    wire N__5628;
    wire N__5625;
    wire N__5624;
    wire N__5623;
    wire N__5622;
    wire N__5621;
    wire N__5618;
    wire N__5615;
    wire N__5610;
    wire N__5605;
    wire N__5596;
    wire N__5595;
    wire N__5592;
    wire N__5591;
    wire N__5590;
    wire N__5589;
    wire N__5586;
    wire N__5583;
    wire N__5580;
    wire N__5575;
    wire N__5566;
    wire N__5565;
    wire N__5564;
    wire N__5563;
    wire N__5556;
    wire N__5555;
    wire N__5552;
    wire N__5549;
    wire N__5546;
    wire N__5543;
    wire N__5540;
    wire N__5537;
    wire N__5530;
    wire N__5527;
    wire N__5524;
    wire N__5521;
    wire N__5518;
    wire N__5515;
    wire N__5512;
    wire N__5509;
    wire N__5506;
    wire N__5503;
    wire N__5500;
    wire N__5497;
    wire N__5494;
    wire N__5491;
    wire N__5488;
    wire N__5485;
    wire N__5482;
    wire N__5479;
    wire N__5476;
    wire N__5473;
    wire N__5470;
    wire N__5467;
    wire N__5464;
    wire N__5461;
    wire N__5458;
    wire N__5455;
    wire N__5452;
    wire N__5449;
    wire N__5446;
    wire N__5443;
    wire N__5440;
    wire N__5437;
    wire N__5434;
    wire N__5431;
    wire N__5428;
    wire N__5425;
    wire N__5422;
    wire N__5419;
    wire N__5416;
    wire N__5413;
    wire N__5410;
    wire N__5407;
    wire N__5404;
    wire N__5401;
    wire N__5398;
    wire N__5395;
    wire N__5392;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5371;
    wire N__5368;
    wire N__5365;
    wire N__5362;
    wire N__5359;
    wire N__5356;
    wire N__5353;
    wire N__5350;
    wire N__5347;
    wire N__5344;
    wire N__5341;
    wire N__5338;
    wire N__5335;
    wire N__5332;
    wire N__5329;
    wire N__5326;
    wire N__5323;
    wire N__5320;
    wire N__5317;
    wire N__5316;
    wire N__5313;
    wire N__5310;
    wire N__5305;
    wire N__5302;
    wire N__5301;
    wire N__5298;
    wire N__5295;
    wire N__5290;
    wire N__5287;
    wire N__5284;
    wire N__5281;
    wire N__5278;
    wire N__5275;
    wire N__5272;
    wire N__5269;
    wire N__5266;
    wire N__5263;
    wire N__5260;
    wire N__5257;
    wire N__5254;
    wire N__5251;
    wire N__5248;
    wire N__5245;
    wire N__5242;
    wire N__5239;
    wire N__5236;
    wire N__5233;
    wire N__5230;
    wire N__5227;
    wire N__5224;
    wire N__5221;
    wire N__5218;
    wire N__5215;
    wire N__5212;
    wire N__5209;
    wire N__5206;
    wire N__5203;
    wire N__5200;
    wire N__5197;
    wire N__5194;
    wire N__5191;
    wire N__5188;
    wire N__5185;
    wire N__5182;
    wire N__5179;
    wire N__5176;
    wire N__5173;
    wire N__5170;
    wire N__5167;
    wire N__5164;
    wire N__5161;
    wire N__5158;
    wire N__5155;
    wire N__5152;
    wire N__5149;
    wire N__5146;
    wire N__5143;
    wire N__5140;
    wire N__5137;
    wire N__5134;
    wire N__5131;
    wire N__5128;
    wire N__5125;
    wire N__5122;
    wire N__5119;
    wire N__5116;
    wire N__5113;
    wire N__5110;
    wire N__5107;
    wire N__5104;
    wire N__5101;
    wire N__5098;
    wire N__5095;
    wire N__5092;
    wire N__5089;
    wire N__5086;
    wire N__5083;
    wire N__5080;
    wire N__5077;
    wire BTN_N_c;
    wire VCCG0;
    wire GNDG0;
    wire \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_0 ;
    wire bfn_12_4_0_;
    wire \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0 ;
    wire \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1 ;
    wire un1_oRxFlag_0_i_cascade_;
    wire \DUT.fifo_rx_inst.rFifoCount_RNITA8H2Z0Z_1 ;
    wire rFifoCount_RNIHH0D1_0_cascade_;
    wire \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0 ;
    wire ioFifoData_in_6;
    wire ioFifoData_in_0;
    wire ioFifoData_in_4;
    wire wRxFifoData_0;
    wire \DUT.rFifoDatarx_0 ;
    wire wRxFifoData_4;
    wire wRxFifoData_6;
    wire \DUT.rFifoDatarx_6 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_7 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_7 ;
    wire \DUT.fifo_rx_inst.rFifoDataro_0 ;
    wire \DUT.fifo_rx_inst.rFifoDataro_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_6 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_7 ;
    wire \DUT.fifo_rx_inst.rReadPtr_RNIDU4H2Z0Z_0_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_6 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6 ;
    wire \DUT.fifo_rx_inst.rReadPtr_RNIDU4H2Z0Z_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_4 ;
    wire \DUT.rFifoDatarx_0_4 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_5 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_5 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_6 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_4 ;
    wire wPllLocked_i;
    wire \DUT.uart_inst0.N_275_cascade_ ;
    wire \DUT.uart_inst0.g0_0_5_cascade_ ;
    wire \DUT.uart_inst0.g0_6_cascade_ ;
    wire \DUT.uart_inst0.g0_1_0 ;
    wire \DUT.uart_inst0.g3_0_cascade_ ;
    wire \DUT.uart_inst0.g0_0_4 ;
    wire \DUT.fifo_rx_inst.rFifoCountZ0Z_1 ;
    wire \DUT.fifo_rx_inst.N_148 ;
    wire ioFifoData_in_7;
    wire ioFifoData_in_1;
    wire ioFifoData_in_3;
    wire ioFifoData_in_5;
    wire ioFifoData_in_2;
    wire wRxFifoData_1;
    wire wRxFifoData_2;
    wire wRxFifoData_3;
    wire \DUT.rFifoDatarx_0_5 ;
    wire wRxFifoData_5;
    wire \DUT.rFifoDatarx_0_7 ;
    wire wRxFifoData_7;
    wire un1_oRxFlag_0_i_0;
    wire \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1 ;
    wire \DUT.rFifoDatarx_0_1 ;
    wire \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1 ;
    wire \DUT.wRcvd ;
    wire \DUT.fifo_rx_inst.rFifoCountZ0Z_2 ;
    wire \DUT.fifo_rx_inst.N_194_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_2 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_2 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2_cascade_ ;
    wire \DUT.rFifoDatarx_0_2 ;
    wire \DUT.rFifoDataror_0_0_cascade_ ;
    wire \DUT.rFifoDataror_1 ;
    wire \DUT.uart_inst0.N_257 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_3 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_3 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ;
    wire \DUT.rFifoDatarx_3 ;
    wire \DUT.fifo_rx_inst.rReadPtrZ0Z_0 ;
    wire \DUT.fifo_rx_inst.rReadPtrZ0Z_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_2 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_3 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_4 ;
    wire \DUT.fifo_rx_inst.rFifoData_awe0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_2 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_5 ;
    wire \DUT.uart_inst0.rx_clk_divider_5_i_a2_1_3 ;
    wire \DUT.uart_inst0.N_222_cascade_ ;
    wire \DUT.uart_inst0.rx_clk_divider_5_i_a2_11_0_5_cascade_ ;
    wire \DUT.uart_inst0.rx_clk_divider_5_i_a2_11_5 ;
    wire \DUT.uart_inst0.rx_clk_divider_5_i_a2_11_5_cascade_ ;
    wire \DUT.uart_inst0.N_221 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_0_0_c_RNOZ0 ;
    wire bfn_14_3_0_;
    wire \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_0Z0Z_0 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_0 ;
    wire \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_1Z0Z_0 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_1 ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_3 ;
    wire \DUT.uart_inst0.rx_clk_divider_RNIP8N2BZ0Z_0 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_2 ;
    wire \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_2Z0Z_0 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_3 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_4 ;
    wire \DUT.uart_inst0.rx_countdown_3_5_cascade_ ;
    wire \DUT.uart_inst0.g3_4 ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_0 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_i_3 ;
    wire \DUT.uart_inst0.N_275 ;
    wire \DUT.uart_inst0.N_196_cascade_ ;
    wire \DUT.uart_inst0.N_33_cascade_ ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_3_0_c_RNIP8IZ0Z482 ;
    wire \DUT.uart_inst0.rx_bits_remaining_RNO_0Z0Z_1 ;
    wire \DUT.uart_inst0.g0_8_1 ;
    wire P1A2_c_0_0;
    wire \DUT.uart_inst0.recv_stateZ0Z_4 ;
    wire \fifo_inst.ftdi_output_inst.rFifoState_0_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_6 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_7 ;
    wire \DUT.fifo_rx_inst.rFifoData_awe3 ;
    wire \DUT.fifo_rx_inst.rFifoDataro_3 ;
    wire \DUT.fifo_rx_inst.rFifoData_awe2 ;
    wire \DUT.fifo_rx_inst.rFifoDataro_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_awe1 ;
    wire \DUT.fifo_tx_inst.rFifoData_awe3_cascade_ ;
    wire \DUT.fifo_tx_inst.un1_i11_i ;
    wire \DUT.fifo_tx_inst.un1_i11_i_cascade_ ;
    wire \DUT.fifo_rx_inst.N_194 ;
    wire \DUT.fifo_rx_inst.rWritePtrZ0Z_0 ;
    wire \DUT.fifo_rx_inst.rWritePtrZ0Z_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_5 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_3 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_4 ;
    wire \DUT.fifo_rx_inst.rFifoData_awe1 ;
    wire bfn_15_1_0_;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_0 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_1 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_3 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_3 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_2 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_4 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_4 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_3 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_5 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_5 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_4 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_6 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_6 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_5 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_7 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_6 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_7 ;
    wire bfn_15_2_0_;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_8 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_9 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_10 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_11 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_12 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_14 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_13 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_15 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_15 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_14 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_15 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_16 ;
    wire bfn_15_3_0_;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_16 ;
    wire \DUT.uart_inst0.recv_state_RNO_2Z0Z_4_cascade_ ;
    wire \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa_0_a2_0_a2_0_a3_1 ;
    wire \DUT.uart_inst0.rx_countdown_8_i_0_o2_1_2_2_cascade_ ;
    wire \DUT.uart_inst0.recv_state_ns_0_i_0_0_o2_0_3 ;
    wire \DUT.uart_inst0.G_9_1_cascade_ ;
    wire \DUT.uart_inst0.G_11_i_a4_0_4 ;
    wire \DUT.uart_inst0.N_4_i_1 ;
    wire \DUT.wRxByte_1 ;
    wire \DUT.wRxByte_0 ;
    wire \DUT.wRxByte_4 ;
    wire \DUT.wRxByte_5 ;
    wire \DUT.wRxByte_6 ;
    wire \DUT.wRxByte_7 ;
    wire \DUT.fifo_tx_inst.rFifoData_awe3 ;
    wire rTxByteZ0Z_0;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_0 ;
    wire rTxByteZ0Z_1;
    wire rTxByteZ0Z_3;
    wire rTxByteZ0Z_6;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_4 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_4 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_ ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_4 ;
    wire rTxByteZ0Z_4;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_4 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_5 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_5 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_5 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ;
    wire rTxByteZ0Z_5;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_5 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_6 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_6 ;
    wire \DUT.fifo_tx_inst.rFifoDataro_3 ;
    wire \DUT.fifo_tx_inst.rFifoDataro_0 ;
    wire \DUT.fifo_tx_inst.rFifoDataro_1 ;
    wire \DUT.rFifoDataror_0_0_0 ;
    wire \DUT.rFifoDataror_1_0_cascade_ ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_6 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_6 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6 ;
    wire \DUT.fifo_tx_inst.rWritePtrZ0Z_0 ;
    wire \DUT.fifo_tx_inst.N_79_cascade_ ;
    wire \DUT.fifo_tx_inst.rWritePtrZ0Z_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_awe2 ;
    wire \DUT.fifo_tx_inst.rFifoDataro_2 ;
    wire \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4 ;
    wire \fifo_inst.ftdi_output_inst.rWrDelayZ0 ;
    wire \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_3 ;
    wire P1A4_c;
    wire rTxBusReady;
    wire \DUT.uart_inst0.rx_clk_divider_1_8 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_8 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_9 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_9 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_11 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_11 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_12 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_12 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_1 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_7 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_1 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ1Z_1 ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_5 ;
    wire \DUT.uart_inst0.rx_countdown_3_1 ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_1 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_2 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_2 ;
    wire \DUT.uart_inst0.g0_0_3 ;
    wire \DUT.uart_inst0.g1 ;
    wire \DUT.uart_inst0.g0_0_0 ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_2 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_17 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_17 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_10 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_10 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_13 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_13 ;
    wire \DUT.uart_inst0.N_199_0 ;
    wire N_1239_i;
    wire \DUT.uart_inst0.recv_stateZ0Z_0 ;
    wire \DUT.uart_inst0.rx_clk_divider_5_i_a2_12_1_5 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_16 ;
    wire \DUT.uart_inst0.rx_clk_divider_5_i_a2_12_4_5 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_14 ;
    wire \DUT.uart_inst0.rx_clk_divider_5_i_a2_12_5 ;
    wire \DUT.uart_inst0.N_31_0 ;
    wire \DUT.uart_inst0.N_203 ;
    wire \DUT.uart_inst0.recv_state_ns_0_i_0_0_a3_0_0_3 ;
    wire \DUT.uart_inst0.rx_bits_remainingZ0Z_2 ;
    wire \DUT.uart_inst0.rx_bits_remainingZ0Z_1 ;
    wire \DUT.uart_inst0.rx_bits_remainingZ0Z_3 ;
    wire \DUT.uart_inst0.rx_bits_remainingZ0Z_0 ;
    wire \DUT.uart_inst0.N_215_4 ;
    wire \DUT.uart_inst0.N_215_4_cascade_ ;
    wire \DUT.uart_inst0.recv_state_srsts_1_2_cascade_ ;
    wire \DUT.uart_inst0.N_193 ;
    wire \DUT.uart_inst0.recv_stateZ0Z_2 ;
    wire \DUT.uart_inst0.g0_0 ;
    wire \DUT.wRxByte_3 ;
    wire \DUT.wRxByte_2 ;
    wire \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_3 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_3 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_3 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_3 ;
    wire \DUT.rFifoDatarx_0_0 ;
    wire \DUT.uart_inst0.tx_out_6_iv_0_1 ;
    wire \DUT.rFifoDatarx_1 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_1 ;
    wire \DUT.rFifoDatarx_2 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_2 ;
    wire \DUT.rFifoDatarx_0_3 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_3 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_7 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_7 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_ ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_7 ;
    wire \DUT.uart_inst0.tx_out_6_iv_0_a3_0_1 ;
    wire \DUT.uart_inst0.N_101 ;
    wire \DUT.rFifoDatarx_5 ;
    wire \DUT.rFifoDatarx_0_6 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_6 ;
    wire \DUT.rFifoDatarx_4 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_5 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_4 ;
    wire \DUT.rFifoDatarx_7 ;
    wire \DUT.uart_inst0.N_145 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_7 ;
    wire \DUT.uart_inst0.N_22_i ;
    wire \DUT.fifo_tx_inst.N_83_cascade_ ;
    wire \DUT.uart_inst0.tx_dataZ0Z_0 ;
    wire P1A7_c;
    wire \DUT.uart_inst0.N_98 ;
    wire \fifo_inst.ftdi_output_inst.rFifoStatec_0 ;
    wire \DUT.fifo_tx_inst.N_79 ;
    wire \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0 ;
    wire \DUT.fifo_tx_inst.rFifoCountZ0Z_0 ;
    wire bfn_16_11_0_;
    wire \DUT.fifo_tx_inst.rFifoCount_RNISSQ21Z0Z_1 ;
    wire \DUT.fifo_tx_inst.rFifoCountZ0Z_1 ;
    wire \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0 ;
    wire \DUT.fifo_tx_inst.N_83 ;
    wire \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1 ;
    wire \DUT.fifo_tx_inst.rFifoCountZ0Z_2 ;
    wire P1A1_c;
    wire \DUT.uart_inst0.recv_stateZ0Z_3 ;
    wire \DUT.uart_inst0.g0_1 ;
    wire \DUT.uart_inst0.recv_stateZ0Z_5 ;
    wire \DUT.uart_inst0.rx_countdown_3_4 ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_4 ;
    wire \DUT.uart_inst0.rx_countdown_3_5 ;
    wire \DUT.uart_inst0.recv_state_RNO_2Z0Z_1 ;
    wire \DUT.uart_inst0.rx_countdown_3_0 ;
    wire \DUT.uart_inst0.rx_countdown_3_2 ;
    wire \DUT.uart_inst0.G_10_i_a4_0_4_cascade_ ;
    wire \DUT.uart_inst0.rx_countdown_3_3 ;
    wire \DUT.uart_inst0.N_4_i_0_1_cascade_ ;
    wire \DUT.uart_inst0.N_149 ;
    wire \DUT.uart_inst0.recv_stateZ0Z_1 ;
    wire rRxReadZ0;
    wire \DUT.fifo_rx_inst.N_206 ;
    wire \DUT.fifo_rx_inst.rFifoCountZ0Z_0 ;
    wire \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1 ;
    wire P1A2_c;
    wire rFifoCount_RNIHH0D1_0;
    wire rTxWriteZ0;
    wire P1A3_c;
    wire rTxByteZ0Z_2;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_2 ;
    wire rTxByteZ0Z_7;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_7 ;
    wire \DUT.fifo_tx_inst.rFifoData_awe0 ;
    wire \DUT.uart_inst0.tx_bits_remainingZ0Z_2 ;
    wire \DUT.uart_inst0.tx_bits_remainingZ0Z_1 ;
    wire \DUT.uart_inst0.tx_bits_remainingZ0Z_0 ;
    wire \DUT.uart_inst0.N_142_cascade_ ;
    wire wPllLocked;
    wire \DUT.uart_inst0.N_84_cascade_ ;
    wire \DUT.uart_inst0.N_22 ;
    wire \DUT.uart_inst0.N_22_cascade_ ;
    wire \DUT.uart_inst0.un1_tx_bits_remaining_c3 ;
    wire \DUT.uart_inst0.tx_bits_remainingZ0Z_3 ;
    wire \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2 ;
    wire \fifo_inst.ftdi_output_inst.N_78_cascade_ ;
    wire \DUT.uart_inst0.N_142 ;
    wire \DUT.uart_inst0.N_144 ;
    wire \DUT.uart_inst0.N_74_cascade_ ;
    wire \DUT.uart_inst0.N_143 ;
    wire \DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0_cascade_ ;
    wire \DUT.uart_inst0.N_75 ;
    wire \DUT.uart_inst0.N_75_cascade_ ;
    wire \DUT.uart_inst0.tx_countdown_7s2_0_0 ;
    wire \DUT.uart_inst0.tx_state_ns_i_i_o2_a0_3_0_cascade_ ;
    wire \DUT.uart_inst0.N_69_i ;
    wire \DUT.uart_inst0.tx_countdown_30_3_cascade_ ;
    wire \DUT.uart_inst0.N_84 ;
    wire \DUT.uart_inst0.N_30_1 ;
    wire N_1242_i;
    wire N_1240_i;
    wire rTxBusReady_rep1_i_ess;
    wire rTxBusReady_rep3_i_ess;
    wire rTxBusReady_rep0_i_ess;
    wire iTxE_n_c;
    wire \fifo_inst.ftdi_output_inst.N_68_0 ;
    wire wPllLocked_i_g;
    wire \fifo_inst.ftdi_output_inst.un1_oTx_n_1_sqmuxa_0_i_cascade_ ;
    wire \fifo_inst.ftdi_output_inst.un1_oTx_n_1_sqmuxa_0_i_0 ;
    wire iRxF_n_c;
    wire \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0 ;
    wire \fifo_inst.ftdi_output_inst.N_80 ;
    wire \DUT.uart_inst0.N_77_cascade_ ;
    wire \DUT.uart_inst0.tx_state_RNI8CH01Z0Z_1 ;
    wire \DUT.uart_inst0.tx_state_RNI8CH01Z0Z_1_cascade_ ;
    wire \DUT.uart_inst0.N_59_i ;
    wire \DUT.N_93 ;
    wire \DUT.tx_state_1 ;
    wire \DUT.rTransmitZ0 ;
    wire \DUT.fifo_tx_inst.rReadPtrZ0Z_1 ;
    wire \DUT.fifo_tx_inst.un1_i11_2_i ;
    wire \DUT.fifo_tx_inst.rReadPtr11 ;
    wire \DUT.fifo_tx_inst.un1_i11_2_i_cascade_ ;
    wire \DUT.fifo_tx_inst.rReadPtrZ0Z_0 ;
    wire \DUT.uart_inst0.N_74 ;
    wire \DUT.tx_state_0 ;
    wire \DUT.uart_inst0.tx_countdown_7_1_2 ;
    wire \DUT.uart_inst0.N_91 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_2 ;
    wire \DUT.uart_inst0.tx_countdown_0_c4_cascade_ ;
    wire \DUT.uart_inst0.tx_countdown_7_ns_1_4 ;
    wire \DUT.uart_inst0.tx_countdown_7_ns_1_1_cascade_ ;
    wire \DUT.uart_inst0.tx_countdown_0_c4 ;
    wire \DUT.uart_inst0.tx_countdown_7_ns_1_5 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_0 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_1 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_5 ;
    wire \DUT.uart_inst0.tx_countdown_7_m1_0_o2_1_2_cascade_ ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_4 ;
    wire \DUT.uart_inst0.N_68 ;
    wire \DUT.uart_inst0.N_146 ;
    wire \DUT.uart_inst0.tx_countdown_7_sm0_0 ;
    wire \DUT.uart_inst0.tx_countdown_7_ns_1_3 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_3 ;
    wire rTxBusReady_rep2_i_ess;
    wire N_1241_i;
    wire \DUT.uart_inst0.un1_tx_clk_divider_9 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_6_cascade_ ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_0_cascade_ ;
    wire wPllLocked_g;
    wire \DUT.uart_inst0.un1_tx_clk_divider_8 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_7 ;
    wire \DUT.uart_inst0.N_77 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_0 ;
    wire \DUT.uart_inst0.N_147 ;
    wire bfn_21_9_0_;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_1 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_0 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_2 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_1 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_3 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_2 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_4 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_3 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_5 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_4 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_6 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_5 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_7 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_6 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_7 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_8 ;
    wire bfn_21_10_0_;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_9 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_8 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_10 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_9 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_11 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_10 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_12 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_11 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_12 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_13 ;
    wire CONSTANT_ONE_NET;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_0 ;
    wire _gnd_net_;
    wire clk_48mhz;
    wire \DUT.uart_inst0.N_20 ;

    defparam \top_pll_inst.top_pll_inst_pll .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \top_pll_inst.top_pll_inst_pll .TEST_MODE=1'b0;
    defparam \top_pll_inst.top_pll_inst_pll .SHIFTREG_DIV_MODE=2'b00;
    defparam \top_pll_inst.top_pll_inst_pll .PLLOUT_SELECT="GENCLK";
    defparam \top_pll_inst.top_pll_inst_pll .FILTER_RANGE=3'b001;
    defparam \top_pll_inst.top_pll_inst_pll .FEEDBACK_PATH="SIMPLE";
    defparam \top_pll_inst.top_pll_inst_pll .FDA_RELATIVE=4'b0000;
    defparam \top_pll_inst.top_pll_inst_pll .FDA_FEEDBACK=4'b0000;
    defparam \top_pll_inst.top_pll_inst_pll .ENABLE_ICEGATE=1'b0;
    defparam \top_pll_inst.top_pll_inst_pll .DIVR=4'b0000;
    defparam \top_pll_inst.top_pll_inst_pll .DIVQ=3'b100;
    defparam \top_pll_inst.top_pll_inst_pll .DIVF=7'b0111111;
    defparam \top_pll_inst.top_pll_inst_pll .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    PLL40 \top_pll_inst.top_pll_inst_pll  (
            .PLLOUTGLOBAL(clk_48mhz),
            .SDI(GNDG0),
            .BYPASS(GNDG0),
            .RESETB(N__5089),
            .PLLOUTCORE(),
            .LOCK(\PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO ),
            .SDO(),
            .SCLK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .EXTFEEDBACK(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLIN(N__13366));
    IO_PAD \top_pll_inst.top_pll_inst_iopad  (
            .OE(VCCG0),
            .DIN(),
            .DOUT(N__13366),
            .PACKAGEPIN(iClk));
    IO_PAD P1A8_obuft_iopad (
            .OE(N__13352),
            .DIN(N__13351),
            .DOUT(N__13350),
            .PACKAGEPIN(P1A8));
    defparam P1A8_obuft_preio.NEG_TRIGGER=1'b0;
    defparam P1A8_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO P1A8_obuft_preio (
            .PADOEN(N__13352),
            .PADOUT(N__13351),
            .PADIN(N__13350),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_6_iopad (
            .OE(N__13343),
            .DIN(N__13342),
            .DOUT(N__13341),
            .PACKAGEPIN(ioFifoData[6]));
    defparam ioFifoData_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_6_preio (
            .PADOEN(N__13343),
            .PADOUT(N__13342),
            .PADIN(N__13341),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7830),
            .DIN0(ioFifoData_in_6),
            .DOUT0(N__12960),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_3_iopad (
            .OE(N__13334),
            .DIN(N__13333),
            .DOUT(N__13332),
            .PACKAGEPIN(ioFifoData[3]));
    defparam ioFifoData_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_3_preio (
            .PADOEN(N__13334),
            .PADOUT(N__13333),
            .PADIN(N__13332),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10819),
            .DIN0(ioFifoData_in_3),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A4_obuf_iopad (
            .OE(N__13325),
            .DIN(N__13324),
            .DOUT(N__13323),
            .PACKAGEPIN(P1A4));
    defparam P1A4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO P1A4_obuf_preio (
            .PADOEN(N__13325),
            .PADOUT(N__13324),
            .PADIN(N__13323),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7873),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD oRx_n_obuf_iopad (
            .OE(N__13316),
            .DIN(N__13315),
            .DOUT(N__13314),
            .PACKAGEPIN(oRx_n));
    defparam oRx_n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam oRx_n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO oRx_n_obuf_preio (
            .PADOEN(N__13316),
            .PADOUT(N__13315),
            .PADIN(N__13314),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10182),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A2_obuf_iopad (
            .OE(N__13307),
            .DIN(N__13306),
            .DOUT(N__13305),
            .PACKAGEPIN(P1A2));
    defparam P1A2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO P1A2_obuf_preio (
            .PADOEN(N__13307),
            .PADOUT(N__13306),
            .PADIN(N__13305),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10351),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_0_iopad (
            .OE(N__13298),
            .DIN(N__13297),
            .DOUT(N__13296),
            .PACKAGEPIN(ioFifoData[0]));
    defparam ioFifoData_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_0_preio (
            .PADOEN(N__13298),
            .PADOUT(N__13297),
            .PADIN(N__13296),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__8296),
            .DIN0(ioFifoData_in_0),
            .DOUT0(N__13041),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD iRxF_n_ibuf_iopad (
            .OE(N__13289),
            .DIN(N__13288),
            .DOUT(N__13287),
            .PACKAGEPIN(iRxF_n));
    defparam iRxF_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam iRxF_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO iRxF_n_ibuf_preio (
            .PADOEN(N__13289),
            .PADOUT(N__13288),
            .PADIN(N__13287),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(iRxF_n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A3_obuf_iopad (
            .OE(N__13280),
            .DIN(N__13279),
            .DOUT(N__13278),
            .PACKAGEPIN(P1A3));
    defparam P1A3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO P1A3_obuf_preio (
            .PADOEN(N__13280),
            .PADOUT(N__13279),
            .PADIN(N__13278),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10195),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A7_obuf_iopad (
            .OE(N__13271),
            .DIN(N__13270),
            .DOUT(N__13269),
            .PACKAGEPIN(P1A7));
    defparam P1A7_obuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A7_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO P1A7_obuf_preio (
            .PADOEN(N__13271),
            .PADOUT(N__13270),
            .PADIN(N__13269),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9060),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_7_iopad (
            .OE(N__13262),
            .DIN(N__13261),
            .DOUT(N__13260),
            .PACKAGEPIN(ioFifoData[7]));
    defparam ioFifoData_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_7_preio (
            .PADOEN(N__13262),
            .PADOUT(N__13261),
            .PADIN(N__13260),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7831),
            .DIN0(ioFifoData_in_7),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BTN_N_ibuf_iopad (
            .OE(N__13253),
            .DIN(N__13252),
            .DOUT(N__13251),
            .PACKAGEPIN(BTN_N));
    defparam BTN_N_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam BTN_N_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO BTN_N_ibuf_preio (
            .PADOEN(N__13253),
            .PADOUT(N__13252),
            .PADIN(N__13251),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(BTN_N_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_4_iopad (
            .OE(N__13244),
            .DIN(N__13243),
            .DOUT(N__13242),
            .PACKAGEPIN(ioFifoData[4]));
    defparam ioFifoData_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_4_preio (
            .PADOEN(N__13244),
            .PADOUT(N__13243),
            .PADIN(N__13242),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7829),
            .DIN0(ioFifoData_in_4),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_1_iopad (
            .OE(N__13235),
            .DIN(N__13234),
            .DOUT(N__13233),
            .PACKAGEPIN(ioFifoData[1]));
    defparam ioFifoData_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_1_preio (
            .PADOEN(N__13235),
            .PADOUT(N__13234),
            .PADIN(N__13233),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10807),
            .DIN0(ioFifoData_in_1),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_5_iopad (
            .OE(N__13226),
            .DIN(N__13225),
            .DOUT(N__13224),
            .PACKAGEPIN(ioFifoData[5]));
    defparam ioFifoData_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_5_preio (
            .PADOEN(N__13226),
            .PADOUT(N__13225),
            .PADIN(N__13224),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__7819),
            .DIN0(ioFifoData_in_5),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD oTx_n_obuf_iopad (
            .OE(N__13217),
            .DIN(N__13216),
            .DOUT(N__13215),
            .PACKAGEPIN(oTx_n));
    defparam oTx_n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam oTx_n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO oTx_n_obuf_preio (
            .PADOEN(N__13217),
            .PADOUT(N__13216),
            .PADIN(N__13215),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7869),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD iTxE_n_ibuf_iopad (
            .OE(N__13208),
            .DIN(N__13207),
            .DOUT(N__13206),
            .PACKAGEPIN(iTxE_n));
    defparam iTxE_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam iTxE_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO iTxE_n_ibuf_preio (
            .PADOEN(N__13208),
            .PADOUT(N__13207),
            .PADIN(N__13206),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(iTxE_n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A1_ibuf_iopad (
            .OE(N__13199),
            .DIN(N__13198),
            .DOUT(N__13197),
            .PACKAGEPIN(P1A1));
    defparam P1A1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO P1A1_ibuf_preio (
            .PADOEN(N__13199),
            .PADOUT(N__13198),
            .PADIN(N__13197),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(P1A1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_2_iopad (
            .OE(N__13190),
            .DIN(N__13189),
            .DOUT(N__13188),
            .PACKAGEPIN(ioFifoData[2]));
    defparam ioFifoData_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_2_preio (
            .PADOEN(N__13190),
            .PADOUT(N__13189),
            .PADIN(N__13188),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__12466),
            .DIN0(ioFifoData_in_2),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A9_obuft_iopad (
            .OE(N__13181),
            .DIN(N__13180),
            .DOUT(N__13179),
            .PACKAGEPIN(P1A9));
    defparam P1A9_obuft_preio.NEG_TRIGGER=1'b0;
    defparam P1A9_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO P1A9_obuft_preio (
            .PADOEN(N__13181),
            .PADOUT(N__13180),
            .PADIN(N__13179),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__3123 (
            .O(N__13162),
            .I(N__13159));
    InMux I__3122 (
            .O(N__13159),
            .I(N__13155));
    InMux I__3121 (
            .O(N__13158),
            .I(N__13152));
    LocalMux I__3120 (
            .O(N__13155),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_9 ));
    LocalMux I__3119 (
            .O(N__13152),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_9 ));
    InMux I__3118 (
            .O(N__13147),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_8 ));
    InMux I__3117 (
            .O(N__13144),
            .I(N__13140));
    InMux I__3116 (
            .O(N__13143),
            .I(N__13137));
    LocalMux I__3115 (
            .O(N__13140),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_10 ));
    LocalMux I__3114 (
            .O(N__13137),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_10 ));
    InMux I__3113 (
            .O(N__13132),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_9 ));
    CascadeMux I__3112 (
            .O(N__13129),
            .I(N__13125));
    CascadeMux I__3111 (
            .O(N__13128),
            .I(N__13122));
    InMux I__3110 (
            .O(N__13125),
            .I(N__13119));
    InMux I__3109 (
            .O(N__13122),
            .I(N__13116));
    LocalMux I__3108 (
            .O(N__13119),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_11 ));
    LocalMux I__3107 (
            .O(N__13116),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_11 ));
    InMux I__3106 (
            .O(N__13111),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_10 ));
    InMux I__3105 (
            .O(N__13108),
            .I(N__13104));
    InMux I__3104 (
            .O(N__13107),
            .I(N__13101));
    LocalMux I__3103 (
            .O(N__13104),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_12 ));
    LocalMux I__3102 (
            .O(N__13101),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_12 ));
    InMux I__3101 (
            .O(N__13096),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_11 ));
    InMux I__3100 (
            .O(N__13093),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_12 ));
    InMux I__3099 (
            .O(N__13090),
            .I(N__13086));
    InMux I__3098 (
            .O(N__13089),
            .I(N__13083));
    LocalMux I__3097 (
            .O(N__13086),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_13 ));
    LocalMux I__3096 (
            .O(N__13083),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_13 ));
    CascadeMux I__3095 (
            .O(N__13078),
            .I(N__13068));
    CascadeMux I__3094 (
            .O(N__13077),
            .I(N__13065));
    CascadeMux I__3093 (
            .O(N__13076),
            .I(N__13062));
    CascadeMux I__3092 (
            .O(N__13075),
            .I(N__13059));
    CascadeMux I__3091 (
            .O(N__13074),
            .I(N__13056));
    CascadeMux I__3090 (
            .O(N__13073),
            .I(N__13052));
    CascadeMux I__3089 (
            .O(N__13072),
            .I(N__13049));
    CascadeMux I__3088 (
            .O(N__13071),
            .I(N__13046));
    InMux I__3087 (
            .O(N__13068),
            .I(N__13034));
    InMux I__3086 (
            .O(N__13065),
            .I(N__13034));
    InMux I__3085 (
            .O(N__13062),
            .I(N__13034));
    InMux I__3084 (
            .O(N__13059),
            .I(N__13023));
    InMux I__3083 (
            .O(N__13056),
            .I(N__13023));
    InMux I__3082 (
            .O(N__13055),
            .I(N__13023));
    InMux I__3081 (
            .O(N__13052),
            .I(N__13023));
    InMux I__3080 (
            .O(N__13049),
            .I(N__13023));
    InMux I__3079 (
            .O(N__13046),
            .I(N__13020));
    CascadeMux I__3078 (
            .O(N__13045),
            .I(N__13017));
    CascadeMux I__3077 (
            .O(N__13044),
            .I(N__13013));
    CascadeMux I__3076 (
            .O(N__13043),
            .I(N__13009));
    CascadeMux I__3075 (
            .O(N__13042),
            .I(N__13005));
    IoInMux I__3074 (
            .O(N__13041),
            .I(N__12999));
    LocalMux I__3073 (
            .O(N__13034),
            .I(N__12993));
    LocalMux I__3072 (
            .O(N__13023),
            .I(N__12988));
    LocalMux I__3071 (
            .O(N__13020),
            .I(N__12988));
    InMux I__3070 (
            .O(N__13017),
            .I(N__12973));
    InMux I__3069 (
            .O(N__13016),
            .I(N__12973));
    InMux I__3068 (
            .O(N__13013),
            .I(N__12973));
    InMux I__3067 (
            .O(N__13012),
            .I(N__12973));
    InMux I__3066 (
            .O(N__13009),
            .I(N__12973));
    InMux I__3065 (
            .O(N__13008),
            .I(N__12973));
    InMux I__3064 (
            .O(N__13005),
            .I(N__12973));
    CascadeMux I__3063 (
            .O(N__13004),
            .I(N__12969));
    CascadeMux I__3062 (
            .O(N__13003),
            .I(N__12966));
    CascadeMux I__3061 (
            .O(N__13002),
            .I(N__12962));
    LocalMux I__3060 (
            .O(N__12999),
            .I(N__12957));
    CascadeMux I__3059 (
            .O(N__12998),
            .I(N__12954));
    CascadeMux I__3058 (
            .O(N__12997),
            .I(N__12950));
    CascadeMux I__3057 (
            .O(N__12996),
            .I(N__12946));
    Span4Mux_v I__3056 (
            .O(N__12993),
            .I(N__12939));
    Span4Mux_v I__3055 (
            .O(N__12988),
            .I(N__12939));
    LocalMux I__3054 (
            .O(N__12973),
            .I(N__12936));
    InMux I__3053 (
            .O(N__12972),
            .I(N__12923));
    InMux I__3052 (
            .O(N__12969),
            .I(N__12923));
    InMux I__3051 (
            .O(N__12966),
            .I(N__12923));
    InMux I__3050 (
            .O(N__12965),
            .I(N__12923));
    InMux I__3049 (
            .O(N__12962),
            .I(N__12923));
    InMux I__3048 (
            .O(N__12961),
            .I(N__12923));
    IoInMux I__3047 (
            .O(N__12960),
            .I(N__12920));
    Span4Mux_s0_v I__3046 (
            .O(N__12957),
            .I(N__12917));
    InMux I__3045 (
            .O(N__12954),
            .I(N__12912));
    InMux I__3044 (
            .O(N__12953),
            .I(N__12912));
    InMux I__3043 (
            .O(N__12950),
            .I(N__12901));
    InMux I__3042 (
            .O(N__12949),
            .I(N__12901));
    InMux I__3041 (
            .O(N__12946),
            .I(N__12901));
    InMux I__3040 (
            .O(N__12945),
            .I(N__12901));
    InMux I__3039 (
            .O(N__12944),
            .I(N__12901));
    Span4Mux_v I__3038 (
            .O(N__12939),
            .I(N__12898));
    Span4Mux_h I__3037 (
            .O(N__12936),
            .I(N__12893));
    LocalMux I__3036 (
            .O(N__12923),
            .I(N__12893));
    LocalMux I__3035 (
            .O(N__12920),
            .I(N__12890));
    Sp12to4 I__3034 (
            .O(N__12917),
            .I(N__12883));
    LocalMux I__3033 (
            .O(N__12912),
            .I(N__12883));
    LocalMux I__3032 (
            .O(N__12901),
            .I(N__12883));
    Span4Mux_v I__3031 (
            .O(N__12898),
            .I(N__12880));
    Span4Mux_v I__3030 (
            .O(N__12893),
            .I(N__12877));
    IoSpan4Mux I__3029 (
            .O(N__12890),
            .I(N__12874));
    Span12Mux_s11_h I__3028 (
            .O(N__12883),
            .I(N__12871));
    Sp12to4 I__3027 (
            .O(N__12880),
            .I(N__12866));
    Sp12to4 I__3026 (
            .O(N__12877),
            .I(N__12866));
    Span4Mux_s3_v I__3025 (
            .O(N__12874),
            .I(N__12863));
    Span12Mux_v I__3024 (
            .O(N__12871),
            .I(N__12858));
    Span12Mux_s11_h I__3023 (
            .O(N__12866),
            .I(N__12858));
    Span4Mux_v I__3022 (
            .O(N__12863),
            .I(N__12855));
    Odrv12 I__3021 (
            .O(N__12858),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3020 (
            .O(N__12855),
            .I(CONSTANT_ONE_NET));
    InMux I__3019 (
            .O(N__12850),
            .I(N__12845));
    InMux I__3018 (
            .O(N__12849),
            .I(N__12842));
    InMux I__3017 (
            .O(N__12848),
            .I(N__12839));
    LocalMux I__3016 (
            .O(N__12845),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_0 ));
    LocalMux I__3015 (
            .O(N__12842),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_0 ));
    LocalMux I__3014 (
            .O(N__12839),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_0 ));
    ClkMux I__3013 (
            .O(N__12832),
            .I(N__12640));
    ClkMux I__3012 (
            .O(N__12831),
            .I(N__12640));
    ClkMux I__3011 (
            .O(N__12830),
            .I(N__12640));
    ClkMux I__3010 (
            .O(N__12829),
            .I(N__12640));
    ClkMux I__3009 (
            .O(N__12828),
            .I(N__12640));
    ClkMux I__3008 (
            .O(N__12827),
            .I(N__12640));
    ClkMux I__3007 (
            .O(N__12826),
            .I(N__12640));
    ClkMux I__3006 (
            .O(N__12825),
            .I(N__12640));
    ClkMux I__3005 (
            .O(N__12824),
            .I(N__12640));
    ClkMux I__3004 (
            .O(N__12823),
            .I(N__12640));
    ClkMux I__3003 (
            .O(N__12822),
            .I(N__12640));
    ClkMux I__3002 (
            .O(N__12821),
            .I(N__12640));
    ClkMux I__3001 (
            .O(N__12820),
            .I(N__12640));
    ClkMux I__3000 (
            .O(N__12819),
            .I(N__12640));
    ClkMux I__2999 (
            .O(N__12818),
            .I(N__12640));
    ClkMux I__2998 (
            .O(N__12817),
            .I(N__12640));
    ClkMux I__2997 (
            .O(N__12816),
            .I(N__12640));
    ClkMux I__2996 (
            .O(N__12815),
            .I(N__12640));
    ClkMux I__2995 (
            .O(N__12814),
            .I(N__12640));
    ClkMux I__2994 (
            .O(N__12813),
            .I(N__12640));
    ClkMux I__2993 (
            .O(N__12812),
            .I(N__12640));
    ClkMux I__2992 (
            .O(N__12811),
            .I(N__12640));
    ClkMux I__2991 (
            .O(N__12810),
            .I(N__12640));
    ClkMux I__2990 (
            .O(N__12809),
            .I(N__12640));
    ClkMux I__2989 (
            .O(N__12808),
            .I(N__12640));
    ClkMux I__2988 (
            .O(N__12807),
            .I(N__12640));
    ClkMux I__2987 (
            .O(N__12806),
            .I(N__12640));
    ClkMux I__2986 (
            .O(N__12805),
            .I(N__12640));
    ClkMux I__2985 (
            .O(N__12804),
            .I(N__12640));
    ClkMux I__2984 (
            .O(N__12803),
            .I(N__12640));
    ClkMux I__2983 (
            .O(N__12802),
            .I(N__12640));
    ClkMux I__2982 (
            .O(N__12801),
            .I(N__12640));
    ClkMux I__2981 (
            .O(N__12800),
            .I(N__12640));
    ClkMux I__2980 (
            .O(N__12799),
            .I(N__12640));
    ClkMux I__2979 (
            .O(N__12798),
            .I(N__12640));
    ClkMux I__2978 (
            .O(N__12797),
            .I(N__12640));
    ClkMux I__2977 (
            .O(N__12796),
            .I(N__12640));
    ClkMux I__2976 (
            .O(N__12795),
            .I(N__12640));
    ClkMux I__2975 (
            .O(N__12794),
            .I(N__12640));
    ClkMux I__2974 (
            .O(N__12793),
            .I(N__12640));
    ClkMux I__2973 (
            .O(N__12792),
            .I(N__12640));
    ClkMux I__2972 (
            .O(N__12791),
            .I(N__12640));
    ClkMux I__2971 (
            .O(N__12790),
            .I(N__12640));
    ClkMux I__2970 (
            .O(N__12789),
            .I(N__12640));
    ClkMux I__2969 (
            .O(N__12788),
            .I(N__12640));
    ClkMux I__2968 (
            .O(N__12787),
            .I(N__12640));
    ClkMux I__2967 (
            .O(N__12786),
            .I(N__12640));
    ClkMux I__2966 (
            .O(N__12785),
            .I(N__12640));
    ClkMux I__2965 (
            .O(N__12784),
            .I(N__12640));
    ClkMux I__2964 (
            .O(N__12783),
            .I(N__12640));
    ClkMux I__2963 (
            .O(N__12782),
            .I(N__12640));
    ClkMux I__2962 (
            .O(N__12781),
            .I(N__12640));
    ClkMux I__2961 (
            .O(N__12780),
            .I(N__12640));
    ClkMux I__2960 (
            .O(N__12779),
            .I(N__12640));
    ClkMux I__2959 (
            .O(N__12778),
            .I(N__12640));
    ClkMux I__2958 (
            .O(N__12777),
            .I(N__12640));
    ClkMux I__2957 (
            .O(N__12776),
            .I(N__12640));
    ClkMux I__2956 (
            .O(N__12775),
            .I(N__12640));
    ClkMux I__2955 (
            .O(N__12774),
            .I(N__12640));
    ClkMux I__2954 (
            .O(N__12773),
            .I(N__12640));
    ClkMux I__2953 (
            .O(N__12772),
            .I(N__12640));
    ClkMux I__2952 (
            .O(N__12771),
            .I(N__12640));
    ClkMux I__2951 (
            .O(N__12770),
            .I(N__12640));
    ClkMux I__2950 (
            .O(N__12769),
            .I(N__12640));
    GlobalMux I__2949 (
            .O(N__12640),
            .I(clk_48mhz));
    SRMux I__2948 (
            .O(N__12637),
            .I(N__12633));
    SRMux I__2947 (
            .O(N__12636),
            .I(N__12630));
    LocalMux I__2946 (
            .O(N__12633),
            .I(N__12627));
    LocalMux I__2945 (
            .O(N__12630),
            .I(N__12624));
    Span4Mux_v I__2944 (
            .O(N__12627),
            .I(N__12621));
    Span4Mux_h I__2943 (
            .O(N__12624),
            .I(N__12618));
    Odrv4 I__2942 (
            .O(N__12621),
            .I(\DUT.uart_inst0.N_20 ));
    Odrv4 I__2941 (
            .O(N__12618),
            .I(\DUT.uart_inst0.N_20 ));
    InMux I__2940 (
            .O(N__12613),
            .I(N__12609));
    InMux I__2939 (
            .O(N__12612),
            .I(N__12606));
    LocalMux I__2938 (
            .O(N__12609),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_1 ));
    LocalMux I__2937 (
            .O(N__12606),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_1 ));
    InMux I__2936 (
            .O(N__12601),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_0 ));
    CascadeMux I__2935 (
            .O(N__12598),
            .I(N__12595));
    InMux I__2934 (
            .O(N__12595),
            .I(N__12591));
    InMux I__2933 (
            .O(N__12594),
            .I(N__12588));
    LocalMux I__2932 (
            .O(N__12591),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_2 ));
    LocalMux I__2931 (
            .O(N__12588),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_2 ));
    InMux I__2930 (
            .O(N__12583),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_1 ));
    CascadeMux I__2929 (
            .O(N__12580),
            .I(N__12576));
    InMux I__2928 (
            .O(N__12579),
            .I(N__12573));
    InMux I__2927 (
            .O(N__12576),
            .I(N__12570));
    LocalMux I__2926 (
            .O(N__12573),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_3 ));
    LocalMux I__2925 (
            .O(N__12570),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_3 ));
    InMux I__2924 (
            .O(N__12565),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_2 ));
    CascadeMux I__2923 (
            .O(N__12562),
            .I(N__12559));
    InMux I__2922 (
            .O(N__12559),
            .I(N__12555));
    InMux I__2921 (
            .O(N__12558),
            .I(N__12552));
    LocalMux I__2920 (
            .O(N__12555),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_4 ));
    LocalMux I__2919 (
            .O(N__12552),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_4 ));
    InMux I__2918 (
            .O(N__12547),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_3 ));
    InMux I__2917 (
            .O(N__12544),
            .I(N__12540));
    InMux I__2916 (
            .O(N__12543),
            .I(N__12537));
    LocalMux I__2915 (
            .O(N__12540),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_5 ));
    LocalMux I__2914 (
            .O(N__12537),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_5 ));
    InMux I__2913 (
            .O(N__12532),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_4 ));
    CascadeMux I__2912 (
            .O(N__12529),
            .I(N__12526));
    InMux I__2911 (
            .O(N__12526),
            .I(N__12522));
    InMux I__2910 (
            .O(N__12525),
            .I(N__12519));
    LocalMux I__2909 (
            .O(N__12522),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_6 ));
    LocalMux I__2908 (
            .O(N__12519),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_6 ));
    InMux I__2907 (
            .O(N__12514),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_5 ));
    CascadeMux I__2906 (
            .O(N__12511),
            .I(N__12507));
    InMux I__2905 (
            .O(N__12510),
            .I(N__12504));
    InMux I__2904 (
            .O(N__12507),
            .I(N__12501));
    LocalMux I__2903 (
            .O(N__12504),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_7 ));
    LocalMux I__2902 (
            .O(N__12501),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_7 ));
    InMux I__2901 (
            .O(N__12496),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_6 ));
    InMux I__2900 (
            .O(N__12493),
            .I(N__12489));
    InMux I__2899 (
            .O(N__12492),
            .I(N__12486));
    LocalMux I__2898 (
            .O(N__12489),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_8 ));
    LocalMux I__2897 (
            .O(N__12486),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_8 ));
    InMux I__2896 (
            .O(N__12481),
            .I(bfn_21_10_0_));
    InMux I__2895 (
            .O(N__12478),
            .I(N__12475));
    LocalMux I__2894 (
            .O(N__12475),
            .I(N__12472));
    Span4Mux_s3_v I__2893 (
            .O(N__12472),
            .I(N__12469));
    Odrv4 I__2892 (
            .O(N__12469),
            .I(rTxBusReady_rep2_i_ess));
    IoInMux I__2891 (
            .O(N__12466),
            .I(N__12463));
    LocalMux I__2890 (
            .O(N__12463),
            .I(N__12460));
    Span4Mux_s1_v I__2889 (
            .O(N__12460),
            .I(N__12457));
    Odrv4 I__2888 (
            .O(N__12457),
            .I(N_1241_i));
    InMux I__2887 (
            .O(N__12454),
            .I(N__12451));
    LocalMux I__2886 (
            .O(N__12451),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_9 ));
    CascadeMux I__2885 (
            .O(N__12448),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_6_cascade_ ));
    CascadeMux I__2884 (
            .O(N__12445),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0_cascade_ ));
    CascadeMux I__2883 (
            .O(N__12442),
            .I(N__12434));
    CascadeMux I__2882 (
            .O(N__12441),
            .I(N__12429));
    CascadeMux I__2881 (
            .O(N__12440),
            .I(N__12425));
    InMux I__2880 (
            .O(N__12439),
            .I(N__12418));
    InMux I__2879 (
            .O(N__12438),
            .I(N__12415));
    InMux I__2878 (
            .O(N__12437),
            .I(N__12410));
    InMux I__2877 (
            .O(N__12434),
            .I(N__12410));
    InMux I__2876 (
            .O(N__12433),
            .I(N__12407));
    InMux I__2875 (
            .O(N__12432),
            .I(N__12404));
    InMux I__2874 (
            .O(N__12429),
            .I(N__12401));
    InMux I__2873 (
            .O(N__12428),
            .I(N__12398));
    InMux I__2872 (
            .O(N__12425),
            .I(N__12395));
    InMux I__2871 (
            .O(N__12424),
            .I(N__12392));
    InMux I__2870 (
            .O(N__12423),
            .I(N__12389));
    InMux I__2869 (
            .O(N__12422),
            .I(N__12386));
    InMux I__2868 (
            .O(N__12421),
            .I(N__12383));
    LocalMux I__2867 (
            .O(N__12418),
            .I(N__12380));
    LocalMux I__2866 (
            .O(N__12415),
            .I(N__12377));
    LocalMux I__2865 (
            .O(N__12410),
            .I(N__12372));
    LocalMux I__2864 (
            .O(N__12407),
            .I(N__12369));
    LocalMux I__2863 (
            .O(N__12404),
            .I(N__12366));
    LocalMux I__2862 (
            .O(N__12401),
            .I(N__12363));
    LocalMux I__2861 (
            .O(N__12398),
            .I(N__12360));
    LocalMux I__2860 (
            .O(N__12395),
            .I(N__12357));
    LocalMux I__2859 (
            .O(N__12392),
            .I(N__12354));
    LocalMux I__2858 (
            .O(N__12389),
            .I(N__12350));
    LocalMux I__2857 (
            .O(N__12386),
            .I(N__12347));
    LocalMux I__2856 (
            .O(N__12383),
            .I(N__12341));
    Glb2LocalMux I__2855 (
            .O(N__12380),
            .I(N__12301));
    Glb2LocalMux I__2854 (
            .O(N__12377),
            .I(N__12301));
    CEMux I__2853 (
            .O(N__12376),
            .I(N__12301));
    CEMux I__2852 (
            .O(N__12375),
            .I(N__12301));
    Glb2LocalMux I__2851 (
            .O(N__12372),
            .I(N__12301));
    Glb2LocalMux I__2850 (
            .O(N__12369),
            .I(N__12301));
    Glb2LocalMux I__2849 (
            .O(N__12366),
            .I(N__12301));
    Glb2LocalMux I__2848 (
            .O(N__12363),
            .I(N__12301));
    Glb2LocalMux I__2847 (
            .O(N__12360),
            .I(N__12301));
    Glb2LocalMux I__2846 (
            .O(N__12357),
            .I(N__12301));
    Glb2LocalMux I__2845 (
            .O(N__12354),
            .I(N__12301));
    CEMux I__2844 (
            .O(N__12353),
            .I(N__12301));
    Glb2LocalMux I__2843 (
            .O(N__12350),
            .I(N__12301));
    Glb2LocalMux I__2842 (
            .O(N__12347),
            .I(N__12301));
    CEMux I__2841 (
            .O(N__12346),
            .I(N__12301));
    CEMux I__2840 (
            .O(N__12345),
            .I(N__12301));
    CEMux I__2839 (
            .O(N__12344),
            .I(N__12301));
    Glb2LocalMux I__2838 (
            .O(N__12341),
            .I(N__12301));
    CEMux I__2837 (
            .O(N__12340),
            .I(N__12301));
    GlobalMux I__2836 (
            .O(N__12301),
            .I(N__12298));
    gio2CtrlBuf I__2835 (
            .O(N__12298),
            .I(wPllLocked_g));
    InMux I__2834 (
            .O(N__12295),
            .I(N__12292));
    LocalMux I__2833 (
            .O(N__12292),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_8 ));
    InMux I__2832 (
            .O(N__12289),
            .I(N__12286));
    LocalMux I__2831 (
            .O(N__12286),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_7 ));
    InMux I__2830 (
            .O(N__12283),
            .I(N__12278));
    InMux I__2829 (
            .O(N__12282),
            .I(N__12275));
    InMux I__2828 (
            .O(N__12281),
            .I(N__12272));
    LocalMux I__2827 (
            .O(N__12278),
            .I(N__12269));
    LocalMux I__2826 (
            .O(N__12275),
            .I(N__12266));
    LocalMux I__2825 (
            .O(N__12272),
            .I(N__12263));
    Span4Mux_v I__2824 (
            .O(N__12269),
            .I(N__12260));
    Span4Mux_h I__2823 (
            .O(N__12266),
            .I(N__12257));
    Odrv4 I__2822 (
            .O(N__12263),
            .I(\DUT.uart_inst0.N_77 ));
    Odrv4 I__2821 (
            .O(N__12260),
            .I(\DUT.uart_inst0.N_77 ));
    Odrv4 I__2820 (
            .O(N__12257),
            .I(\DUT.uart_inst0.N_77 ));
    CascadeMux I__2819 (
            .O(N__12250),
            .I(N__12240));
    InMux I__2818 (
            .O(N__12249),
            .I(N__12237));
    CascadeMux I__2817 (
            .O(N__12248),
            .I(N__12234));
    CascadeMux I__2816 (
            .O(N__12247),
            .I(N__12231));
    InMux I__2815 (
            .O(N__12246),
            .I(N__12225));
    InMux I__2814 (
            .O(N__12245),
            .I(N__12225));
    InMux I__2813 (
            .O(N__12244),
            .I(N__12218));
    InMux I__2812 (
            .O(N__12243),
            .I(N__12218));
    InMux I__2811 (
            .O(N__12240),
            .I(N__12215));
    LocalMux I__2810 (
            .O(N__12237),
            .I(N__12212));
    InMux I__2809 (
            .O(N__12234),
            .I(N__12205));
    InMux I__2808 (
            .O(N__12231),
            .I(N__12205));
    InMux I__2807 (
            .O(N__12230),
            .I(N__12205));
    LocalMux I__2806 (
            .O(N__12225),
            .I(N__12202));
    InMux I__2805 (
            .O(N__12224),
            .I(N__12197));
    InMux I__2804 (
            .O(N__12223),
            .I(N__12197));
    LocalMux I__2803 (
            .O(N__12218),
            .I(N__12193));
    LocalMux I__2802 (
            .O(N__12215),
            .I(N__12190));
    Span4Mux_h I__2801 (
            .O(N__12212),
            .I(N__12187));
    LocalMux I__2800 (
            .O(N__12205),
            .I(N__12180));
    Span4Mux_v I__2799 (
            .O(N__12202),
            .I(N__12180));
    LocalMux I__2798 (
            .O(N__12197),
            .I(N__12180));
    InMux I__2797 (
            .O(N__12196),
            .I(N__12177));
    Span4Mux_h I__2796 (
            .O(N__12193),
            .I(N__12174));
    Odrv12 I__2795 (
            .O(N__12190),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0 ));
    Odrv4 I__2794 (
            .O(N__12187),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0 ));
    Odrv4 I__2793 (
            .O(N__12180),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0 ));
    LocalMux I__2792 (
            .O(N__12177),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0 ));
    Odrv4 I__2791 (
            .O(N__12174),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0 ));
    CascadeMux I__2790 (
            .O(N__12163),
            .I(N__12159));
    InMux I__2789 (
            .O(N__12162),
            .I(N__12154));
    InMux I__2788 (
            .O(N__12159),
            .I(N__12147));
    InMux I__2787 (
            .O(N__12158),
            .I(N__12147));
    InMux I__2786 (
            .O(N__12157),
            .I(N__12147));
    LocalMux I__2785 (
            .O(N__12154),
            .I(N__12142));
    LocalMux I__2784 (
            .O(N__12147),
            .I(N__12142));
    Odrv4 I__2783 (
            .O(N__12142),
            .I(\DUT.uart_inst0.N_147 ));
    CascadeMux I__2782 (
            .O(N__12139),
            .I(N__12136));
    InMux I__2781 (
            .O(N__12136),
            .I(N__12127));
    InMux I__2780 (
            .O(N__12135),
            .I(N__12127));
    InMux I__2779 (
            .O(N__12134),
            .I(N__12124));
    InMux I__2778 (
            .O(N__12133),
            .I(N__12119));
    InMux I__2777 (
            .O(N__12132),
            .I(N__12119));
    LocalMux I__2776 (
            .O(N__12127),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_2 ));
    LocalMux I__2775 (
            .O(N__12124),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_2 ));
    LocalMux I__2774 (
            .O(N__12119),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_2 ));
    CascadeMux I__2773 (
            .O(N__12112),
            .I(\DUT.uart_inst0.tx_countdown_0_c4_cascade_ ));
    InMux I__2772 (
            .O(N__12109),
            .I(N__12106));
    LocalMux I__2771 (
            .O(N__12106),
            .I(\DUT.uart_inst0.tx_countdown_7_ns_1_4 ));
    CascadeMux I__2770 (
            .O(N__12103),
            .I(\DUT.uart_inst0.tx_countdown_7_ns_1_1_cascade_ ));
    CascadeMux I__2769 (
            .O(N__12100),
            .I(N__12097));
    InMux I__2768 (
            .O(N__12097),
            .I(N__12094));
    LocalMux I__2767 (
            .O(N__12094),
            .I(\DUT.uart_inst0.tx_countdown_0_c4 ));
    InMux I__2766 (
            .O(N__12091),
            .I(N__12088));
    LocalMux I__2765 (
            .O(N__12088),
            .I(\DUT.uart_inst0.tx_countdown_7_ns_1_5 ));
    InMux I__2764 (
            .O(N__12085),
            .I(N__12075));
    InMux I__2763 (
            .O(N__12084),
            .I(N__12070));
    InMux I__2762 (
            .O(N__12083),
            .I(N__12070));
    InMux I__2761 (
            .O(N__12082),
            .I(N__12063));
    InMux I__2760 (
            .O(N__12081),
            .I(N__12063));
    InMux I__2759 (
            .O(N__12080),
            .I(N__12063));
    InMux I__2758 (
            .O(N__12079),
            .I(N__12058));
    InMux I__2757 (
            .O(N__12078),
            .I(N__12058));
    LocalMux I__2756 (
            .O(N__12075),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_0 ));
    LocalMux I__2755 (
            .O(N__12070),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_0 ));
    LocalMux I__2754 (
            .O(N__12063),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_0 ));
    LocalMux I__2753 (
            .O(N__12058),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_0 ));
    CascadeMux I__2752 (
            .O(N__12049),
            .I(N__12039));
    InMux I__2751 (
            .O(N__12048),
            .I(N__12034));
    InMux I__2750 (
            .O(N__12047),
            .I(N__12034));
    InMux I__2749 (
            .O(N__12046),
            .I(N__12029));
    InMux I__2748 (
            .O(N__12045),
            .I(N__12029));
    InMux I__2747 (
            .O(N__12044),
            .I(N__12024));
    InMux I__2746 (
            .O(N__12043),
            .I(N__12024));
    InMux I__2745 (
            .O(N__12042),
            .I(N__12019));
    InMux I__2744 (
            .O(N__12039),
            .I(N__12019));
    LocalMux I__2743 (
            .O(N__12034),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_1 ));
    LocalMux I__2742 (
            .O(N__12029),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_1 ));
    LocalMux I__2741 (
            .O(N__12024),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_1 ));
    LocalMux I__2740 (
            .O(N__12019),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_1 ));
    CascadeMux I__2739 (
            .O(N__12010),
            .I(N__12003));
    InMux I__2738 (
            .O(N__12009),
            .I(N__12000));
    InMux I__2737 (
            .O(N__12008),
            .I(N__11995));
    InMux I__2736 (
            .O(N__12007),
            .I(N__11995));
    InMux I__2735 (
            .O(N__12006),
            .I(N__11990));
    InMux I__2734 (
            .O(N__12003),
            .I(N__11990));
    LocalMux I__2733 (
            .O(N__12000),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_5 ));
    LocalMux I__2732 (
            .O(N__11995),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_5 ));
    LocalMux I__2731 (
            .O(N__11990),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_5 ));
    CascadeMux I__2730 (
            .O(N__11983),
            .I(\DUT.uart_inst0.tx_countdown_7_m1_0_o2_1_2_cascade_ ));
    InMux I__2729 (
            .O(N__11980),
            .I(N__11972));
    InMux I__2728 (
            .O(N__11979),
            .I(N__11965));
    InMux I__2727 (
            .O(N__11978),
            .I(N__11965));
    InMux I__2726 (
            .O(N__11977),
            .I(N__11965));
    InMux I__2725 (
            .O(N__11976),
            .I(N__11960));
    InMux I__2724 (
            .O(N__11975),
            .I(N__11960));
    LocalMux I__2723 (
            .O(N__11972),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_4 ));
    LocalMux I__2722 (
            .O(N__11965),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_4 ));
    LocalMux I__2721 (
            .O(N__11960),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_4 ));
    InMux I__2720 (
            .O(N__11953),
            .I(N__11950));
    LocalMux I__2719 (
            .O(N__11950),
            .I(N__11947));
    Odrv4 I__2718 (
            .O(N__11947),
            .I(\DUT.uart_inst0.N_68 ));
    InMux I__2717 (
            .O(N__11944),
            .I(N__11935));
    InMux I__2716 (
            .O(N__11943),
            .I(N__11935));
    InMux I__2715 (
            .O(N__11942),
            .I(N__11935));
    LocalMux I__2714 (
            .O(N__11935),
            .I(N__11932));
    Span4Mux_h I__2713 (
            .O(N__11932),
            .I(N__11929));
    Odrv4 I__2712 (
            .O(N__11929),
            .I(\DUT.uart_inst0.N_146 ));
    CascadeMux I__2711 (
            .O(N__11926),
            .I(N__11922));
    InMux I__2710 (
            .O(N__11925),
            .I(N__11914));
    InMux I__2709 (
            .O(N__11922),
            .I(N__11911));
    InMux I__2708 (
            .O(N__11921),
            .I(N__11902));
    InMux I__2707 (
            .O(N__11920),
            .I(N__11902));
    InMux I__2706 (
            .O(N__11919),
            .I(N__11902));
    InMux I__2705 (
            .O(N__11918),
            .I(N__11902));
    InMux I__2704 (
            .O(N__11917),
            .I(N__11899));
    LocalMux I__2703 (
            .O(N__11914),
            .I(\DUT.uart_inst0.tx_countdown_7_sm0_0 ));
    LocalMux I__2702 (
            .O(N__11911),
            .I(\DUT.uart_inst0.tx_countdown_7_sm0_0 ));
    LocalMux I__2701 (
            .O(N__11902),
            .I(\DUT.uart_inst0.tx_countdown_7_sm0_0 ));
    LocalMux I__2700 (
            .O(N__11899),
            .I(\DUT.uart_inst0.tx_countdown_7_sm0_0 ));
    InMux I__2699 (
            .O(N__11890),
            .I(N__11887));
    LocalMux I__2698 (
            .O(N__11887),
            .I(\DUT.uart_inst0.tx_countdown_7_ns_1_3 ));
    CascadeMux I__2697 (
            .O(N__11884),
            .I(N__11879));
    CascadeMux I__2696 (
            .O(N__11883),
            .I(N__11876));
    InMux I__2695 (
            .O(N__11882),
            .I(N__11870));
    InMux I__2694 (
            .O(N__11879),
            .I(N__11867));
    InMux I__2693 (
            .O(N__11876),
            .I(N__11862));
    InMux I__2692 (
            .O(N__11875),
            .I(N__11862));
    InMux I__2691 (
            .O(N__11874),
            .I(N__11857));
    InMux I__2690 (
            .O(N__11873),
            .I(N__11857));
    LocalMux I__2689 (
            .O(N__11870),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_3 ));
    LocalMux I__2688 (
            .O(N__11867),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_3 ));
    LocalMux I__2687 (
            .O(N__11862),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_3 ));
    LocalMux I__2686 (
            .O(N__11857),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_3 ));
    CascadeMux I__2685 (
            .O(N__11848),
            .I(\DUT.uart_inst0.tx_state_RNI8CH01Z0Z_1_cascade_ ));
    SRMux I__2684 (
            .O(N__11845),
            .I(N__11842));
    LocalMux I__2683 (
            .O(N__11842),
            .I(\DUT.uart_inst0.N_59_i ));
    InMux I__2682 (
            .O(N__11839),
            .I(N__11836));
    LocalMux I__2681 (
            .O(N__11836),
            .I(N__11833));
    Span4Mux_h I__2680 (
            .O(N__11833),
            .I(N__11829));
    InMux I__2679 (
            .O(N__11832),
            .I(N__11826));
    Odrv4 I__2678 (
            .O(N__11829),
            .I(\DUT.N_93 ));
    LocalMux I__2677 (
            .O(N__11826),
            .I(\DUT.N_93 ));
    InMux I__2676 (
            .O(N__11821),
            .I(N__11815));
    CascadeMux I__2675 (
            .O(N__11820),
            .I(N__11812));
    CascadeMux I__2674 (
            .O(N__11819),
            .I(N__11809));
    CascadeMux I__2673 (
            .O(N__11818),
            .I(N__11805));
    LocalMux I__2672 (
            .O(N__11815),
            .I(N__11798));
    InMux I__2671 (
            .O(N__11812),
            .I(N__11795));
    InMux I__2670 (
            .O(N__11809),
            .I(N__11792));
    InMux I__2669 (
            .O(N__11808),
            .I(N__11789));
    InMux I__2668 (
            .O(N__11805),
            .I(N__11784));
    InMux I__2667 (
            .O(N__11804),
            .I(N__11784));
    InMux I__2666 (
            .O(N__11803),
            .I(N__11779));
    InMux I__2665 (
            .O(N__11802),
            .I(N__11779));
    InMux I__2664 (
            .O(N__11801),
            .I(N__11776));
    Span4Mux_v I__2663 (
            .O(N__11798),
            .I(N__11773));
    LocalMux I__2662 (
            .O(N__11795),
            .I(N__11764));
    LocalMux I__2661 (
            .O(N__11792),
            .I(N__11764));
    LocalMux I__2660 (
            .O(N__11789),
            .I(N__11764));
    LocalMux I__2659 (
            .O(N__11784),
            .I(N__11764));
    LocalMux I__2658 (
            .O(N__11779),
            .I(\DUT.tx_state_1 ));
    LocalMux I__2657 (
            .O(N__11776),
            .I(\DUT.tx_state_1 ));
    Odrv4 I__2656 (
            .O(N__11773),
            .I(\DUT.tx_state_1 ));
    Odrv4 I__2655 (
            .O(N__11764),
            .I(\DUT.tx_state_1 ));
    CascadeMux I__2654 (
            .O(N__11755),
            .I(N__11750));
    InMux I__2653 (
            .O(N__11754),
            .I(N__11743));
    InMux I__2652 (
            .O(N__11753),
            .I(N__11740));
    InMux I__2651 (
            .O(N__11750),
            .I(N__11737));
    InMux I__2650 (
            .O(N__11749),
            .I(N__11730));
    InMux I__2649 (
            .O(N__11748),
            .I(N__11730));
    InMux I__2648 (
            .O(N__11747),
            .I(N__11730));
    InMux I__2647 (
            .O(N__11746),
            .I(N__11727));
    LocalMux I__2646 (
            .O(N__11743),
            .I(N__11724));
    LocalMux I__2645 (
            .O(N__11740),
            .I(N__11719));
    LocalMux I__2644 (
            .O(N__11737),
            .I(N__11719));
    LocalMux I__2643 (
            .O(N__11730),
            .I(N__11716));
    LocalMux I__2642 (
            .O(N__11727),
            .I(N__11713));
    Span4Mux_v I__2641 (
            .O(N__11724),
            .I(N__11708));
    Span4Mux_v I__2640 (
            .O(N__11719),
            .I(N__11705));
    Span4Mux_h I__2639 (
            .O(N__11716),
            .I(N__11702));
    Span4Mux_h I__2638 (
            .O(N__11713),
            .I(N__11699));
    InMux I__2637 (
            .O(N__11712),
            .I(N__11696));
    InMux I__2636 (
            .O(N__11711),
            .I(N__11693));
    Odrv4 I__2635 (
            .O(N__11708),
            .I(\DUT.rTransmitZ0 ));
    Odrv4 I__2634 (
            .O(N__11705),
            .I(\DUT.rTransmitZ0 ));
    Odrv4 I__2633 (
            .O(N__11702),
            .I(\DUT.rTransmitZ0 ));
    Odrv4 I__2632 (
            .O(N__11699),
            .I(\DUT.rTransmitZ0 ));
    LocalMux I__2631 (
            .O(N__11696),
            .I(\DUT.rTransmitZ0 ));
    LocalMux I__2630 (
            .O(N__11693),
            .I(\DUT.rTransmitZ0 ));
    CascadeMux I__2629 (
            .O(N__11680),
            .I(N__11671));
    CascadeMux I__2628 (
            .O(N__11679),
            .I(N__11667));
    CascadeMux I__2627 (
            .O(N__11678),
            .I(N__11662));
    CascadeMux I__2626 (
            .O(N__11677),
            .I(N__11653));
    CascadeMux I__2625 (
            .O(N__11676),
            .I(N__11648));
    InMux I__2624 (
            .O(N__11675),
            .I(N__11641));
    InMux I__2623 (
            .O(N__11674),
            .I(N__11641));
    InMux I__2622 (
            .O(N__11671),
            .I(N__11641));
    InMux I__2621 (
            .O(N__11670),
            .I(N__11636));
    InMux I__2620 (
            .O(N__11667),
            .I(N__11636));
    InMux I__2619 (
            .O(N__11666),
            .I(N__11625));
    InMux I__2618 (
            .O(N__11665),
            .I(N__11625));
    InMux I__2617 (
            .O(N__11662),
            .I(N__11625));
    InMux I__2616 (
            .O(N__11661),
            .I(N__11625));
    InMux I__2615 (
            .O(N__11660),
            .I(N__11625));
    InMux I__2614 (
            .O(N__11659),
            .I(N__11614));
    InMux I__2613 (
            .O(N__11658),
            .I(N__11614));
    InMux I__2612 (
            .O(N__11657),
            .I(N__11614));
    InMux I__2611 (
            .O(N__11656),
            .I(N__11614));
    InMux I__2610 (
            .O(N__11653),
            .I(N__11614));
    InMux I__2609 (
            .O(N__11652),
            .I(N__11607));
    InMux I__2608 (
            .O(N__11651),
            .I(N__11607));
    InMux I__2607 (
            .O(N__11648),
            .I(N__11607));
    LocalMux I__2606 (
            .O(N__11641),
            .I(N__11604));
    LocalMux I__2605 (
            .O(N__11636),
            .I(N__11595));
    LocalMux I__2604 (
            .O(N__11625),
            .I(N__11595));
    LocalMux I__2603 (
            .O(N__11614),
            .I(N__11595));
    LocalMux I__2602 (
            .O(N__11607),
            .I(N__11592));
    Span4Mux_v I__2601 (
            .O(N__11604),
            .I(N__11589));
    InMux I__2600 (
            .O(N__11603),
            .I(N__11584));
    InMux I__2599 (
            .O(N__11602),
            .I(N__11584));
    Span4Mux_v I__2598 (
            .O(N__11595),
            .I(N__11581));
    Span4Mux_h I__2597 (
            .O(N__11592),
            .I(N__11576));
    Span4Mux_h I__2596 (
            .O(N__11589),
            .I(N__11576));
    LocalMux I__2595 (
            .O(N__11584),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    Odrv4 I__2594 (
            .O(N__11581),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    Odrv4 I__2593 (
            .O(N__11576),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    InMux I__2592 (
            .O(N__11569),
            .I(N__11566));
    LocalMux I__2591 (
            .O(N__11566),
            .I(\DUT.fifo_tx_inst.un1_i11_2_i ));
    InMux I__2590 (
            .O(N__11563),
            .I(N__11554));
    InMux I__2589 (
            .O(N__11562),
            .I(N__11554));
    InMux I__2588 (
            .O(N__11561),
            .I(N__11554));
    LocalMux I__2587 (
            .O(N__11554),
            .I(N__11551));
    Span4Mux_h I__2586 (
            .O(N__11551),
            .I(N__11548));
    Odrv4 I__2585 (
            .O(N__11548),
            .I(\DUT.fifo_tx_inst.rReadPtr11 ));
    CascadeMux I__2584 (
            .O(N__11545),
            .I(\DUT.fifo_tx_inst.un1_i11_2_i_cascade_ ));
    InMux I__2583 (
            .O(N__11542),
            .I(N__11531));
    InMux I__2582 (
            .O(N__11541),
            .I(N__11524));
    InMux I__2581 (
            .O(N__11540),
            .I(N__11524));
    InMux I__2580 (
            .O(N__11539),
            .I(N__11524));
    InMux I__2579 (
            .O(N__11538),
            .I(N__11517));
    InMux I__2578 (
            .O(N__11537),
            .I(N__11517));
    InMux I__2577 (
            .O(N__11536),
            .I(N__11512));
    InMux I__2576 (
            .O(N__11535),
            .I(N__11512));
    CascadeMux I__2575 (
            .O(N__11534),
            .I(N__11508));
    LocalMux I__2574 (
            .O(N__11531),
            .I(N__11504));
    LocalMux I__2573 (
            .O(N__11524),
            .I(N__11501));
    InMux I__2572 (
            .O(N__11523),
            .I(N__11496));
    InMux I__2571 (
            .O(N__11522),
            .I(N__11496));
    LocalMux I__2570 (
            .O(N__11517),
            .I(N__11491));
    LocalMux I__2569 (
            .O(N__11512),
            .I(N__11491));
    InMux I__2568 (
            .O(N__11511),
            .I(N__11488));
    InMux I__2567 (
            .O(N__11508),
            .I(N__11483));
    InMux I__2566 (
            .O(N__11507),
            .I(N__11483));
    Span4Mux_h I__2565 (
            .O(N__11504),
            .I(N__11480));
    Span4Mux_v I__2564 (
            .O(N__11501),
            .I(N__11475));
    LocalMux I__2563 (
            .O(N__11496),
            .I(N__11475));
    Span4Mux_h I__2562 (
            .O(N__11491),
            .I(N__11472));
    LocalMux I__2561 (
            .O(N__11488),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__2560 (
            .O(N__11483),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    Odrv4 I__2559 (
            .O(N__11480),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    Odrv4 I__2558 (
            .O(N__11475),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    Odrv4 I__2557 (
            .O(N__11472),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    InMux I__2556 (
            .O(N__11461),
            .I(N__11456));
    InMux I__2555 (
            .O(N__11460),
            .I(N__11453));
    InMux I__2554 (
            .O(N__11459),
            .I(N__11450));
    LocalMux I__2553 (
            .O(N__11456),
            .I(\DUT.uart_inst0.N_74 ));
    LocalMux I__2552 (
            .O(N__11453),
            .I(\DUT.uart_inst0.N_74 ));
    LocalMux I__2551 (
            .O(N__11450),
            .I(\DUT.uart_inst0.N_74 ));
    CascadeMux I__2550 (
            .O(N__11443),
            .I(N__11438));
    CascadeMux I__2549 (
            .O(N__11442),
            .I(N__11429));
    InMux I__2548 (
            .O(N__11441),
            .I(N__11424));
    InMux I__2547 (
            .O(N__11438),
            .I(N__11419));
    InMux I__2546 (
            .O(N__11437),
            .I(N__11412));
    InMux I__2545 (
            .O(N__11436),
            .I(N__11412));
    InMux I__2544 (
            .O(N__11435),
            .I(N__11412));
    InMux I__2543 (
            .O(N__11434),
            .I(N__11409));
    InMux I__2542 (
            .O(N__11433),
            .I(N__11399));
    InMux I__2541 (
            .O(N__11432),
            .I(N__11399));
    InMux I__2540 (
            .O(N__11429),
            .I(N__11399));
    InMux I__2539 (
            .O(N__11428),
            .I(N__11396));
    CascadeMux I__2538 (
            .O(N__11427),
            .I(N__11388));
    LocalMux I__2537 (
            .O(N__11424),
            .I(N__11385));
    InMux I__2536 (
            .O(N__11423),
            .I(N__11380));
    InMux I__2535 (
            .O(N__11422),
            .I(N__11380));
    LocalMux I__2534 (
            .O(N__11419),
            .I(N__11375));
    LocalMux I__2533 (
            .O(N__11412),
            .I(N__11375));
    LocalMux I__2532 (
            .O(N__11409),
            .I(N__11372));
    InMux I__2531 (
            .O(N__11408),
            .I(N__11363));
    InMux I__2530 (
            .O(N__11407),
            .I(N__11363));
    InMux I__2529 (
            .O(N__11406),
            .I(N__11363));
    LocalMux I__2528 (
            .O(N__11399),
            .I(N__11360));
    LocalMux I__2527 (
            .O(N__11396),
            .I(N__11357));
    InMux I__2526 (
            .O(N__11395),
            .I(N__11350));
    InMux I__2525 (
            .O(N__11394),
            .I(N__11350));
    InMux I__2524 (
            .O(N__11393),
            .I(N__11350));
    InMux I__2523 (
            .O(N__11392),
            .I(N__11345));
    InMux I__2522 (
            .O(N__11391),
            .I(N__11345));
    InMux I__2521 (
            .O(N__11388),
            .I(N__11342));
    Span12Mux_s10_v I__2520 (
            .O(N__11385),
            .I(N__11339));
    LocalMux I__2519 (
            .O(N__11380),
            .I(N__11336));
    Span4Mux_v I__2518 (
            .O(N__11375),
            .I(N__11331));
    Span4Mux_h I__2517 (
            .O(N__11372),
            .I(N__11331));
    InMux I__2516 (
            .O(N__11371),
            .I(N__11328));
    InMux I__2515 (
            .O(N__11370),
            .I(N__11325));
    LocalMux I__2514 (
            .O(N__11363),
            .I(N__11318));
    Span4Mux_h I__2513 (
            .O(N__11360),
            .I(N__11318));
    Span4Mux_h I__2512 (
            .O(N__11357),
            .I(N__11318));
    LocalMux I__2511 (
            .O(N__11350),
            .I(N__11313));
    LocalMux I__2510 (
            .O(N__11345),
            .I(N__11313));
    LocalMux I__2509 (
            .O(N__11342),
            .I(\DUT.tx_state_0 ));
    Odrv12 I__2508 (
            .O(N__11339),
            .I(\DUT.tx_state_0 ));
    Odrv4 I__2507 (
            .O(N__11336),
            .I(\DUT.tx_state_0 ));
    Odrv4 I__2506 (
            .O(N__11331),
            .I(\DUT.tx_state_0 ));
    LocalMux I__2505 (
            .O(N__11328),
            .I(\DUT.tx_state_0 ));
    LocalMux I__2504 (
            .O(N__11325),
            .I(\DUT.tx_state_0 ));
    Odrv4 I__2503 (
            .O(N__11318),
            .I(\DUT.tx_state_0 ));
    Odrv12 I__2502 (
            .O(N__11313),
            .I(\DUT.tx_state_0 ));
    InMux I__2501 (
            .O(N__11296),
            .I(N__11293));
    LocalMux I__2500 (
            .O(N__11293),
            .I(\DUT.uart_inst0.tx_countdown_7_1_2 ));
    CascadeMux I__2499 (
            .O(N__11290),
            .I(N__11287));
    InMux I__2498 (
            .O(N__11287),
            .I(N__11284));
    LocalMux I__2497 (
            .O(N__11284),
            .I(\DUT.uart_inst0.N_91 ));
    InMux I__2496 (
            .O(N__11281),
            .I(N__11278));
    LocalMux I__2495 (
            .O(N__11278),
            .I(rTxBusReady_rep1_i_ess));
    InMux I__2494 (
            .O(N__11275),
            .I(N__11272));
    LocalMux I__2493 (
            .O(N__11272),
            .I(N__11269));
    Odrv12 I__2492 (
            .O(N__11269),
            .I(rTxBusReady_rep3_i_ess));
    InMux I__2491 (
            .O(N__11266),
            .I(N__11263));
    LocalMux I__2490 (
            .O(N__11263),
            .I(N__11260));
    Span4Mux_s3_v I__2489 (
            .O(N__11260),
            .I(N__11257));
    Odrv4 I__2488 (
            .O(N__11257),
            .I(rTxBusReady_rep0_i_ess));
    InMux I__2487 (
            .O(N__11254),
            .I(N__11251));
    LocalMux I__2486 (
            .O(N__11251),
            .I(N__11245));
    InMux I__2485 (
            .O(N__11250),
            .I(N__11242));
    CascadeMux I__2484 (
            .O(N__11249),
            .I(N__11236));
    CascadeMux I__2483 (
            .O(N__11248),
            .I(N__11232));
    Span4Mux_h I__2482 (
            .O(N__11245),
            .I(N__11227));
    LocalMux I__2481 (
            .O(N__11242),
            .I(N__11227));
    InMux I__2480 (
            .O(N__11241),
            .I(N__11224));
    InMux I__2479 (
            .O(N__11240),
            .I(N__11215));
    InMux I__2478 (
            .O(N__11239),
            .I(N__11215));
    InMux I__2477 (
            .O(N__11236),
            .I(N__11215));
    InMux I__2476 (
            .O(N__11235),
            .I(N__11215));
    InMux I__2475 (
            .O(N__11232),
            .I(N__11212));
    Span4Mux_v I__2474 (
            .O(N__11227),
            .I(N__11209));
    LocalMux I__2473 (
            .O(N__11224),
            .I(N__11206));
    LocalMux I__2472 (
            .O(N__11215),
            .I(N__11201));
    LocalMux I__2471 (
            .O(N__11212),
            .I(N__11201));
    Sp12to4 I__2470 (
            .O(N__11209),
            .I(N__11198));
    Span4Mux_h I__2469 (
            .O(N__11206),
            .I(N__11195));
    Span12Mux_v I__2468 (
            .O(N__11201),
            .I(N__11188));
    Span12Mux_s7_h I__2467 (
            .O(N__11198),
            .I(N__11188));
    Sp12to4 I__2466 (
            .O(N__11195),
            .I(N__11188));
    Span12Mux_v I__2465 (
            .O(N__11188),
            .I(N__11185));
    Odrv12 I__2464 (
            .O(N__11185),
            .I(iTxE_n_c));
    InMux I__2463 (
            .O(N__11182),
            .I(N__11178));
    InMux I__2462 (
            .O(N__11181),
            .I(N__11175));
    LocalMux I__2461 (
            .O(N__11178),
            .I(N__11172));
    LocalMux I__2460 (
            .O(N__11175),
            .I(N__11167));
    Span4Mux_h I__2459 (
            .O(N__11172),
            .I(N__11164));
    InMux I__2458 (
            .O(N__11171),
            .I(N__11159));
    InMux I__2457 (
            .O(N__11170),
            .I(N__11159));
    Span12Mux_s9_v I__2456 (
            .O(N__11167),
            .I(N__11156));
    Odrv4 I__2455 (
            .O(N__11164),
            .I(\fifo_inst.ftdi_output_inst.N_68_0 ));
    LocalMux I__2454 (
            .O(N__11159),
            .I(\fifo_inst.ftdi_output_inst.N_68_0 ));
    Odrv12 I__2453 (
            .O(N__11156),
            .I(\fifo_inst.ftdi_output_inst.N_68_0 ));
    InMux I__2452 (
            .O(N__11149),
            .I(N__11143));
    InMux I__2451 (
            .O(N__11148),
            .I(N__11138));
    InMux I__2450 (
            .O(N__11147),
            .I(N__11138));
    InMux I__2449 (
            .O(N__11146),
            .I(N__11135));
    LocalMux I__2448 (
            .O(N__11143),
            .I(N__11131));
    LocalMux I__2447 (
            .O(N__11138),
            .I(N__11126));
    LocalMux I__2446 (
            .O(N__11135),
            .I(N__11120));
    SRMux I__2445 (
            .O(N__11134),
            .I(N__11074));
    Glb2LocalMux I__2444 (
            .O(N__11131),
            .I(N__11074));
    SRMux I__2443 (
            .O(N__11130),
            .I(N__11074));
    SRMux I__2442 (
            .O(N__11129),
            .I(N__11074));
    Glb2LocalMux I__2441 (
            .O(N__11126),
            .I(N__11074));
    SRMux I__2440 (
            .O(N__11125),
            .I(N__11074));
    SRMux I__2439 (
            .O(N__11124),
            .I(N__11074));
    SRMux I__2438 (
            .O(N__11123),
            .I(N__11074));
    Glb2LocalMux I__2437 (
            .O(N__11120),
            .I(N__11074));
    SRMux I__2436 (
            .O(N__11119),
            .I(N__11074));
    SRMux I__2435 (
            .O(N__11118),
            .I(N__11074));
    SRMux I__2434 (
            .O(N__11117),
            .I(N__11074));
    SRMux I__2433 (
            .O(N__11116),
            .I(N__11074));
    SRMux I__2432 (
            .O(N__11115),
            .I(N__11074));
    SRMux I__2431 (
            .O(N__11114),
            .I(N__11074));
    SRMux I__2430 (
            .O(N__11113),
            .I(N__11074));
    SRMux I__2429 (
            .O(N__11112),
            .I(N__11074));
    SRMux I__2428 (
            .O(N__11111),
            .I(N__11074));
    GlobalMux I__2427 (
            .O(N__11074),
            .I(N__11071));
    gio2CtrlBuf I__2426 (
            .O(N__11071),
            .I(wPllLocked_i_g));
    CascadeMux I__2425 (
            .O(N__11068),
            .I(\fifo_inst.ftdi_output_inst.un1_oTx_n_1_sqmuxa_0_i_cascade_ ));
    CEMux I__2424 (
            .O(N__11065),
            .I(N__11062));
    LocalMux I__2423 (
            .O(N__11062),
            .I(\fifo_inst.ftdi_output_inst.un1_oTx_n_1_sqmuxa_0_i_0 ));
    InMux I__2422 (
            .O(N__11059),
            .I(N__11056));
    LocalMux I__2421 (
            .O(N__11056),
            .I(N__11051));
    InMux I__2420 (
            .O(N__11055),
            .I(N__11048));
    InMux I__2419 (
            .O(N__11054),
            .I(N__11045));
    Span4Mux_v I__2418 (
            .O(N__11051),
            .I(N__11031));
    LocalMux I__2417 (
            .O(N__11048),
            .I(N__11031));
    LocalMux I__2416 (
            .O(N__11045),
            .I(N__11031));
    InMux I__2415 (
            .O(N__11044),
            .I(N__11028));
    InMux I__2414 (
            .O(N__11043),
            .I(N__11019));
    InMux I__2413 (
            .O(N__11042),
            .I(N__11019));
    InMux I__2412 (
            .O(N__11041),
            .I(N__11019));
    InMux I__2411 (
            .O(N__11040),
            .I(N__11019));
    InMux I__2410 (
            .O(N__11039),
            .I(N__11016));
    InMux I__2409 (
            .O(N__11038),
            .I(N__11013));
    Span4Mux_v I__2408 (
            .O(N__11031),
            .I(N__11010));
    LocalMux I__2407 (
            .O(N__11028),
            .I(N__11007));
    LocalMux I__2406 (
            .O(N__11019),
            .I(N__11000));
    LocalMux I__2405 (
            .O(N__11016),
            .I(N__11000));
    LocalMux I__2404 (
            .O(N__11013),
            .I(N__11000));
    Sp12to4 I__2403 (
            .O(N__11010),
            .I(N__10997));
    Span4Mux_h I__2402 (
            .O(N__11007),
            .I(N__10994));
    Span12Mux_v I__2401 (
            .O(N__11000),
            .I(N__10991));
    Span12Mux_h I__2400 (
            .O(N__10997),
            .I(N__10986));
    Sp12to4 I__2399 (
            .O(N__10994),
            .I(N__10986));
    Span12Mux_v I__2398 (
            .O(N__10991),
            .I(N__10983));
    Span12Mux_v I__2397 (
            .O(N__10986),
            .I(N__10980));
    Odrv12 I__2396 (
            .O(N__10983),
            .I(iRxF_n_c));
    Odrv12 I__2395 (
            .O(N__10980),
            .I(iRxF_n_c));
    InMux I__2394 (
            .O(N__10975),
            .I(N__10966));
    InMux I__2393 (
            .O(N__10974),
            .I(N__10957));
    InMux I__2392 (
            .O(N__10973),
            .I(N__10957));
    InMux I__2391 (
            .O(N__10972),
            .I(N__10957));
    InMux I__2390 (
            .O(N__10971),
            .I(N__10957));
    InMux I__2389 (
            .O(N__10970),
            .I(N__10953));
    InMux I__2388 (
            .O(N__10969),
            .I(N__10950));
    LocalMux I__2387 (
            .O(N__10966),
            .I(N__10947));
    LocalMux I__2386 (
            .O(N__10957),
            .I(N__10943));
    InMux I__2385 (
            .O(N__10956),
            .I(N__10940));
    LocalMux I__2384 (
            .O(N__10953),
            .I(N__10934));
    LocalMux I__2383 (
            .O(N__10950),
            .I(N__10934));
    Span4Mux_h I__2382 (
            .O(N__10947),
            .I(N__10931));
    InMux I__2381 (
            .O(N__10946),
            .I(N__10928));
    Span4Mux_v I__2380 (
            .O(N__10943),
            .I(N__10923));
    LocalMux I__2379 (
            .O(N__10940),
            .I(N__10923));
    InMux I__2378 (
            .O(N__10939),
            .I(N__10920));
    Span4Mux_h I__2377 (
            .O(N__10934),
            .I(N__10917));
    Odrv4 I__2376 (
            .O(N__10931),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0 ));
    LocalMux I__2375 (
            .O(N__10928),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0 ));
    Odrv4 I__2374 (
            .O(N__10923),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0 ));
    LocalMux I__2373 (
            .O(N__10920),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0 ));
    Odrv4 I__2372 (
            .O(N__10917),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0 ));
    InMux I__2371 (
            .O(N__10906),
            .I(N__10903));
    LocalMux I__2370 (
            .O(N__10903),
            .I(\fifo_inst.ftdi_output_inst.N_80 ));
    CascadeMux I__2369 (
            .O(N__10900),
            .I(\DUT.uart_inst0.N_77_cascade_ ));
    InMux I__2368 (
            .O(N__10897),
            .I(N__10894));
    LocalMux I__2367 (
            .O(N__10894),
            .I(\DUT.uart_inst0.tx_state_RNI8CH01Z0Z_1 ));
    CascadeMux I__2366 (
            .O(N__10891),
            .I(\DUT.uart_inst0.tx_state_ns_i_i_o2_a0_3_0_cascade_ ));
    CascadeMux I__2365 (
            .O(N__10888),
            .I(N__10884));
    InMux I__2364 (
            .O(N__10887),
            .I(N__10880));
    InMux I__2363 (
            .O(N__10884),
            .I(N__10875));
    InMux I__2362 (
            .O(N__10883),
            .I(N__10875));
    LocalMux I__2361 (
            .O(N__10880),
            .I(\DUT.uart_inst0.N_69_i ));
    LocalMux I__2360 (
            .O(N__10875),
            .I(\DUT.uart_inst0.N_69_i ));
    CascadeMux I__2359 (
            .O(N__10870),
            .I(\DUT.uart_inst0.tx_countdown_30_3_cascade_ ));
    InMux I__2358 (
            .O(N__10867),
            .I(N__10864));
    LocalMux I__2357 (
            .O(N__10864),
            .I(N__10861));
    Span4Mux_h I__2356 (
            .O(N__10861),
            .I(N__10856));
    InMux I__2355 (
            .O(N__10860),
            .I(N__10853));
    InMux I__2354 (
            .O(N__10859),
            .I(N__10849));
    Span4Mux_v I__2353 (
            .O(N__10856),
            .I(N__10846));
    LocalMux I__2352 (
            .O(N__10853),
            .I(N__10843));
    InMux I__2351 (
            .O(N__10852),
            .I(N__10840));
    LocalMux I__2350 (
            .O(N__10849),
            .I(N__10837));
    Odrv4 I__2349 (
            .O(N__10846),
            .I(\DUT.uart_inst0.N_84 ));
    Odrv4 I__2348 (
            .O(N__10843),
            .I(\DUT.uart_inst0.N_84 ));
    LocalMux I__2347 (
            .O(N__10840),
            .I(\DUT.uart_inst0.N_84 ));
    Odrv4 I__2346 (
            .O(N__10837),
            .I(\DUT.uart_inst0.N_84 ));
    InMux I__2345 (
            .O(N__10828),
            .I(N__10822));
    InMux I__2344 (
            .O(N__10827),
            .I(N__10822));
    LocalMux I__2343 (
            .O(N__10822),
            .I(\DUT.uart_inst0.N_30_1 ));
    IoInMux I__2342 (
            .O(N__10819),
            .I(N__10816));
    LocalMux I__2341 (
            .O(N__10816),
            .I(N__10813));
    Span4Mux_s0_v I__2340 (
            .O(N__10813),
            .I(N__10810));
    Odrv4 I__2339 (
            .O(N__10810),
            .I(N_1242_i));
    IoInMux I__2338 (
            .O(N__10807),
            .I(N__10804));
    LocalMux I__2337 (
            .O(N__10804),
            .I(N__10801));
    Span4Mux_s2_v I__2336 (
            .O(N__10801),
            .I(N__10798));
    Odrv4 I__2335 (
            .O(N__10798),
            .I(N_1240_i));
    InMux I__2334 (
            .O(N__10795),
            .I(N__10792));
    LocalMux I__2333 (
            .O(N__10792),
            .I(N__10787));
    InMux I__2332 (
            .O(N__10791),
            .I(N__10784));
    InMux I__2331 (
            .O(N__10790),
            .I(N__10781));
    Odrv12 I__2330 (
            .O(N__10787),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2 ));
    LocalMux I__2329 (
            .O(N__10784),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2 ));
    LocalMux I__2328 (
            .O(N__10781),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2 ));
    CascadeMux I__2327 (
            .O(N__10774),
            .I(\fifo_inst.ftdi_output_inst.N_78_cascade_ ));
    InMux I__2326 (
            .O(N__10771),
            .I(N__10764));
    InMux I__2325 (
            .O(N__10770),
            .I(N__10759));
    InMux I__2324 (
            .O(N__10769),
            .I(N__10759));
    InMux I__2323 (
            .O(N__10768),
            .I(N__10754));
    InMux I__2322 (
            .O(N__10767),
            .I(N__10754));
    LocalMux I__2321 (
            .O(N__10764),
            .I(\DUT.uart_inst0.N_142 ));
    LocalMux I__2320 (
            .O(N__10759),
            .I(\DUT.uart_inst0.N_142 ));
    LocalMux I__2319 (
            .O(N__10754),
            .I(\DUT.uart_inst0.N_142 ));
    InMux I__2318 (
            .O(N__10747),
            .I(N__10744));
    LocalMux I__2317 (
            .O(N__10744),
            .I(\DUT.uart_inst0.N_144 ));
    CascadeMux I__2316 (
            .O(N__10741),
            .I(\DUT.uart_inst0.N_74_cascade_ ));
    CascadeMux I__2315 (
            .O(N__10738),
            .I(N__10735));
    InMux I__2314 (
            .O(N__10735),
            .I(N__10732));
    LocalMux I__2313 (
            .O(N__10732),
            .I(\DUT.uart_inst0.N_143 ));
    CascadeMux I__2312 (
            .O(N__10729),
            .I(\DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0_cascade_ ));
    InMux I__2311 (
            .O(N__10726),
            .I(N__10722));
    InMux I__2310 (
            .O(N__10725),
            .I(N__10718));
    LocalMux I__2309 (
            .O(N__10722),
            .I(N__10715));
    InMux I__2308 (
            .O(N__10721),
            .I(N__10712));
    LocalMux I__2307 (
            .O(N__10718),
            .I(\DUT.uart_inst0.N_75 ));
    Odrv4 I__2306 (
            .O(N__10715),
            .I(\DUT.uart_inst0.N_75 ));
    LocalMux I__2305 (
            .O(N__10712),
            .I(\DUT.uart_inst0.N_75 ));
    CascadeMux I__2304 (
            .O(N__10705),
            .I(\DUT.uart_inst0.N_75_cascade_ ));
    InMux I__2303 (
            .O(N__10702),
            .I(N__10699));
    LocalMux I__2302 (
            .O(N__10699),
            .I(\DUT.uart_inst0.tx_countdown_7s2_0_0 ));
    InMux I__2301 (
            .O(N__10696),
            .I(N__10687));
    InMux I__2300 (
            .O(N__10695),
            .I(N__10687));
    InMux I__2299 (
            .O(N__10694),
            .I(N__10687));
    LocalMux I__2298 (
            .O(N__10687),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_2 ));
    CascadeMux I__2297 (
            .O(N__10684),
            .I(N__10679));
    CascadeMux I__2296 (
            .O(N__10683),
            .I(N__10676));
    InMux I__2295 (
            .O(N__10682),
            .I(N__10666));
    InMux I__2294 (
            .O(N__10679),
            .I(N__10666));
    InMux I__2293 (
            .O(N__10676),
            .I(N__10666));
    InMux I__2292 (
            .O(N__10675),
            .I(N__10666));
    LocalMux I__2291 (
            .O(N__10666),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_1 ));
    InMux I__2290 (
            .O(N__10663),
            .I(N__10648));
    InMux I__2289 (
            .O(N__10662),
            .I(N__10648));
    InMux I__2288 (
            .O(N__10661),
            .I(N__10648));
    InMux I__2287 (
            .O(N__10660),
            .I(N__10648));
    InMux I__2286 (
            .O(N__10659),
            .I(N__10648));
    LocalMux I__2285 (
            .O(N__10648),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_0 ));
    CascadeMux I__2284 (
            .O(N__10645),
            .I(\DUT.uart_inst0.N_142_cascade_ ));
    CascadeMux I__2283 (
            .O(N__10642),
            .I(N__10635));
    InMux I__2282 (
            .O(N__10641),
            .I(N__10630));
    CascadeMux I__2281 (
            .O(N__10640),
            .I(N__10627));
    IoInMux I__2280 (
            .O(N__10639),
            .I(N__10622));
    InMux I__2279 (
            .O(N__10638),
            .I(N__10619));
    InMux I__2278 (
            .O(N__10635),
            .I(N__10616));
    InMux I__2277 (
            .O(N__10634),
            .I(N__10613));
    InMux I__2276 (
            .O(N__10633),
            .I(N__10610));
    LocalMux I__2275 (
            .O(N__10630),
            .I(N__10607));
    InMux I__2274 (
            .O(N__10627),
            .I(N__10604));
    CascadeMux I__2273 (
            .O(N__10626),
            .I(N__10601));
    InMux I__2272 (
            .O(N__10625),
            .I(N__10598));
    LocalMux I__2271 (
            .O(N__10622),
            .I(N__10595));
    LocalMux I__2270 (
            .O(N__10619),
            .I(N__10592));
    LocalMux I__2269 (
            .O(N__10616),
            .I(N__10585));
    LocalMux I__2268 (
            .O(N__10613),
            .I(N__10585));
    LocalMux I__2267 (
            .O(N__10610),
            .I(N__10585));
    Span4Mux_v I__2266 (
            .O(N__10607),
            .I(N__10582));
    LocalMux I__2265 (
            .O(N__10604),
            .I(N__10579));
    InMux I__2264 (
            .O(N__10601),
            .I(N__10576));
    LocalMux I__2263 (
            .O(N__10598),
            .I(N__10573));
    Span4Mux_s1_v I__2262 (
            .O(N__10595),
            .I(N__10570));
    Span4Mux_v I__2261 (
            .O(N__10592),
            .I(N__10567));
    Span4Mux_v I__2260 (
            .O(N__10585),
            .I(N__10564));
    Span4Mux_h I__2259 (
            .O(N__10582),
            .I(N__10559));
    Span4Mux_v I__2258 (
            .O(N__10579),
            .I(N__10559));
    LocalMux I__2257 (
            .O(N__10576),
            .I(N__10556));
    Span4Mux_v I__2256 (
            .O(N__10573),
            .I(N__10553));
    Span4Mux_v I__2255 (
            .O(N__10570),
            .I(N__10546));
    Span4Mux_h I__2254 (
            .O(N__10567),
            .I(N__10546));
    Span4Mux_h I__2253 (
            .O(N__10564),
            .I(N__10546));
    Span4Mux_h I__2252 (
            .O(N__10559),
            .I(N__10543));
    Sp12to4 I__2251 (
            .O(N__10556),
            .I(N__10540));
    Span4Mux_h I__2250 (
            .O(N__10553),
            .I(N__10537));
    Sp12to4 I__2249 (
            .O(N__10546),
            .I(N__10532));
    Sp12to4 I__2248 (
            .O(N__10543),
            .I(N__10532));
    Span12Mux_v I__2247 (
            .O(N__10540),
            .I(N__10529));
    Sp12to4 I__2246 (
            .O(N__10537),
            .I(N__10526));
    Span12Mux_h I__2245 (
            .O(N__10532),
            .I(N__10523));
    Span12Mux_h I__2244 (
            .O(N__10529),
            .I(N__10520));
    Span12Mux_v I__2243 (
            .O(N__10526),
            .I(N__10517));
    Span12Mux_v I__2242 (
            .O(N__10523),
            .I(N__10514));
    Span12Mux_v I__2241 (
            .O(N__10520),
            .I(N__10509));
    Span12Mux_h I__2240 (
            .O(N__10517),
            .I(N__10509));
    Odrv12 I__2239 (
            .O(N__10514),
            .I(wPllLocked));
    Odrv12 I__2238 (
            .O(N__10509),
            .I(wPllLocked));
    CascadeMux I__2237 (
            .O(N__10504),
            .I(\DUT.uart_inst0.N_84_cascade_ ));
    CascadeMux I__2236 (
            .O(N__10501),
            .I(N__10498));
    InMux I__2235 (
            .O(N__10498),
            .I(N__10486));
    InMux I__2234 (
            .O(N__10497),
            .I(N__10486));
    InMux I__2233 (
            .O(N__10496),
            .I(N__10486));
    InMux I__2232 (
            .O(N__10495),
            .I(N__10486));
    LocalMux I__2231 (
            .O(N__10486),
            .I(N__10483));
    Odrv4 I__2230 (
            .O(N__10483),
            .I(\DUT.uart_inst0.N_22 ));
    CascadeMux I__2229 (
            .O(N__10480),
            .I(\DUT.uart_inst0.N_22_cascade_ ));
    InMux I__2228 (
            .O(N__10477),
            .I(N__10474));
    LocalMux I__2227 (
            .O(N__10474),
            .I(\DUT.uart_inst0.un1_tx_bits_remaining_c3 ));
    CascadeMux I__2226 (
            .O(N__10471),
            .I(N__10467));
    InMux I__2225 (
            .O(N__10470),
            .I(N__10464));
    InMux I__2224 (
            .O(N__10467),
            .I(N__10461));
    LocalMux I__2223 (
            .O(N__10464),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_3 ));
    LocalMux I__2222 (
            .O(N__10461),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_3 ));
    InMux I__2221 (
            .O(N__10456),
            .I(N__10453));
    LocalMux I__2220 (
            .O(N__10453),
            .I(N__10447));
    InMux I__2219 (
            .O(N__10452),
            .I(N__10444));
    InMux I__2218 (
            .O(N__10451),
            .I(N__10439));
    InMux I__2217 (
            .O(N__10450),
            .I(N__10439));
    Odrv12 I__2216 (
            .O(N__10447),
            .I(rRxReadZ0));
    LocalMux I__2215 (
            .O(N__10444),
            .I(rRxReadZ0));
    LocalMux I__2214 (
            .O(N__10439),
            .I(rRxReadZ0));
    InMux I__2213 (
            .O(N__10432),
            .I(N__10429));
    LocalMux I__2212 (
            .O(N__10429),
            .I(N__10425));
    InMux I__2211 (
            .O(N__10428),
            .I(N__10422));
    Odrv12 I__2210 (
            .O(N__10425),
            .I(\DUT.fifo_rx_inst.N_206 ));
    LocalMux I__2209 (
            .O(N__10422),
            .I(\DUT.fifo_rx_inst.N_206 ));
    CascadeMux I__2208 (
            .O(N__10417),
            .I(N__10414));
    InMux I__2207 (
            .O(N__10414),
            .I(N__10409));
    CascadeMux I__2206 (
            .O(N__10413),
            .I(N__10405));
    InMux I__2205 (
            .O(N__10412),
            .I(N__10400));
    LocalMux I__2204 (
            .O(N__10409),
            .I(N__10397));
    InMux I__2203 (
            .O(N__10408),
            .I(N__10392));
    InMux I__2202 (
            .O(N__10405),
            .I(N__10392));
    InMux I__2201 (
            .O(N__10404),
            .I(N__10389));
    InMux I__2200 (
            .O(N__10403),
            .I(N__10386));
    LocalMux I__2199 (
            .O(N__10400),
            .I(N__10377));
    Span4Mux_v I__2198 (
            .O(N__10397),
            .I(N__10377));
    LocalMux I__2197 (
            .O(N__10392),
            .I(N__10377));
    LocalMux I__2196 (
            .O(N__10389),
            .I(N__10377));
    LocalMux I__2195 (
            .O(N__10386),
            .I(N__10372));
    Span4Mux_h I__2194 (
            .O(N__10377),
            .I(N__10372));
    Odrv4 I__2193 (
            .O(N__10372),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_0 ));
    InMux I__2192 (
            .O(N__10369),
            .I(N__10364));
    InMux I__2191 (
            .O(N__10368),
            .I(N__10359));
    InMux I__2190 (
            .O(N__10367),
            .I(N__10359));
    LocalMux I__2189 (
            .O(N__10364),
            .I(N__10356));
    LocalMux I__2188 (
            .O(N__10359),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1 ));
    Odrv12 I__2187 (
            .O(N__10356),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1 ));
    IoInMux I__2186 (
            .O(N__10351),
            .I(N__10348));
    LocalMux I__2185 (
            .O(N__10348),
            .I(N__10344));
    CascadeMux I__2184 (
            .O(N__10347),
            .I(N__10337));
    Span4Mux_s2_v I__2183 (
            .O(N__10344),
            .I(N__10330));
    InMux I__2182 (
            .O(N__10343),
            .I(N__10323));
    InMux I__2181 (
            .O(N__10342),
            .I(N__10323));
    InMux I__2180 (
            .O(N__10341),
            .I(N__10323));
    InMux I__2179 (
            .O(N__10340),
            .I(N__10316));
    InMux I__2178 (
            .O(N__10337),
            .I(N__10316));
    InMux I__2177 (
            .O(N__10336),
            .I(N__10309));
    InMux I__2176 (
            .O(N__10335),
            .I(N__10309));
    InMux I__2175 (
            .O(N__10334),
            .I(N__10309));
    InMux I__2174 (
            .O(N__10333),
            .I(N__10306));
    Sp12to4 I__2173 (
            .O(N__10330),
            .I(N__10303));
    LocalMux I__2172 (
            .O(N__10323),
            .I(N__10298));
    InMux I__2171 (
            .O(N__10322),
            .I(N__10295));
    InMux I__2170 (
            .O(N__10321),
            .I(N__10292));
    LocalMux I__2169 (
            .O(N__10316),
            .I(N__10285));
    LocalMux I__2168 (
            .O(N__10309),
            .I(N__10285));
    LocalMux I__2167 (
            .O(N__10306),
            .I(N__10285));
    Span12Mux_h I__2166 (
            .O(N__10303),
            .I(N__10282));
    InMux I__2165 (
            .O(N__10302),
            .I(N__10279));
    InMux I__2164 (
            .O(N__10301),
            .I(N__10276));
    Span12Mux_h I__2163 (
            .O(N__10298),
            .I(N__10273));
    LocalMux I__2162 (
            .O(N__10295),
            .I(N__10270));
    LocalMux I__2161 (
            .O(N__10292),
            .I(N__10265));
    Span4Mux_v I__2160 (
            .O(N__10285),
            .I(N__10265));
    Odrv12 I__2159 (
            .O(N__10282),
            .I(P1A2_c));
    LocalMux I__2158 (
            .O(N__10279),
            .I(P1A2_c));
    LocalMux I__2157 (
            .O(N__10276),
            .I(P1A2_c));
    Odrv12 I__2156 (
            .O(N__10273),
            .I(P1A2_c));
    Odrv12 I__2155 (
            .O(N__10270),
            .I(P1A2_c));
    Odrv4 I__2154 (
            .O(N__10265),
            .I(P1A2_c));
    CascadeMux I__2153 (
            .O(N__10252),
            .I(N__10248));
    InMux I__2152 (
            .O(N__10251),
            .I(N__10245));
    InMux I__2151 (
            .O(N__10248),
            .I(N__10242));
    LocalMux I__2150 (
            .O(N__10245),
            .I(N__10239));
    LocalMux I__2149 (
            .O(N__10242),
            .I(N__10234));
    Span4Mux_v I__2148 (
            .O(N__10239),
            .I(N__10234));
    Span4Mux_h I__2147 (
            .O(N__10234),
            .I(N__10230));
    InMux I__2146 (
            .O(N__10233),
            .I(N__10227));
    Odrv4 I__2145 (
            .O(N__10230),
            .I(rFifoCount_RNIHH0D1_0));
    LocalMux I__2144 (
            .O(N__10227),
            .I(rFifoCount_RNIHH0D1_0));
    InMux I__2143 (
            .O(N__10222),
            .I(N__10219));
    LocalMux I__2142 (
            .O(N__10219),
            .I(N__10214));
    InMux I__2141 (
            .O(N__10218),
            .I(N__10211));
    InMux I__2140 (
            .O(N__10217),
            .I(N__10208));
    Span4Mux_h I__2139 (
            .O(N__10214),
            .I(N__10201));
    LocalMux I__2138 (
            .O(N__10211),
            .I(N__10201));
    LocalMux I__2137 (
            .O(N__10208),
            .I(N__10201));
    Span4Mux_v I__2136 (
            .O(N__10201),
            .I(N__10198));
    Odrv4 I__2135 (
            .O(N__10198),
            .I(rTxWriteZ0));
    IoInMux I__2134 (
            .O(N__10195),
            .I(N__10192));
    LocalMux I__2133 (
            .O(N__10192),
            .I(N__10189));
    IoSpan4Mux I__2132 (
            .O(N__10189),
            .I(N__10186));
    Span4Mux_s3_v I__2131 (
            .O(N__10186),
            .I(N__10183));
    Span4Mux_h I__2130 (
            .O(N__10183),
            .I(N__10179));
    IoInMux I__2129 (
            .O(N__10182),
            .I(N__10176));
    Span4Mux_h I__2128 (
            .O(N__10179),
            .I(N__10172));
    LocalMux I__2127 (
            .O(N__10176),
            .I(N__10169));
    InMux I__2126 (
            .O(N__10175),
            .I(N__10166));
    Odrv4 I__2125 (
            .O(N__10172),
            .I(P1A3_c));
    Odrv12 I__2124 (
            .O(N__10169),
            .I(P1A3_c));
    LocalMux I__2123 (
            .O(N__10166),
            .I(P1A3_c));
    InMux I__2122 (
            .O(N__10159),
            .I(N__10155));
    InMux I__2121 (
            .O(N__10158),
            .I(N__10152));
    LocalMux I__2120 (
            .O(N__10155),
            .I(N__10148));
    LocalMux I__2119 (
            .O(N__10152),
            .I(N__10145));
    InMux I__2118 (
            .O(N__10151),
            .I(N__10142));
    Span4Mux_h I__2117 (
            .O(N__10148),
            .I(N__10134));
    Span4Mux_v I__2116 (
            .O(N__10145),
            .I(N__10134));
    LocalMux I__2115 (
            .O(N__10142),
            .I(N__10134));
    InMux I__2114 (
            .O(N__10141),
            .I(N__10131));
    Odrv4 I__2113 (
            .O(N__10134),
            .I(rTxByteZ0Z_2));
    LocalMux I__2112 (
            .O(N__10131),
            .I(rTxByteZ0Z_2));
    InMux I__2111 (
            .O(N__10126),
            .I(N__10123));
    LocalMux I__2110 (
            .O(N__10123),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_2 ));
    InMux I__2109 (
            .O(N__10120),
            .I(N__10117));
    LocalMux I__2108 (
            .O(N__10117),
            .I(N__10113));
    InMux I__2107 (
            .O(N__10116),
            .I(N__10109));
    Span4Mux_v I__2106 (
            .O(N__10113),
            .I(N__10106));
    InMux I__2105 (
            .O(N__10112),
            .I(N__10103));
    LocalMux I__2104 (
            .O(N__10109),
            .I(N__10095));
    Sp12to4 I__2103 (
            .O(N__10106),
            .I(N__10095));
    LocalMux I__2102 (
            .O(N__10103),
            .I(N__10095));
    InMux I__2101 (
            .O(N__10102),
            .I(N__10092));
    Odrv12 I__2100 (
            .O(N__10095),
            .I(rTxByteZ0Z_7));
    LocalMux I__2099 (
            .O(N__10092),
            .I(rTxByteZ0Z_7));
    InMux I__2098 (
            .O(N__10087),
            .I(N__10084));
    LocalMux I__2097 (
            .O(N__10084),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_7 ));
    CEMux I__2096 (
            .O(N__10081),
            .I(N__10075));
    CEMux I__2095 (
            .O(N__10080),
            .I(N__10072));
    CEMux I__2094 (
            .O(N__10079),
            .I(N__10068));
    CEMux I__2093 (
            .O(N__10078),
            .I(N__10065));
    LocalMux I__2092 (
            .O(N__10075),
            .I(N__10062));
    LocalMux I__2091 (
            .O(N__10072),
            .I(N__10058));
    CEMux I__2090 (
            .O(N__10071),
            .I(N__10055));
    LocalMux I__2089 (
            .O(N__10068),
            .I(N__10052));
    LocalMux I__2088 (
            .O(N__10065),
            .I(N__10049));
    Span4Mux_v I__2087 (
            .O(N__10062),
            .I(N__10046));
    CEMux I__2086 (
            .O(N__10061),
            .I(N__10043));
    Span4Mux_v I__2085 (
            .O(N__10058),
            .I(N__10038));
    LocalMux I__2084 (
            .O(N__10055),
            .I(N__10038));
    Span4Mux_v I__2083 (
            .O(N__10052),
            .I(N__10033));
    Span4Mux_h I__2082 (
            .O(N__10049),
            .I(N__10033));
    Sp12to4 I__2081 (
            .O(N__10046),
            .I(N__10028));
    LocalMux I__2080 (
            .O(N__10043),
            .I(N__10028));
    Span4Mux_h I__2079 (
            .O(N__10038),
            .I(N__10024));
    Sp12to4 I__2078 (
            .O(N__10033),
            .I(N__10019));
    Span12Mux_s11_h I__2077 (
            .O(N__10028),
            .I(N__10019));
    InMux I__2076 (
            .O(N__10027),
            .I(N__10016));
    Odrv4 I__2075 (
            .O(N__10024),
            .I(\DUT.fifo_tx_inst.rFifoData_awe0 ));
    Odrv12 I__2074 (
            .O(N__10019),
            .I(\DUT.fifo_tx_inst.rFifoData_awe0 ));
    LocalMux I__2073 (
            .O(N__10016),
            .I(\DUT.fifo_tx_inst.rFifoData_awe0 ));
    InMux I__2072 (
            .O(N__10009),
            .I(N__10006));
    LocalMux I__2071 (
            .O(N__10006),
            .I(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0 ));
    CascadeMux I__2070 (
            .O(N__10003),
            .I(N__9998));
    CascadeMux I__2069 (
            .O(N__10002),
            .I(N__9995));
    InMux I__2068 (
            .O(N__10001),
            .I(N__9990));
    InMux I__2067 (
            .O(N__9998),
            .I(N__9987));
    InMux I__2066 (
            .O(N__9995),
            .I(N__9980));
    InMux I__2065 (
            .O(N__9994),
            .I(N__9980));
    InMux I__2064 (
            .O(N__9993),
            .I(N__9980));
    LocalMux I__2063 (
            .O(N__9990),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_0 ));
    LocalMux I__2062 (
            .O(N__9987),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_0 ));
    LocalMux I__2061 (
            .O(N__9980),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_0 ));
    CascadeMux I__2060 (
            .O(N__9973),
            .I(N__9970));
    InMux I__2059 (
            .O(N__9970),
            .I(N__9967));
    LocalMux I__2058 (
            .O(N__9967),
            .I(\DUT.fifo_tx_inst.rFifoCount_RNISSQ21Z0Z_1 ));
    InMux I__2057 (
            .O(N__9964),
            .I(N__9958));
    InMux I__2056 (
            .O(N__9963),
            .I(N__9953));
    InMux I__2055 (
            .O(N__9962),
            .I(N__9953));
    InMux I__2054 (
            .O(N__9961),
            .I(N__9950));
    LocalMux I__2053 (
            .O(N__9958),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_1 ));
    LocalMux I__2052 (
            .O(N__9953),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_1 ));
    LocalMux I__2051 (
            .O(N__9950),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_1 ));
    InMux I__2050 (
            .O(N__9943),
            .I(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0 ));
    InMux I__2049 (
            .O(N__9940),
            .I(N__9935));
    InMux I__2048 (
            .O(N__9939),
            .I(N__9932));
    InMux I__2047 (
            .O(N__9938),
            .I(N__9929));
    LocalMux I__2046 (
            .O(N__9935),
            .I(\DUT.fifo_tx_inst.N_83 ));
    LocalMux I__2045 (
            .O(N__9932),
            .I(\DUT.fifo_tx_inst.N_83 ));
    LocalMux I__2044 (
            .O(N__9929),
            .I(\DUT.fifo_tx_inst.N_83 ));
    InMux I__2043 (
            .O(N__9922),
            .I(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1 ));
    InMux I__2042 (
            .O(N__9919),
            .I(N__9916));
    LocalMux I__2041 (
            .O(N__9916),
            .I(N__9911));
    CascadeMux I__2040 (
            .O(N__9915),
            .I(N__9907));
    InMux I__2039 (
            .O(N__9914),
            .I(N__9903));
    Span4Mux_h I__2038 (
            .O(N__9911),
            .I(N__9900));
    InMux I__2037 (
            .O(N__9910),
            .I(N__9897));
    InMux I__2036 (
            .O(N__9907),
            .I(N__9892));
    InMux I__2035 (
            .O(N__9906),
            .I(N__9892));
    LocalMux I__2034 (
            .O(N__9903),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_2 ));
    Odrv4 I__2033 (
            .O(N__9900),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_2 ));
    LocalMux I__2032 (
            .O(N__9897),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_2 ));
    LocalMux I__2031 (
            .O(N__9892),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_2 ));
    CascadeMux I__2030 (
            .O(N__9883),
            .I(N__9878));
    InMux I__2029 (
            .O(N__9882),
            .I(N__9871));
    InMux I__2028 (
            .O(N__9881),
            .I(N__9871));
    InMux I__2027 (
            .O(N__9878),
            .I(N__9871));
    LocalMux I__2026 (
            .O(N__9871),
            .I(N__9866));
    InMux I__2025 (
            .O(N__9870),
            .I(N__9863));
    CascadeMux I__2024 (
            .O(N__9869),
            .I(N__9857));
    Span4Mux_v I__2023 (
            .O(N__9866),
            .I(N__9852));
    LocalMux I__2022 (
            .O(N__9863),
            .I(N__9849));
    InMux I__2021 (
            .O(N__9862),
            .I(N__9844));
    InMux I__2020 (
            .O(N__9861),
            .I(N__9844));
    InMux I__2019 (
            .O(N__9860),
            .I(N__9839));
    InMux I__2018 (
            .O(N__9857),
            .I(N__9839));
    CascadeMux I__2017 (
            .O(N__9856),
            .I(N__9836));
    InMux I__2016 (
            .O(N__9855),
            .I(N__9833));
    Span4Mux_h I__2015 (
            .O(N__9852),
            .I(N__9824));
    Span4Mux_s2_v I__2014 (
            .O(N__9849),
            .I(N__9824));
    LocalMux I__2013 (
            .O(N__9844),
            .I(N__9824));
    LocalMux I__2012 (
            .O(N__9839),
            .I(N__9824));
    InMux I__2011 (
            .O(N__9836),
            .I(N__9821));
    LocalMux I__2010 (
            .O(N__9833),
            .I(N__9818));
    Span4Mux_h I__2009 (
            .O(N__9824),
            .I(N__9813));
    LocalMux I__2008 (
            .O(N__9821),
            .I(N__9813));
    Span12Mux_h I__2007 (
            .O(N__9818),
            .I(N__9810));
    IoSpan4Mux I__2006 (
            .O(N__9813),
            .I(N__9807));
    Odrv12 I__2005 (
            .O(N__9810),
            .I(P1A1_c));
    Odrv4 I__2004 (
            .O(N__9807),
            .I(P1A1_c));
    InMux I__2003 (
            .O(N__9802),
            .I(N__9797));
    InMux I__2002 (
            .O(N__9801),
            .I(N__9794));
    InMux I__2001 (
            .O(N__9800),
            .I(N__9791));
    LocalMux I__2000 (
            .O(N__9797),
            .I(\DUT.uart_inst0.recv_stateZ0Z_3 ));
    LocalMux I__1999 (
            .O(N__9794),
            .I(\DUT.uart_inst0.recv_stateZ0Z_3 ));
    LocalMux I__1998 (
            .O(N__9791),
            .I(\DUT.uart_inst0.recv_stateZ0Z_3 ));
    InMux I__1997 (
            .O(N__9784),
            .I(N__9781));
    LocalMux I__1996 (
            .O(N__9781),
            .I(N__9778));
    Span4Mux_h I__1995 (
            .O(N__9778),
            .I(N__9775));
    Odrv4 I__1994 (
            .O(N__9775),
            .I(\DUT.uart_inst0.g0_1 ));
    InMux I__1993 (
            .O(N__9772),
            .I(N__9765));
    InMux I__1992 (
            .O(N__9771),
            .I(N__9765));
    InMux I__1991 (
            .O(N__9770),
            .I(N__9762));
    LocalMux I__1990 (
            .O(N__9765),
            .I(N__9756));
    LocalMux I__1989 (
            .O(N__9762),
            .I(N__9753));
    InMux I__1988 (
            .O(N__9761),
            .I(N__9748));
    InMux I__1987 (
            .O(N__9760),
            .I(N__9748));
    InMux I__1986 (
            .O(N__9759),
            .I(N__9743));
    Span4Mux_s2_v I__1985 (
            .O(N__9756),
            .I(N__9738));
    Span4Mux_h I__1984 (
            .O(N__9753),
            .I(N__9738));
    LocalMux I__1983 (
            .O(N__9748),
            .I(N__9735));
    InMux I__1982 (
            .O(N__9747),
            .I(N__9730));
    InMux I__1981 (
            .O(N__9746),
            .I(N__9730));
    LocalMux I__1980 (
            .O(N__9743),
            .I(\DUT.uart_inst0.recv_stateZ0Z_5 ));
    Odrv4 I__1979 (
            .O(N__9738),
            .I(\DUT.uart_inst0.recv_stateZ0Z_5 ));
    Odrv4 I__1978 (
            .O(N__9735),
            .I(\DUT.uart_inst0.recv_stateZ0Z_5 ));
    LocalMux I__1977 (
            .O(N__9730),
            .I(\DUT.uart_inst0.recv_stateZ0Z_5 ));
    InMux I__1976 (
            .O(N__9721),
            .I(N__9717));
    CascadeMux I__1975 (
            .O(N__9720),
            .I(N__9708));
    LocalMux I__1974 (
            .O(N__9717),
            .I(N__9702));
    InMux I__1973 (
            .O(N__9716),
            .I(N__9697));
    InMux I__1972 (
            .O(N__9715),
            .I(N__9697));
    InMux I__1971 (
            .O(N__9714),
            .I(N__9694));
    InMux I__1970 (
            .O(N__9713),
            .I(N__9689));
    InMux I__1969 (
            .O(N__9712),
            .I(N__9689));
    InMux I__1968 (
            .O(N__9711),
            .I(N__9682));
    InMux I__1967 (
            .O(N__9708),
            .I(N__9682));
    InMux I__1966 (
            .O(N__9707),
            .I(N__9682));
    InMux I__1965 (
            .O(N__9706),
            .I(N__9677));
    InMux I__1964 (
            .O(N__9705),
            .I(N__9677));
    Odrv4 I__1963 (
            .O(N__9702),
            .I(\DUT.uart_inst0.rx_countdown_3_4 ));
    LocalMux I__1962 (
            .O(N__9697),
            .I(\DUT.uart_inst0.rx_countdown_3_4 ));
    LocalMux I__1961 (
            .O(N__9694),
            .I(\DUT.uart_inst0.rx_countdown_3_4 ));
    LocalMux I__1960 (
            .O(N__9689),
            .I(\DUT.uart_inst0.rx_countdown_3_4 ));
    LocalMux I__1959 (
            .O(N__9682),
            .I(\DUT.uart_inst0.rx_countdown_3_4 ));
    LocalMux I__1958 (
            .O(N__9677),
            .I(\DUT.uart_inst0.rx_countdown_3_4 ));
    CascadeMux I__1957 (
            .O(N__9664),
            .I(N__9661));
    InMux I__1956 (
            .O(N__9661),
            .I(N__9658));
    LocalMux I__1955 (
            .O(N__9658),
            .I(N__9655));
    Odrv4 I__1954 (
            .O(N__9655),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_4 ));
    InMux I__1953 (
            .O(N__9652),
            .I(N__9647));
    InMux I__1952 (
            .O(N__9651),
            .I(N__9644));
    InMux I__1951 (
            .O(N__9650),
            .I(N__9641));
    LocalMux I__1950 (
            .O(N__9647),
            .I(N__9634));
    LocalMux I__1949 (
            .O(N__9644),
            .I(N__9634));
    LocalMux I__1948 (
            .O(N__9641),
            .I(N__9631));
    InMux I__1947 (
            .O(N__9640),
            .I(N__9620));
    InMux I__1946 (
            .O(N__9639),
            .I(N__9620));
    Span4Mux_s2_v I__1945 (
            .O(N__9634),
            .I(N__9617));
    Span4Mux_v I__1944 (
            .O(N__9631),
            .I(N__9614));
    InMux I__1943 (
            .O(N__9630),
            .I(N__9607));
    InMux I__1942 (
            .O(N__9629),
            .I(N__9607));
    InMux I__1941 (
            .O(N__9628),
            .I(N__9607));
    InMux I__1940 (
            .O(N__9627),
            .I(N__9602));
    InMux I__1939 (
            .O(N__9626),
            .I(N__9602));
    InMux I__1938 (
            .O(N__9625),
            .I(N__9599));
    LocalMux I__1937 (
            .O(N__9620),
            .I(\DUT.uart_inst0.rx_countdown_3_5 ));
    Odrv4 I__1936 (
            .O(N__9617),
            .I(\DUT.uart_inst0.rx_countdown_3_5 ));
    Odrv4 I__1935 (
            .O(N__9614),
            .I(\DUT.uart_inst0.rx_countdown_3_5 ));
    LocalMux I__1934 (
            .O(N__9607),
            .I(\DUT.uart_inst0.rx_countdown_3_5 ));
    LocalMux I__1933 (
            .O(N__9602),
            .I(\DUT.uart_inst0.rx_countdown_3_5 ));
    LocalMux I__1932 (
            .O(N__9599),
            .I(\DUT.uart_inst0.rx_countdown_3_5 ));
    InMux I__1931 (
            .O(N__9586),
            .I(N__9583));
    LocalMux I__1930 (
            .O(N__9583),
            .I(N__9580));
    Odrv4 I__1929 (
            .O(N__9580),
            .I(\DUT.uart_inst0.recv_state_RNO_2Z0Z_1 ));
    InMux I__1928 (
            .O(N__9577),
            .I(N__9572));
    InMux I__1927 (
            .O(N__9576),
            .I(N__9568));
    InMux I__1926 (
            .O(N__9575),
            .I(N__9565));
    LocalMux I__1925 (
            .O(N__9572),
            .I(N__9562));
    CascadeMux I__1924 (
            .O(N__9571),
            .I(N__9553));
    LocalMux I__1923 (
            .O(N__9568),
            .I(N__9548));
    LocalMux I__1922 (
            .O(N__9565),
            .I(N__9543));
    Span4Mux_h I__1921 (
            .O(N__9562),
            .I(N__9543));
    InMux I__1920 (
            .O(N__9561),
            .I(N__9536));
    InMux I__1919 (
            .O(N__9560),
            .I(N__9536));
    InMux I__1918 (
            .O(N__9559),
            .I(N__9536));
    InMux I__1917 (
            .O(N__9558),
            .I(N__9531));
    InMux I__1916 (
            .O(N__9557),
            .I(N__9531));
    InMux I__1915 (
            .O(N__9556),
            .I(N__9526));
    InMux I__1914 (
            .O(N__9553),
            .I(N__9526));
    InMux I__1913 (
            .O(N__9552),
            .I(N__9523));
    InMux I__1912 (
            .O(N__9551),
            .I(N__9520));
    Odrv4 I__1911 (
            .O(N__9548),
            .I(\DUT.uart_inst0.rx_countdown_3_0 ));
    Odrv4 I__1910 (
            .O(N__9543),
            .I(\DUT.uart_inst0.rx_countdown_3_0 ));
    LocalMux I__1909 (
            .O(N__9536),
            .I(\DUT.uart_inst0.rx_countdown_3_0 ));
    LocalMux I__1908 (
            .O(N__9531),
            .I(\DUT.uart_inst0.rx_countdown_3_0 ));
    LocalMux I__1907 (
            .O(N__9526),
            .I(\DUT.uart_inst0.rx_countdown_3_0 ));
    LocalMux I__1906 (
            .O(N__9523),
            .I(\DUT.uart_inst0.rx_countdown_3_0 ));
    LocalMux I__1905 (
            .O(N__9520),
            .I(\DUT.uart_inst0.rx_countdown_3_0 ));
    InMux I__1904 (
            .O(N__9505),
            .I(N__9500));
    CascadeMux I__1903 (
            .O(N__9504),
            .I(N__9494));
    CascadeMux I__1902 (
            .O(N__9503),
            .I(N__9491));
    LocalMux I__1901 (
            .O(N__9500),
            .I(N__9488));
    CascadeMux I__1900 (
            .O(N__9499),
            .I(N__9483));
    CascadeMux I__1899 (
            .O(N__9498),
            .I(N__9480));
    CascadeMux I__1898 (
            .O(N__9497),
            .I(N__9476));
    InMux I__1897 (
            .O(N__9494),
            .I(N__9471));
    InMux I__1896 (
            .O(N__9491),
            .I(N__9471));
    Span4Mux_h I__1895 (
            .O(N__9488),
            .I(N__9468));
    InMux I__1894 (
            .O(N__9487),
            .I(N__9465));
    InMux I__1893 (
            .O(N__9486),
            .I(N__9462));
    InMux I__1892 (
            .O(N__9483),
            .I(N__9459));
    InMux I__1891 (
            .O(N__9480),
            .I(N__9452));
    InMux I__1890 (
            .O(N__9479),
            .I(N__9452));
    InMux I__1889 (
            .O(N__9476),
            .I(N__9452));
    LocalMux I__1888 (
            .O(N__9471),
            .I(\DUT.uart_inst0.rx_countdown_3_2 ));
    Odrv4 I__1887 (
            .O(N__9468),
            .I(\DUT.uart_inst0.rx_countdown_3_2 ));
    LocalMux I__1886 (
            .O(N__9465),
            .I(\DUT.uart_inst0.rx_countdown_3_2 ));
    LocalMux I__1885 (
            .O(N__9462),
            .I(\DUT.uart_inst0.rx_countdown_3_2 ));
    LocalMux I__1884 (
            .O(N__9459),
            .I(\DUT.uart_inst0.rx_countdown_3_2 ));
    LocalMux I__1883 (
            .O(N__9452),
            .I(\DUT.uart_inst0.rx_countdown_3_2 ));
    CascadeMux I__1882 (
            .O(N__9439),
            .I(\DUT.uart_inst0.G_10_i_a4_0_4_cascade_ ));
    InMux I__1881 (
            .O(N__9436),
            .I(N__9432));
    InMux I__1880 (
            .O(N__9435),
            .I(N__9425));
    LocalMux I__1879 (
            .O(N__9432),
            .I(N__9422));
    CascadeMux I__1878 (
            .O(N__9431),
            .I(N__9413));
    CascadeMux I__1877 (
            .O(N__9430),
            .I(N__9410));
    InMux I__1876 (
            .O(N__9429),
            .I(N__9405));
    InMux I__1875 (
            .O(N__9428),
            .I(N__9405));
    LocalMux I__1874 (
            .O(N__9425),
            .I(N__9400));
    Span4Mux_h I__1873 (
            .O(N__9422),
            .I(N__9400));
    InMux I__1872 (
            .O(N__9421),
            .I(N__9397));
    InMux I__1871 (
            .O(N__9420),
            .I(N__9388));
    InMux I__1870 (
            .O(N__9419),
            .I(N__9388));
    InMux I__1869 (
            .O(N__9418),
            .I(N__9388));
    InMux I__1868 (
            .O(N__9417),
            .I(N__9388));
    InMux I__1867 (
            .O(N__9416),
            .I(N__9385));
    InMux I__1866 (
            .O(N__9413),
            .I(N__9380));
    InMux I__1865 (
            .O(N__9410),
            .I(N__9380));
    LocalMux I__1864 (
            .O(N__9405),
            .I(\DUT.uart_inst0.rx_countdown_3_3 ));
    Odrv4 I__1863 (
            .O(N__9400),
            .I(\DUT.uart_inst0.rx_countdown_3_3 ));
    LocalMux I__1862 (
            .O(N__9397),
            .I(\DUT.uart_inst0.rx_countdown_3_3 ));
    LocalMux I__1861 (
            .O(N__9388),
            .I(\DUT.uart_inst0.rx_countdown_3_3 ));
    LocalMux I__1860 (
            .O(N__9385),
            .I(\DUT.uart_inst0.rx_countdown_3_3 ));
    LocalMux I__1859 (
            .O(N__9380),
            .I(\DUT.uart_inst0.rx_countdown_3_3 ));
    CascadeMux I__1858 (
            .O(N__9367),
            .I(\DUT.uart_inst0.N_4_i_0_1_cascade_ ));
    InMux I__1857 (
            .O(N__9364),
            .I(N__9355));
    InMux I__1856 (
            .O(N__9363),
            .I(N__9355));
    InMux I__1855 (
            .O(N__9362),
            .I(N__9355));
    LocalMux I__1854 (
            .O(N__9355),
            .I(N__9343));
    InMux I__1853 (
            .O(N__9354),
            .I(N__9332));
    InMux I__1852 (
            .O(N__9353),
            .I(N__9332));
    InMux I__1851 (
            .O(N__9352),
            .I(N__9332));
    InMux I__1850 (
            .O(N__9351),
            .I(N__9332));
    InMux I__1849 (
            .O(N__9350),
            .I(N__9332));
    InMux I__1848 (
            .O(N__9349),
            .I(N__9327));
    InMux I__1847 (
            .O(N__9348),
            .I(N__9327));
    CascadeMux I__1846 (
            .O(N__9347),
            .I(N__9324));
    CascadeMux I__1845 (
            .O(N__9346),
            .I(N__9321));
    Span4Mux_s2_v I__1844 (
            .O(N__9343),
            .I(N__9305));
    LocalMux I__1843 (
            .O(N__9332),
            .I(N__9300));
    LocalMux I__1842 (
            .O(N__9327),
            .I(N__9300));
    InMux I__1841 (
            .O(N__9324),
            .I(N__9287));
    InMux I__1840 (
            .O(N__9321),
            .I(N__9287));
    InMux I__1839 (
            .O(N__9320),
            .I(N__9287));
    InMux I__1838 (
            .O(N__9319),
            .I(N__9287));
    InMux I__1837 (
            .O(N__9318),
            .I(N__9287));
    InMux I__1836 (
            .O(N__9317),
            .I(N__9287));
    InMux I__1835 (
            .O(N__9316),
            .I(N__9284));
    InMux I__1834 (
            .O(N__9315),
            .I(N__9281));
    InMux I__1833 (
            .O(N__9314),
            .I(N__9278));
    InMux I__1832 (
            .O(N__9313),
            .I(N__9271));
    InMux I__1831 (
            .O(N__9312),
            .I(N__9271));
    InMux I__1830 (
            .O(N__9311),
            .I(N__9271));
    InMux I__1829 (
            .O(N__9310),
            .I(N__9264));
    InMux I__1828 (
            .O(N__9309),
            .I(N__9264));
    InMux I__1827 (
            .O(N__9308),
            .I(N__9264));
    Span4Mux_h I__1826 (
            .O(N__9305),
            .I(N__9259));
    Span4Mux_s2_v I__1825 (
            .O(N__9300),
            .I(N__9259));
    LocalMux I__1824 (
            .O(N__9287),
            .I(N__9254));
    LocalMux I__1823 (
            .O(N__9284),
            .I(N__9254));
    LocalMux I__1822 (
            .O(N__9281),
            .I(\DUT.uart_inst0.N_149 ));
    LocalMux I__1821 (
            .O(N__9278),
            .I(\DUT.uart_inst0.N_149 ));
    LocalMux I__1820 (
            .O(N__9271),
            .I(\DUT.uart_inst0.N_149 ));
    LocalMux I__1819 (
            .O(N__9264),
            .I(\DUT.uart_inst0.N_149 ));
    Odrv4 I__1818 (
            .O(N__9259),
            .I(\DUT.uart_inst0.N_149 ));
    Odrv4 I__1817 (
            .O(N__9254),
            .I(\DUT.uart_inst0.N_149 ));
    InMux I__1816 (
            .O(N__9241),
            .I(N__9238));
    LocalMux I__1815 (
            .O(N__9238),
            .I(N__9231));
    InMux I__1814 (
            .O(N__9237),
            .I(N__9224));
    InMux I__1813 (
            .O(N__9236),
            .I(N__9224));
    InMux I__1812 (
            .O(N__9235),
            .I(N__9224));
    InMux I__1811 (
            .O(N__9234),
            .I(N__9216));
    Span4Mux_h I__1810 (
            .O(N__9231),
            .I(N__9213));
    LocalMux I__1809 (
            .O(N__9224),
            .I(N__9210));
    InMux I__1808 (
            .O(N__9223),
            .I(N__9205));
    InMux I__1807 (
            .O(N__9222),
            .I(N__9205));
    InMux I__1806 (
            .O(N__9221),
            .I(N__9198));
    InMux I__1805 (
            .O(N__9220),
            .I(N__9198));
    InMux I__1804 (
            .O(N__9219),
            .I(N__9198));
    LocalMux I__1803 (
            .O(N__9216),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    Odrv4 I__1802 (
            .O(N__9213),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    Odrv4 I__1801 (
            .O(N__9210),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    LocalMux I__1800 (
            .O(N__9205),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    LocalMux I__1799 (
            .O(N__9198),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    InMux I__1798 (
            .O(N__9187),
            .I(N__9184));
    LocalMux I__1797 (
            .O(N__9184),
            .I(\DUT.rFifoDatarx_4 ));
    CascadeMux I__1796 (
            .O(N__9181),
            .I(N__9178));
    InMux I__1795 (
            .O(N__9178),
            .I(N__9175));
    LocalMux I__1794 (
            .O(N__9175),
            .I(\DUT.uart_inst0.tx_dataZ0Z_5 ));
    CascadeMux I__1793 (
            .O(N__9172),
            .I(N__9169));
    InMux I__1792 (
            .O(N__9169),
            .I(N__9166));
    LocalMux I__1791 (
            .O(N__9166),
            .I(N__9163));
    Odrv12 I__1790 (
            .O(N__9163),
            .I(\DUT.uart_inst0.tx_dataZ0Z_4 ));
    InMux I__1789 (
            .O(N__9160),
            .I(N__9157));
    LocalMux I__1788 (
            .O(N__9157),
            .I(\DUT.rFifoDatarx_7 ));
    CascadeMux I__1787 (
            .O(N__9154),
            .I(N__9150));
    InMux I__1786 (
            .O(N__9153),
            .I(N__9139));
    InMux I__1785 (
            .O(N__9150),
            .I(N__9139));
    InMux I__1784 (
            .O(N__9149),
            .I(N__9139));
    InMux I__1783 (
            .O(N__9148),
            .I(N__9139));
    LocalMux I__1782 (
            .O(N__9139),
            .I(N__9132));
    InMux I__1781 (
            .O(N__9138),
            .I(N__9123));
    InMux I__1780 (
            .O(N__9137),
            .I(N__9123));
    InMux I__1779 (
            .O(N__9136),
            .I(N__9123));
    InMux I__1778 (
            .O(N__9135),
            .I(N__9123));
    Odrv4 I__1777 (
            .O(N__9132),
            .I(\DUT.uart_inst0.N_145 ));
    LocalMux I__1776 (
            .O(N__9123),
            .I(\DUT.uart_inst0.N_145 ));
    CascadeMux I__1775 (
            .O(N__9118),
            .I(N__9115));
    InMux I__1774 (
            .O(N__9115),
            .I(N__9112));
    LocalMux I__1773 (
            .O(N__9112),
            .I(\DUT.uart_inst0.tx_dataZ0Z_7 ));
    CEMux I__1772 (
            .O(N__9109),
            .I(N__9106));
    LocalMux I__1771 (
            .O(N__9106),
            .I(N__9103));
    Span4Mux_v I__1770 (
            .O(N__9103),
            .I(N__9099));
    CEMux I__1769 (
            .O(N__9102),
            .I(N__9096));
    Span4Mux_h I__1768 (
            .O(N__9099),
            .I(N__9093));
    LocalMux I__1767 (
            .O(N__9096),
            .I(N__9090));
    Odrv4 I__1766 (
            .O(N__9093),
            .I(\DUT.uart_inst0.N_22_i ));
    Odrv12 I__1765 (
            .O(N__9090),
            .I(\DUT.uart_inst0.N_22_i ));
    CascadeMux I__1764 (
            .O(N__9085),
            .I(\DUT.fifo_tx_inst.N_83_cascade_ ));
    InMux I__1763 (
            .O(N__9082),
            .I(N__9078));
    CascadeMux I__1762 (
            .O(N__9081),
            .I(N__9075));
    LocalMux I__1761 (
            .O(N__9078),
            .I(N__9072));
    InMux I__1760 (
            .O(N__9075),
            .I(N__9069));
    Odrv12 I__1759 (
            .O(N__9072),
            .I(\DUT.uart_inst0.tx_dataZ0Z_0 ));
    LocalMux I__1758 (
            .O(N__9069),
            .I(\DUT.uart_inst0.tx_dataZ0Z_0 ));
    CascadeMux I__1757 (
            .O(N__9064),
            .I(N__9061));
    InMux I__1756 (
            .O(N__9061),
            .I(N__9057));
    IoInMux I__1755 (
            .O(N__9060),
            .I(N__9054));
    LocalMux I__1754 (
            .O(N__9057),
            .I(N__9050));
    LocalMux I__1753 (
            .O(N__9054),
            .I(N__9047));
    InMux I__1752 (
            .O(N__9053),
            .I(N__9043));
    Span4Mux_h I__1751 (
            .O(N__9050),
            .I(N__9040));
    Span4Mux_s0_v I__1750 (
            .O(N__9047),
            .I(N__9037));
    CascadeMux I__1749 (
            .O(N__9046),
            .I(N__9034));
    LocalMux I__1748 (
            .O(N__9043),
            .I(N__9031));
    Span4Mux_v I__1747 (
            .O(N__9040),
            .I(N__9028));
    Span4Mux_h I__1746 (
            .O(N__9037),
            .I(N__9025));
    InMux I__1745 (
            .O(N__9034),
            .I(N__9022));
    Span12Mux_s11_h I__1744 (
            .O(N__9031),
            .I(N__9019));
    Span4Mux_v I__1743 (
            .O(N__9028),
            .I(N__9016));
    Odrv4 I__1742 (
            .O(N__9025),
            .I(P1A7_c));
    LocalMux I__1741 (
            .O(N__9022),
            .I(P1A7_c));
    Odrv12 I__1740 (
            .O(N__9019),
            .I(P1A7_c));
    Odrv4 I__1739 (
            .O(N__9016),
            .I(P1A7_c));
    CascadeMux I__1738 (
            .O(N__9007),
            .I(N__9004));
    InMux I__1737 (
            .O(N__9004),
            .I(N__9001));
    LocalMux I__1736 (
            .O(N__9001),
            .I(N__8998));
    Odrv4 I__1735 (
            .O(N__8998),
            .I(\DUT.uart_inst0.N_98 ));
    InMux I__1734 (
            .O(N__8995),
            .I(N__8992));
    LocalMux I__1733 (
            .O(N__8992),
            .I(\fifo_inst.ftdi_output_inst.rFifoStatec_0 ));
    CascadeMux I__1732 (
            .O(N__8989),
            .I(N__8986));
    InMux I__1731 (
            .O(N__8986),
            .I(N__8978));
    InMux I__1730 (
            .O(N__8985),
            .I(N__8969));
    InMux I__1729 (
            .O(N__8984),
            .I(N__8969));
    InMux I__1728 (
            .O(N__8983),
            .I(N__8969));
    InMux I__1727 (
            .O(N__8982),
            .I(N__8969));
    InMux I__1726 (
            .O(N__8981),
            .I(N__8966));
    LocalMux I__1725 (
            .O(N__8978),
            .I(\DUT.fifo_tx_inst.N_79 ));
    LocalMux I__1724 (
            .O(N__8969),
            .I(\DUT.fifo_tx_inst.N_79 ));
    LocalMux I__1723 (
            .O(N__8966),
            .I(\DUT.fifo_tx_inst.N_79 ));
    InMux I__1722 (
            .O(N__8959),
            .I(N__8956));
    LocalMux I__1721 (
            .O(N__8956),
            .I(\DUT.uart_inst0.tx_dataZ0Z_2 ));
    InMux I__1720 (
            .O(N__8953),
            .I(N__8950));
    LocalMux I__1719 (
            .O(N__8950),
            .I(\DUT.rFifoDatarx_0_3 ));
    InMux I__1718 (
            .O(N__8947),
            .I(N__8944));
    LocalMux I__1717 (
            .O(N__8944),
            .I(N__8941));
    Odrv4 I__1716 (
            .O(N__8941),
            .I(\DUT.uart_inst0.tx_dataZ0Z_3 ));
    InMux I__1715 (
            .O(N__8938),
            .I(N__8935));
    LocalMux I__1714 (
            .O(N__8935),
            .I(N__8932));
    Span4Mux_h I__1713 (
            .O(N__8932),
            .I(N__8929));
    Odrv4 I__1712 (
            .O(N__8929),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_7 ));
    InMux I__1711 (
            .O(N__8926),
            .I(N__8923));
    LocalMux I__1710 (
            .O(N__8923),
            .I(N__8920));
    Odrv4 I__1709 (
            .O(N__8920),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_7 ));
    CascadeMux I__1708 (
            .O(N__8917),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_ ));
    InMux I__1707 (
            .O(N__8914),
            .I(N__8911));
    LocalMux I__1706 (
            .O(N__8911),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_7 ));
    InMux I__1705 (
            .O(N__8908),
            .I(N__8905));
    LocalMux I__1704 (
            .O(N__8905),
            .I(\DUT.uart_inst0.tx_out_6_iv_0_a3_0_1 ));
    InMux I__1703 (
            .O(N__8902),
            .I(N__8899));
    LocalMux I__1702 (
            .O(N__8899),
            .I(\DUT.uart_inst0.N_101 ));
    InMux I__1701 (
            .O(N__8896),
            .I(N__8893));
    LocalMux I__1700 (
            .O(N__8893),
            .I(\DUT.rFifoDatarx_5 ));
    InMux I__1699 (
            .O(N__8890),
            .I(N__8887));
    LocalMux I__1698 (
            .O(N__8887),
            .I(\DUT.rFifoDatarx_0_6 ));
    CascadeMux I__1697 (
            .O(N__8884),
            .I(N__8881));
    InMux I__1696 (
            .O(N__8881),
            .I(N__8878));
    LocalMux I__1695 (
            .O(N__8878),
            .I(\DUT.uart_inst0.tx_dataZ0Z_6 ));
    InMux I__1694 (
            .O(N__8875),
            .I(N__8872));
    LocalMux I__1693 (
            .O(N__8872),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_2 ));
    CascadeMux I__1692 (
            .O(N__8869),
            .I(N__8866));
    InMux I__1691 (
            .O(N__8866),
            .I(N__8863));
    LocalMux I__1690 (
            .O(N__8863),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_2 ));
    InMux I__1689 (
            .O(N__8860),
            .I(N__8857));
    LocalMux I__1688 (
            .O(N__8857),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_1 ));
    CascadeMux I__1687 (
            .O(N__8854),
            .I(N__8851));
    InMux I__1686 (
            .O(N__8851),
            .I(N__8848));
    LocalMux I__1685 (
            .O(N__8848),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_1 ));
    InMux I__1684 (
            .O(N__8845),
            .I(N__8842));
    LocalMux I__1683 (
            .O(N__8842),
            .I(N__8839));
    Odrv4 I__1682 (
            .O(N__8839),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1 ));
    InMux I__1681 (
            .O(N__8836),
            .I(N__8833));
    LocalMux I__1680 (
            .O(N__8833),
            .I(N__8830));
    Span4Mux_h I__1679 (
            .O(N__8830),
            .I(N__8827));
    Odrv4 I__1678 (
            .O(N__8827),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_2 ));
    InMux I__1677 (
            .O(N__8824),
            .I(N__8821));
    LocalMux I__1676 (
            .O(N__8821),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2 ));
    InMux I__1675 (
            .O(N__8818),
            .I(N__8815));
    LocalMux I__1674 (
            .O(N__8815),
            .I(N__8812));
    Span4Mux_h I__1673 (
            .O(N__8812),
            .I(N__8809));
    Odrv4 I__1672 (
            .O(N__8809),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_3 ));
    CascadeMux I__1671 (
            .O(N__8806),
            .I(N__8803));
    InMux I__1670 (
            .O(N__8803),
            .I(N__8800));
    LocalMux I__1669 (
            .O(N__8800),
            .I(N__8797));
    Span4Mux_v I__1668 (
            .O(N__8797),
            .I(N__8794));
    Odrv4 I__1667 (
            .O(N__8794),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_3 ));
    InMux I__1666 (
            .O(N__8791),
            .I(N__8788));
    LocalMux I__1665 (
            .O(N__8788),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_3 ));
    CascadeMux I__1664 (
            .O(N__8785),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ));
    InMux I__1663 (
            .O(N__8782),
            .I(N__8779));
    LocalMux I__1662 (
            .O(N__8779),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_3 ));
    InMux I__1661 (
            .O(N__8776),
            .I(N__8773));
    LocalMux I__1660 (
            .O(N__8773),
            .I(N__8770));
    Span4Mux_h I__1659 (
            .O(N__8770),
            .I(N__8767));
    Odrv4 I__1658 (
            .O(N__8767),
            .I(\DUT.rFifoDatarx_0_0 ));
    InMux I__1657 (
            .O(N__8764),
            .I(N__8761));
    LocalMux I__1656 (
            .O(N__8761),
            .I(N__8758));
    Span4Mux_s2_v I__1655 (
            .O(N__8758),
            .I(N__8755));
    Span4Mux_v I__1654 (
            .O(N__8755),
            .I(N__8752));
    Odrv4 I__1653 (
            .O(N__8752),
            .I(\DUT.uart_inst0.tx_out_6_iv_0_1 ));
    InMux I__1652 (
            .O(N__8749),
            .I(N__8746));
    LocalMux I__1651 (
            .O(N__8746),
            .I(\DUT.rFifoDatarx_1 ));
    CascadeMux I__1650 (
            .O(N__8743),
            .I(N__8740));
    InMux I__1649 (
            .O(N__8740),
            .I(N__8737));
    LocalMux I__1648 (
            .O(N__8737),
            .I(\DUT.uart_inst0.tx_dataZ0Z_1 ));
    InMux I__1647 (
            .O(N__8734),
            .I(N__8731));
    LocalMux I__1646 (
            .O(N__8731),
            .I(\DUT.rFifoDatarx_2 ));
    InMux I__1645 (
            .O(N__8728),
            .I(N__8725));
    LocalMux I__1644 (
            .O(N__8725),
            .I(N__8722));
    Odrv4 I__1643 (
            .O(N__8722),
            .I(\DUT.uart_inst0.N_31_0 ));
    InMux I__1642 (
            .O(N__8719),
            .I(N__8716));
    LocalMux I__1641 (
            .O(N__8716),
            .I(\DUT.uart_inst0.N_203 ));
    InMux I__1640 (
            .O(N__8713),
            .I(N__8710));
    LocalMux I__1639 (
            .O(N__8710),
            .I(\DUT.uart_inst0.recv_state_ns_0_i_0_0_a3_0_0_3 ));
    InMux I__1638 (
            .O(N__8707),
            .I(N__8703));
    InMux I__1637 (
            .O(N__8706),
            .I(N__8698));
    LocalMux I__1636 (
            .O(N__8703),
            .I(N__8695));
    InMux I__1635 (
            .O(N__8702),
            .I(N__8692));
    InMux I__1634 (
            .O(N__8701),
            .I(N__8689));
    LocalMux I__1633 (
            .O(N__8698),
            .I(N__8686));
    Span4Mux_h I__1632 (
            .O(N__8695),
            .I(N__8683));
    LocalMux I__1631 (
            .O(N__8692),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_2 ));
    LocalMux I__1630 (
            .O(N__8689),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_2 ));
    Odrv4 I__1629 (
            .O(N__8686),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_2 ));
    Odrv4 I__1628 (
            .O(N__8683),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_2 ));
    InMux I__1627 (
            .O(N__8674),
            .I(N__8669));
    InMux I__1626 (
            .O(N__8673),
            .I(N__8666));
    CascadeMux I__1625 (
            .O(N__8672),
            .I(N__8663));
    LocalMux I__1624 (
            .O(N__8669),
            .I(N__8655));
    LocalMux I__1623 (
            .O(N__8666),
            .I(N__8655));
    InMux I__1622 (
            .O(N__8663),
            .I(N__8652));
    InMux I__1621 (
            .O(N__8662),
            .I(N__8645));
    InMux I__1620 (
            .O(N__8661),
            .I(N__8645));
    InMux I__1619 (
            .O(N__8660),
            .I(N__8645));
    Span4Mux_v I__1618 (
            .O(N__8655),
            .I(N__8642));
    LocalMux I__1617 (
            .O(N__8652),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_1 ));
    LocalMux I__1616 (
            .O(N__8645),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_1 ));
    Odrv4 I__1615 (
            .O(N__8642),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_1 ));
    CascadeMux I__1614 (
            .O(N__8635),
            .I(N__8632));
    InMux I__1613 (
            .O(N__8632),
            .I(N__8628));
    InMux I__1612 (
            .O(N__8631),
            .I(N__8625));
    LocalMux I__1611 (
            .O(N__8628),
            .I(N__8622));
    LocalMux I__1610 (
            .O(N__8625),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_3 ));
    Odrv4 I__1609 (
            .O(N__8622),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_3 ));
    CascadeMux I__1608 (
            .O(N__8617),
            .I(N__8614));
    InMux I__1607 (
            .O(N__8614),
            .I(N__8610));
    CascadeMux I__1606 (
            .O(N__8613),
            .I(N__8606));
    LocalMux I__1605 (
            .O(N__8610),
            .I(N__8601));
    InMux I__1604 (
            .O(N__8609),
            .I(N__8598));
    InMux I__1603 (
            .O(N__8606),
            .I(N__8591));
    InMux I__1602 (
            .O(N__8605),
            .I(N__8591));
    InMux I__1601 (
            .O(N__8604),
            .I(N__8591));
    Span4Mux_s3_v I__1600 (
            .O(N__8601),
            .I(N__8586));
    LocalMux I__1599 (
            .O(N__8598),
            .I(N__8586));
    LocalMux I__1598 (
            .O(N__8591),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_0 ));
    Odrv4 I__1597 (
            .O(N__8586),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_0 ));
    InMux I__1596 (
            .O(N__8581),
            .I(N__8578));
    LocalMux I__1595 (
            .O(N__8578),
            .I(\DUT.uart_inst0.N_215_4 ));
    CascadeMux I__1594 (
            .O(N__8575),
            .I(\DUT.uart_inst0.N_215_4_cascade_ ));
    CascadeMux I__1593 (
            .O(N__8572),
            .I(\DUT.uart_inst0.recv_state_srsts_1_2_cascade_ ));
    InMux I__1592 (
            .O(N__8569),
            .I(N__8565));
    InMux I__1591 (
            .O(N__8568),
            .I(N__8562));
    LocalMux I__1590 (
            .O(N__8565),
            .I(\DUT.uart_inst0.N_193 ));
    LocalMux I__1589 (
            .O(N__8562),
            .I(\DUT.uart_inst0.N_193 ));
    InMux I__1588 (
            .O(N__8557),
            .I(N__8548));
    InMux I__1587 (
            .O(N__8556),
            .I(N__8543));
    InMux I__1586 (
            .O(N__8555),
            .I(N__8543));
    InMux I__1585 (
            .O(N__8554),
            .I(N__8540));
    InMux I__1584 (
            .O(N__8553),
            .I(N__8533));
    InMux I__1583 (
            .O(N__8552),
            .I(N__8533));
    InMux I__1582 (
            .O(N__8551),
            .I(N__8533));
    LocalMux I__1581 (
            .O(N__8548),
            .I(\DUT.uart_inst0.recv_stateZ0Z_2 ));
    LocalMux I__1580 (
            .O(N__8543),
            .I(\DUT.uart_inst0.recv_stateZ0Z_2 ));
    LocalMux I__1579 (
            .O(N__8540),
            .I(\DUT.uart_inst0.recv_stateZ0Z_2 ));
    LocalMux I__1578 (
            .O(N__8533),
            .I(\DUT.uart_inst0.recv_stateZ0Z_2 ));
    InMux I__1577 (
            .O(N__8524),
            .I(N__8521));
    LocalMux I__1576 (
            .O(N__8521),
            .I(N__8518));
    Odrv4 I__1575 (
            .O(N__8518),
            .I(\DUT.uart_inst0.g0_0 ));
    InMux I__1574 (
            .O(N__8515),
            .I(N__8511));
    InMux I__1573 (
            .O(N__8514),
            .I(N__8507));
    LocalMux I__1572 (
            .O(N__8511),
            .I(N__8503));
    InMux I__1571 (
            .O(N__8510),
            .I(N__8500));
    LocalMux I__1570 (
            .O(N__8507),
            .I(N__8497));
    InMux I__1569 (
            .O(N__8506),
            .I(N__8494));
    Span4Mux_v I__1568 (
            .O(N__8503),
            .I(N__8491));
    LocalMux I__1567 (
            .O(N__8500),
            .I(N__8488));
    Span4Mux_h I__1566 (
            .O(N__8497),
            .I(N__8483));
    LocalMux I__1565 (
            .O(N__8494),
            .I(N__8483));
    Span4Mux_v I__1564 (
            .O(N__8491),
            .I(N__8479));
    Span4Mux_v I__1563 (
            .O(N__8488),
            .I(N__8476));
    Span4Mux_v I__1562 (
            .O(N__8483),
            .I(N__8473));
    InMux I__1561 (
            .O(N__8482),
            .I(N__8470));
    Odrv4 I__1560 (
            .O(N__8479),
            .I(\DUT.wRxByte_3 ));
    Odrv4 I__1559 (
            .O(N__8476),
            .I(\DUT.wRxByte_3 ));
    Odrv4 I__1558 (
            .O(N__8473),
            .I(\DUT.wRxByte_3 ));
    LocalMux I__1557 (
            .O(N__8470),
            .I(\DUT.wRxByte_3 ));
    InMux I__1556 (
            .O(N__8461),
            .I(N__8456));
    InMux I__1555 (
            .O(N__8460),
            .I(N__8453));
    InMux I__1554 (
            .O(N__8459),
            .I(N__8450));
    LocalMux I__1553 (
            .O(N__8456),
            .I(N__8446));
    LocalMux I__1552 (
            .O(N__8453),
            .I(N__8441));
    LocalMux I__1551 (
            .O(N__8450),
            .I(N__8441));
    InMux I__1550 (
            .O(N__8449),
            .I(N__8438));
    Span4Mux_h I__1549 (
            .O(N__8446),
            .I(N__8431));
    Span4Mux_v I__1548 (
            .O(N__8441),
            .I(N__8431));
    LocalMux I__1547 (
            .O(N__8438),
            .I(N__8431));
    Span4Mux_v I__1546 (
            .O(N__8431),
            .I(N__8427));
    InMux I__1545 (
            .O(N__8430),
            .I(N__8424));
    Odrv4 I__1544 (
            .O(N__8427),
            .I(\DUT.wRxByte_2 ));
    LocalMux I__1543 (
            .O(N__8424),
            .I(\DUT.wRxByte_2 ));
    CEMux I__1542 (
            .O(N__8419),
            .I(N__8415));
    CEMux I__1541 (
            .O(N__8418),
            .I(N__8412));
    LocalMux I__1540 (
            .O(N__8415),
            .I(N__8409));
    LocalMux I__1539 (
            .O(N__8412),
            .I(N__8406));
    Span4Mux_h I__1538 (
            .O(N__8409),
            .I(N__8403));
    Span4Mux_h I__1537 (
            .O(N__8406),
            .I(N__8400));
    Odrv4 I__1536 (
            .O(N__8403),
            .I(\DUT.uart_inst0.rx_bits_remaining_2_sqmuxa ));
    Odrv4 I__1535 (
            .O(N__8400),
            .I(\DUT.uart_inst0.rx_bits_remaining_2_sqmuxa ));
    InMux I__1534 (
            .O(N__8395),
            .I(N__8392));
    LocalMux I__1533 (
            .O(N__8392),
            .I(\DUT.uart_inst0.g0_0_3 ));
    InMux I__1532 (
            .O(N__8389),
            .I(N__8386));
    LocalMux I__1531 (
            .O(N__8386),
            .I(\DUT.uart_inst0.g1 ));
    CascadeMux I__1530 (
            .O(N__8383),
            .I(N__8380));
    InMux I__1529 (
            .O(N__8380),
            .I(N__8377));
    LocalMux I__1528 (
            .O(N__8377),
            .I(\DUT.uart_inst0.g0_0_0 ));
    InMux I__1527 (
            .O(N__8374),
            .I(N__8371));
    LocalMux I__1526 (
            .O(N__8371),
            .I(N__8368));
    Span4Mux_v I__1525 (
            .O(N__8368),
            .I(N__8365));
    Odrv4 I__1524 (
            .O(N__8365),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_2 ));
    InMux I__1523 (
            .O(N__8362),
            .I(N__8358));
    InMux I__1522 (
            .O(N__8361),
            .I(N__8355));
    LocalMux I__1521 (
            .O(N__8358),
            .I(\DUT.uart_inst0.rx_clk_divider_1_17 ));
    LocalMux I__1520 (
            .O(N__8355),
            .I(\DUT.uart_inst0.rx_clk_divider_1_17 ));
    InMux I__1519 (
            .O(N__8350),
            .I(N__8347));
    LocalMux I__1518 (
            .O(N__8347),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_17 ));
    InMux I__1517 (
            .O(N__8344),
            .I(N__8340));
    InMux I__1516 (
            .O(N__8343),
            .I(N__8337));
    LocalMux I__1515 (
            .O(N__8340),
            .I(\DUT.uart_inst0.rx_clk_divider_1_10 ));
    LocalMux I__1514 (
            .O(N__8337),
            .I(\DUT.uart_inst0.rx_clk_divider_1_10 ));
    InMux I__1513 (
            .O(N__8332),
            .I(N__8329));
    LocalMux I__1512 (
            .O(N__8329),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_10 ));
    InMux I__1511 (
            .O(N__8326),
            .I(N__8322));
    InMux I__1510 (
            .O(N__8325),
            .I(N__8319));
    LocalMux I__1509 (
            .O(N__8322),
            .I(\DUT.uart_inst0.rx_clk_divider_1_13 ));
    LocalMux I__1508 (
            .O(N__8319),
            .I(\DUT.uart_inst0.rx_clk_divider_1_13 ));
    InMux I__1507 (
            .O(N__8314),
            .I(N__8311));
    LocalMux I__1506 (
            .O(N__8311),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_13 ));
    InMux I__1505 (
            .O(N__8308),
            .I(N__8305));
    LocalMux I__1504 (
            .O(N__8305),
            .I(N__8302));
    Span4Mux_h I__1503 (
            .O(N__8302),
            .I(N__8299));
    Odrv4 I__1502 (
            .O(N__8299),
            .I(\DUT.uart_inst0.N_199_0 ));
    IoInMux I__1501 (
            .O(N__8296),
            .I(N__8293));
    LocalMux I__1500 (
            .O(N__8293),
            .I(N__8290));
    IoSpan4Mux I__1499 (
            .O(N__8290),
            .I(N__8287));
    Odrv4 I__1498 (
            .O(N__8287),
            .I(N_1239_i));
    CascadeMux I__1497 (
            .O(N__8284),
            .I(N__8281));
    InMux I__1496 (
            .O(N__8281),
            .I(N__8276));
    InMux I__1495 (
            .O(N__8280),
            .I(N__8273));
    InMux I__1494 (
            .O(N__8279),
            .I(N__8270));
    LocalMux I__1493 (
            .O(N__8276),
            .I(N__8265));
    LocalMux I__1492 (
            .O(N__8273),
            .I(N__8265));
    LocalMux I__1491 (
            .O(N__8270),
            .I(\DUT.uart_inst0.recv_stateZ0Z_0 ));
    Odrv12 I__1490 (
            .O(N__8265),
            .I(\DUT.uart_inst0.recv_stateZ0Z_0 ));
    CascadeMux I__1489 (
            .O(N__8260),
            .I(N__8257));
    InMux I__1488 (
            .O(N__8257),
            .I(N__8253));
    InMux I__1487 (
            .O(N__8256),
            .I(N__8250));
    LocalMux I__1486 (
            .O(N__8253),
            .I(N__8247));
    LocalMux I__1485 (
            .O(N__8250),
            .I(N__8244));
    Span4Mux_h I__1484 (
            .O(N__8247),
            .I(N__8241));
    Odrv4 I__1483 (
            .O(N__8244),
            .I(\DUT.uart_inst0.rx_clk_divider_5_i_a2_12_1_5 ));
    Odrv4 I__1482 (
            .O(N__8241),
            .I(\DUT.uart_inst0.rx_clk_divider_5_i_a2_12_1_5 ));
    InMux I__1481 (
            .O(N__8236),
            .I(N__8231));
    InMux I__1480 (
            .O(N__8235),
            .I(N__8226));
    InMux I__1479 (
            .O(N__8234),
            .I(N__8226));
    LocalMux I__1478 (
            .O(N__8231),
            .I(\DUT.uart_inst0.rx_clk_divider_1_16 ));
    LocalMux I__1477 (
            .O(N__8226),
            .I(\DUT.uart_inst0.rx_clk_divider_1_16 ));
    CascadeMux I__1476 (
            .O(N__8221),
            .I(N__8217));
    InMux I__1475 (
            .O(N__8220),
            .I(N__8214));
    InMux I__1474 (
            .O(N__8217),
            .I(N__8211));
    LocalMux I__1473 (
            .O(N__8214),
            .I(N__8208));
    LocalMux I__1472 (
            .O(N__8211),
            .I(N__8205));
    Span4Mux_h I__1471 (
            .O(N__8208),
            .I(N__8202));
    Odrv4 I__1470 (
            .O(N__8205),
            .I(\DUT.uart_inst0.rx_clk_divider_5_i_a2_12_4_5 ));
    Odrv4 I__1469 (
            .O(N__8202),
            .I(\DUT.uart_inst0.rx_clk_divider_5_i_a2_12_4_5 ));
    InMux I__1468 (
            .O(N__8197),
            .I(N__8192));
    InMux I__1467 (
            .O(N__8196),
            .I(N__8187));
    InMux I__1466 (
            .O(N__8195),
            .I(N__8187));
    LocalMux I__1465 (
            .O(N__8192),
            .I(\DUT.uart_inst0.rx_clk_divider_1_14 ));
    LocalMux I__1464 (
            .O(N__8187),
            .I(\DUT.uart_inst0.rx_clk_divider_1_14 ));
    InMux I__1463 (
            .O(N__8182),
            .I(N__8176));
    InMux I__1462 (
            .O(N__8181),
            .I(N__8176));
    LocalMux I__1461 (
            .O(N__8176),
            .I(N__8173));
    Span4Mux_s2_v I__1460 (
            .O(N__8173),
            .I(N__8170));
    Odrv4 I__1459 (
            .O(N__8170),
            .I(\DUT.uart_inst0.rx_clk_divider_5_i_a2_12_5 ));
    CascadeMux I__1458 (
            .O(N__8167),
            .I(N__8163));
    CascadeMux I__1457 (
            .O(N__8166),
            .I(N__8160));
    InMux I__1456 (
            .O(N__8163),
            .I(N__8155));
    InMux I__1455 (
            .O(N__8160),
            .I(N__8155));
    LocalMux I__1454 (
            .O(N__8155),
            .I(\DUT.uart_inst0.rx_clk_divider_1_9 ));
    InMux I__1453 (
            .O(N__8152),
            .I(N__8149));
    LocalMux I__1452 (
            .O(N__8149),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_9 ));
    InMux I__1451 (
            .O(N__8146),
            .I(N__8140));
    InMux I__1450 (
            .O(N__8145),
            .I(N__8140));
    LocalMux I__1449 (
            .O(N__8140),
            .I(\DUT.uart_inst0.rx_clk_divider_1_11 ));
    InMux I__1448 (
            .O(N__8137),
            .I(N__8134));
    LocalMux I__1447 (
            .O(N__8134),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_11 ));
    InMux I__1446 (
            .O(N__8131),
            .I(N__8125));
    InMux I__1445 (
            .O(N__8130),
            .I(N__8125));
    LocalMux I__1444 (
            .O(N__8125),
            .I(\DUT.uart_inst0.rx_clk_divider_1_12 ));
    InMux I__1443 (
            .O(N__8122),
            .I(N__8119));
    LocalMux I__1442 (
            .O(N__8119),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_12 ));
    CascadeMux I__1441 (
            .O(N__8116),
            .I(N__8111));
    CascadeMux I__1440 (
            .O(N__8115),
            .I(N__8108));
    InMux I__1439 (
            .O(N__8114),
            .I(N__8103));
    InMux I__1438 (
            .O(N__8111),
            .I(N__8103));
    InMux I__1437 (
            .O(N__8108),
            .I(N__8100));
    LocalMux I__1436 (
            .O(N__8103),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_1 ));
    LocalMux I__1435 (
            .O(N__8100),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_1 ));
    InMux I__1434 (
            .O(N__8095),
            .I(N__8092));
    LocalMux I__1433 (
            .O(N__8092),
            .I(N__8088));
    InMux I__1432 (
            .O(N__8091),
            .I(N__8085));
    Odrv4 I__1431 (
            .O(N__8088),
            .I(\DUT.uart_inst0.rx_clk_divider_1_7 ));
    LocalMux I__1430 (
            .O(N__8085),
            .I(\DUT.uart_inst0.rx_clk_divider_1_7 ));
    InMux I__1429 (
            .O(N__8080),
            .I(N__8074));
    InMux I__1428 (
            .O(N__8079),
            .I(N__8074));
    LocalMux I__1427 (
            .O(N__8074),
            .I(\DUT.uart_inst0.rx_clk_divider_1_1 ));
    CascadeMux I__1426 (
            .O(N__8071),
            .I(N__8068));
    InMux I__1425 (
            .O(N__8068),
            .I(N__8065));
    LocalMux I__1424 (
            .O(N__8065),
            .I(\DUT.uart_inst0.rx_clk_dividerZ1Z_1 ));
    InMux I__1423 (
            .O(N__8062),
            .I(N__8059));
    LocalMux I__1422 (
            .O(N__8059),
            .I(N__8056));
    Span4Mux_h I__1421 (
            .O(N__8056),
            .I(N__8053));
    Odrv4 I__1420 (
            .O(N__8053),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_5 ));
    InMux I__1419 (
            .O(N__8050),
            .I(N__8047));
    LocalMux I__1418 (
            .O(N__8047),
            .I(N__8043));
    InMux I__1417 (
            .O(N__8046),
            .I(N__8040));
    Span4Mux_s2_v I__1416 (
            .O(N__8043),
            .I(N__8036));
    LocalMux I__1415 (
            .O(N__8040),
            .I(N__8033));
    CascadeMux I__1414 (
            .O(N__8039),
            .I(N__8023));
    Span4Mux_h I__1413 (
            .O(N__8036),
            .I(N__8017));
    Span4Mux_s2_v I__1412 (
            .O(N__8033),
            .I(N__8017));
    InMux I__1411 (
            .O(N__8032),
            .I(N__8012));
    InMux I__1410 (
            .O(N__8031),
            .I(N__8012));
    InMux I__1409 (
            .O(N__8030),
            .I(N__8005));
    InMux I__1408 (
            .O(N__8029),
            .I(N__8005));
    InMux I__1407 (
            .O(N__8028),
            .I(N__8005));
    InMux I__1406 (
            .O(N__8027),
            .I(N__8002));
    InMux I__1405 (
            .O(N__8026),
            .I(N__7995));
    InMux I__1404 (
            .O(N__8023),
            .I(N__7995));
    InMux I__1403 (
            .O(N__8022),
            .I(N__7995));
    Odrv4 I__1402 (
            .O(N__8017),
            .I(\DUT.uart_inst0.rx_countdown_3_1 ));
    LocalMux I__1401 (
            .O(N__8012),
            .I(\DUT.uart_inst0.rx_countdown_3_1 ));
    LocalMux I__1400 (
            .O(N__8005),
            .I(\DUT.uart_inst0.rx_countdown_3_1 ));
    LocalMux I__1399 (
            .O(N__8002),
            .I(\DUT.uart_inst0.rx_countdown_3_1 ));
    LocalMux I__1398 (
            .O(N__7995),
            .I(\DUT.uart_inst0.rx_countdown_3_1 ));
    InMux I__1397 (
            .O(N__7984),
            .I(N__7981));
    LocalMux I__1396 (
            .O(N__7981),
            .I(N__7978));
    Span4Mux_h I__1395 (
            .O(N__7978),
            .I(N__7975));
    Odrv4 I__1394 (
            .O(N__7975),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_1 ));
    InMux I__1393 (
            .O(N__7972),
            .I(N__7969));
    LocalMux I__1392 (
            .O(N__7969),
            .I(N__7965));
    InMux I__1391 (
            .O(N__7968),
            .I(N__7962));
    Odrv4 I__1390 (
            .O(N__7965),
            .I(\DUT.uart_inst0.rx_clk_divider_1_2 ));
    LocalMux I__1389 (
            .O(N__7962),
            .I(\DUT.uart_inst0.rx_clk_divider_1_2 ));
    CascadeMux I__1388 (
            .O(N__7957),
            .I(N__7954));
    InMux I__1387 (
            .O(N__7954),
            .I(N__7951));
    LocalMux I__1386 (
            .O(N__7951),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_2 ));
    CEMux I__1385 (
            .O(N__7948),
            .I(N__7945));
    LocalMux I__1384 (
            .O(N__7945),
            .I(N__7942));
    Span4Mux_h I__1383 (
            .O(N__7942),
            .I(N__7938));
    InMux I__1382 (
            .O(N__7941),
            .I(N__7935));
    Odrv4 I__1381 (
            .O(N__7938),
            .I(\DUT.fifo_tx_inst.rFifoData_awe2 ));
    LocalMux I__1380 (
            .O(N__7935),
            .I(\DUT.fifo_tx_inst.rFifoData_awe2 ));
    InMux I__1379 (
            .O(N__7930),
            .I(N__7926));
    InMux I__1378 (
            .O(N__7929),
            .I(N__7923));
    LocalMux I__1377 (
            .O(N__7926),
            .I(N__7920));
    LocalMux I__1376 (
            .O(N__7923),
            .I(\DUT.fifo_tx_inst.rFifoDataro_2 ));
    Odrv4 I__1375 (
            .O(N__7920),
            .I(\DUT.fifo_tx_inst.rFifoDataro_2 ));
    InMux I__1374 (
            .O(N__7915),
            .I(N__7908));
    InMux I__1373 (
            .O(N__7914),
            .I(N__7908));
    InMux I__1372 (
            .O(N__7913),
            .I(N__7905));
    LocalMux I__1371 (
            .O(N__7908),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4 ));
    LocalMux I__1370 (
            .O(N__7905),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4 ));
    CascadeMux I__1369 (
            .O(N__7900),
            .I(N__7897));
    InMux I__1368 (
            .O(N__7897),
            .I(N__7890));
    InMux I__1367 (
            .O(N__7896),
            .I(N__7890));
    InMux I__1366 (
            .O(N__7895),
            .I(N__7887));
    LocalMux I__1365 (
            .O(N__7890),
            .I(\fifo_inst.ftdi_output_inst.rWrDelayZ0 ));
    LocalMux I__1364 (
            .O(N__7887),
            .I(\fifo_inst.ftdi_output_inst.rWrDelayZ0 ));
    InMux I__1363 (
            .O(N__7882),
            .I(N__7876));
    InMux I__1362 (
            .O(N__7881),
            .I(N__7876));
    LocalMux I__1361 (
            .O(N__7876),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_3 ));
    IoInMux I__1360 (
            .O(N__7873),
            .I(N__7870));
    LocalMux I__1359 (
            .O(N__7870),
            .I(N__7866));
    IoInMux I__1358 (
            .O(N__7869),
            .I(N__7863));
    Span4Mux_s3_v I__1357 (
            .O(N__7866),
            .I(N__7860));
    LocalMux I__1356 (
            .O(N__7863),
            .I(N__7857));
    Span4Mux_v I__1355 (
            .O(N__7860),
            .I(N__7854));
    Span12Mux_s7_v I__1354 (
            .O(N__7857),
            .I(N__7851));
    Span4Mux_h I__1353 (
            .O(N__7854),
            .I(N__7848));
    Span12Mux_v I__1352 (
            .O(N__7851),
            .I(N__7844));
    Span4Mux_h I__1351 (
            .O(N__7848),
            .I(N__7841));
    InMux I__1350 (
            .O(N__7847),
            .I(N__7838));
    Odrv12 I__1349 (
            .O(N__7844),
            .I(P1A4_c));
    Odrv4 I__1348 (
            .O(N__7841),
            .I(P1A4_c));
    LocalMux I__1347 (
            .O(N__7838),
            .I(P1A4_c));
    IoInMux I__1346 (
            .O(N__7831),
            .I(N__7826));
    IoInMux I__1345 (
            .O(N__7830),
            .I(N__7823));
    IoInMux I__1344 (
            .O(N__7829),
            .I(N__7820));
    LocalMux I__1343 (
            .O(N__7826),
            .I(N__7814));
    LocalMux I__1342 (
            .O(N__7823),
            .I(N__7814));
    LocalMux I__1341 (
            .O(N__7820),
            .I(N__7811));
    IoInMux I__1340 (
            .O(N__7819),
            .I(N__7808));
    Span4Mux_s3_v I__1339 (
            .O(N__7814),
            .I(N__7805));
    IoSpan4Mux I__1338 (
            .O(N__7811),
            .I(N__7802));
    LocalMux I__1337 (
            .O(N__7808),
            .I(N__7799));
    Span4Mux_h I__1336 (
            .O(N__7805),
            .I(N__7796));
    Span4Mux_s2_v I__1335 (
            .O(N__7802),
            .I(N__7791));
    Span4Mux_s2_v I__1334 (
            .O(N__7799),
            .I(N__7791));
    Sp12to4 I__1333 (
            .O(N__7796),
            .I(N__7788));
    Span4Mux_v I__1332 (
            .O(N__7791),
            .I(N__7785));
    Span12Mux_v I__1331 (
            .O(N__7788),
            .I(N__7781));
    Span4Mux_v I__1330 (
            .O(N__7785),
            .I(N__7778));
    InMux I__1329 (
            .O(N__7784),
            .I(N__7775));
    Odrv12 I__1328 (
            .O(N__7781),
            .I(rTxBusReady));
    Odrv4 I__1327 (
            .O(N__7778),
            .I(rTxBusReady));
    LocalMux I__1326 (
            .O(N__7775),
            .I(rTxBusReady));
    InMux I__1325 (
            .O(N__7768),
            .I(N__7762));
    InMux I__1324 (
            .O(N__7767),
            .I(N__7762));
    LocalMux I__1323 (
            .O(N__7762),
            .I(\DUT.uart_inst0.rx_clk_divider_1_8 ));
    InMux I__1322 (
            .O(N__7759),
            .I(N__7756));
    LocalMux I__1321 (
            .O(N__7756),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_8 ));
    InMux I__1320 (
            .O(N__7753),
            .I(N__7750));
    LocalMux I__1319 (
            .O(N__7750),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_6 ));
    CascadeMux I__1318 (
            .O(N__7747),
            .I(N__7744));
    InMux I__1317 (
            .O(N__7744),
            .I(N__7741));
    LocalMux I__1316 (
            .O(N__7741),
            .I(N__7738));
    Span4Mux_h I__1315 (
            .O(N__7738),
            .I(N__7735));
    Span4Mux_h I__1314 (
            .O(N__7735),
            .I(N__7732));
    Odrv4 I__1313 (
            .O(N__7732),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_6 ));
    InMux I__1312 (
            .O(N__7729),
            .I(N__7725));
    InMux I__1311 (
            .O(N__7728),
            .I(N__7722));
    LocalMux I__1310 (
            .O(N__7725),
            .I(\DUT.fifo_tx_inst.rFifoDataro_3 ));
    LocalMux I__1309 (
            .O(N__7722),
            .I(\DUT.fifo_tx_inst.rFifoDataro_3 ));
    InMux I__1308 (
            .O(N__7717),
            .I(N__7713));
    InMux I__1307 (
            .O(N__7716),
            .I(N__7710));
    LocalMux I__1306 (
            .O(N__7713),
            .I(\DUT.fifo_tx_inst.rFifoDataro_0 ));
    LocalMux I__1305 (
            .O(N__7710),
            .I(\DUT.fifo_tx_inst.rFifoDataro_0 ));
    CascadeMux I__1304 (
            .O(N__7705),
            .I(N__7701));
    InMux I__1303 (
            .O(N__7704),
            .I(N__7698));
    InMux I__1302 (
            .O(N__7701),
            .I(N__7695));
    LocalMux I__1301 (
            .O(N__7698),
            .I(\DUT.fifo_tx_inst.rFifoDataro_1 ));
    LocalMux I__1300 (
            .O(N__7695),
            .I(\DUT.fifo_tx_inst.rFifoDataro_1 ));
    InMux I__1299 (
            .O(N__7690),
            .I(N__7687));
    LocalMux I__1298 (
            .O(N__7687),
            .I(\DUT.rFifoDataror_0_0_0 ));
    CascadeMux I__1297 (
            .O(N__7684),
            .I(\DUT.rFifoDataror_1_0_cascade_ ));
    InMux I__1296 (
            .O(N__7681),
            .I(N__7678));
    LocalMux I__1295 (
            .O(N__7678),
            .I(N__7675));
    Odrv4 I__1294 (
            .O(N__7675),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_6 ));
    CascadeMux I__1293 (
            .O(N__7672),
            .I(N__7669));
    InMux I__1292 (
            .O(N__7669),
            .I(N__7666));
    LocalMux I__1291 (
            .O(N__7666),
            .I(N__7663));
    Odrv12 I__1290 (
            .O(N__7663),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_6 ));
    InMux I__1289 (
            .O(N__7660),
            .I(N__7657));
    LocalMux I__1288 (
            .O(N__7657),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6 ));
    CascadeMux I__1287 (
            .O(N__7654),
            .I(N__7649));
    CascadeMux I__1286 (
            .O(N__7653),
            .I(N__7643));
    InMux I__1285 (
            .O(N__7652),
            .I(N__7640));
    InMux I__1284 (
            .O(N__7649),
            .I(N__7631));
    InMux I__1283 (
            .O(N__7648),
            .I(N__7631));
    InMux I__1282 (
            .O(N__7647),
            .I(N__7631));
    InMux I__1281 (
            .O(N__7646),
            .I(N__7631));
    InMux I__1280 (
            .O(N__7643),
            .I(N__7628));
    LocalMux I__1279 (
            .O(N__7640),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_0 ));
    LocalMux I__1278 (
            .O(N__7631),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_0 ));
    LocalMux I__1277 (
            .O(N__7628),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_0 ));
    CascadeMux I__1276 (
            .O(N__7621),
            .I(\DUT.fifo_tx_inst.N_79_cascade_ ));
    CascadeMux I__1275 (
            .O(N__7618),
            .I(N__7613));
    InMux I__1274 (
            .O(N__7617),
            .I(N__7608));
    InMux I__1273 (
            .O(N__7616),
            .I(N__7605));
    InMux I__1272 (
            .O(N__7613),
            .I(N__7598));
    InMux I__1271 (
            .O(N__7612),
            .I(N__7598));
    InMux I__1270 (
            .O(N__7611),
            .I(N__7598));
    LocalMux I__1269 (
            .O(N__7608),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_1 ));
    LocalMux I__1268 (
            .O(N__7605),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_1 ));
    LocalMux I__1267 (
            .O(N__7598),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_1 ));
    InMux I__1266 (
            .O(N__7591),
            .I(N__7587));
    InMux I__1265 (
            .O(N__7590),
            .I(N__7584));
    LocalMux I__1264 (
            .O(N__7587),
            .I(N__7579));
    LocalMux I__1263 (
            .O(N__7584),
            .I(N__7576));
    InMux I__1262 (
            .O(N__7583),
            .I(N__7573));
    InMux I__1261 (
            .O(N__7582),
            .I(N__7570));
    Span4Mux_v I__1260 (
            .O(N__7579),
            .I(N__7563));
    Span4Mux_h I__1259 (
            .O(N__7576),
            .I(N__7563));
    LocalMux I__1258 (
            .O(N__7573),
            .I(N__7563));
    LocalMux I__1257 (
            .O(N__7570),
            .I(N__7560));
    Odrv4 I__1256 (
            .O(N__7563),
            .I(rTxByteZ0Z_6));
    Odrv4 I__1255 (
            .O(N__7560),
            .I(rTxByteZ0Z_6));
    InMux I__1254 (
            .O(N__7555),
            .I(N__7552));
    LocalMux I__1253 (
            .O(N__7552),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_4 ));
    InMux I__1252 (
            .O(N__7549),
            .I(N__7546));
    LocalMux I__1251 (
            .O(N__7546),
            .I(N__7543));
    Odrv4 I__1250 (
            .O(N__7543),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_4 ));
    CascadeMux I__1249 (
            .O(N__7540),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_ ));
    InMux I__1248 (
            .O(N__7537),
            .I(N__7534));
    LocalMux I__1247 (
            .O(N__7534),
            .I(N__7531));
    Odrv4 I__1246 (
            .O(N__7531),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_4 ));
    InMux I__1245 (
            .O(N__7528),
            .I(N__7523));
    InMux I__1244 (
            .O(N__7527),
            .I(N__7520));
    InMux I__1243 (
            .O(N__7526),
            .I(N__7517));
    LocalMux I__1242 (
            .O(N__7523),
            .I(N__7513));
    LocalMux I__1241 (
            .O(N__7520),
            .I(N__7510));
    LocalMux I__1240 (
            .O(N__7517),
            .I(N__7507));
    InMux I__1239 (
            .O(N__7516),
            .I(N__7504));
    Span4Mux_v I__1238 (
            .O(N__7513),
            .I(N__7495));
    Span4Mux_v I__1237 (
            .O(N__7510),
            .I(N__7495));
    Span4Mux_h I__1236 (
            .O(N__7507),
            .I(N__7495));
    LocalMux I__1235 (
            .O(N__7504),
            .I(N__7495));
    Odrv4 I__1234 (
            .O(N__7495),
            .I(rTxByteZ0Z_4));
    CascadeMux I__1233 (
            .O(N__7492),
            .I(N__7489));
    InMux I__1232 (
            .O(N__7489),
            .I(N__7486));
    LocalMux I__1231 (
            .O(N__7486),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_4 ));
    InMux I__1230 (
            .O(N__7483),
            .I(N__7480));
    LocalMux I__1229 (
            .O(N__7480),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_5 ));
    InMux I__1228 (
            .O(N__7477),
            .I(N__7474));
    LocalMux I__1227 (
            .O(N__7474),
            .I(N__7471));
    Odrv4 I__1226 (
            .O(N__7471),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_5 ));
    InMux I__1225 (
            .O(N__7468),
            .I(N__7465));
    LocalMux I__1224 (
            .O(N__7465),
            .I(N__7462));
    Odrv4 I__1223 (
            .O(N__7462),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_5 ));
    CascadeMux I__1222 (
            .O(N__7459),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ));
    InMux I__1221 (
            .O(N__7456),
            .I(N__7452));
    InMux I__1220 (
            .O(N__7455),
            .I(N__7449));
    LocalMux I__1219 (
            .O(N__7452),
            .I(N__7445));
    LocalMux I__1218 (
            .O(N__7449),
            .I(N__7442));
    InMux I__1217 (
            .O(N__7448),
            .I(N__7439));
    Span4Mux_v I__1216 (
            .O(N__7445),
            .I(N__7433));
    Span4Mux_v I__1215 (
            .O(N__7442),
            .I(N__7433));
    LocalMux I__1214 (
            .O(N__7439),
            .I(N__7430));
    InMux I__1213 (
            .O(N__7438),
            .I(N__7427));
    Odrv4 I__1212 (
            .O(N__7433),
            .I(rTxByteZ0Z_5));
    Odrv4 I__1211 (
            .O(N__7430),
            .I(rTxByteZ0Z_5));
    LocalMux I__1210 (
            .O(N__7427),
            .I(rTxByteZ0Z_5));
    InMux I__1209 (
            .O(N__7420),
            .I(N__7417));
    LocalMux I__1208 (
            .O(N__7417),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_5 ));
    CEMux I__1207 (
            .O(N__7414),
            .I(N__7409));
    CEMux I__1206 (
            .O(N__7413),
            .I(N__7406));
    CEMux I__1205 (
            .O(N__7412),
            .I(N__7403));
    LocalMux I__1204 (
            .O(N__7409),
            .I(N__7400));
    LocalMux I__1203 (
            .O(N__7406),
            .I(N__7397));
    LocalMux I__1202 (
            .O(N__7403),
            .I(N__7394));
    Span4Mux_h I__1201 (
            .O(N__7400),
            .I(N__7390));
    Span4Mux_v I__1200 (
            .O(N__7397),
            .I(N__7387));
    Span4Mux_h I__1199 (
            .O(N__7394),
            .I(N__7384));
    InMux I__1198 (
            .O(N__7393),
            .I(N__7381));
    Odrv4 I__1197 (
            .O(N__7390),
            .I(\DUT.fifo_tx_inst.rFifoData_awe3 ));
    Odrv4 I__1196 (
            .O(N__7387),
            .I(\DUT.fifo_tx_inst.rFifoData_awe3 ));
    Odrv4 I__1195 (
            .O(N__7384),
            .I(\DUT.fifo_tx_inst.rFifoData_awe3 ));
    LocalMux I__1194 (
            .O(N__7381),
            .I(\DUT.fifo_tx_inst.rFifoData_awe3 ));
    InMux I__1193 (
            .O(N__7372),
            .I(N__7367));
    InMux I__1192 (
            .O(N__7371),
            .I(N__7364));
    InMux I__1191 (
            .O(N__7370),
            .I(N__7361));
    LocalMux I__1190 (
            .O(N__7367),
            .I(N__7357));
    LocalMux I__1189 (
            .O(N__7364),
            .I(N__7354));
    LocalMux I__1188 (
            .O(N__7361),
            .I(N__7351));
    InMux I__1187 (
            .O(N__7360),
            .I(N__7348));
    Span4Mux_v I__1186 (
            .O(N__7357),
            .I(N__7339));
    Span4Mux_v I__1185 (
            .O(N__7354),
            .I(N__7339));
    Span4Mux_h I__1184 (
            .O(N__7351),
            .I(N__7339));
    LocalMux I__1183 (
            .O(N__7348),
            .I(N__7339));
    Odrv4 I__1182 (
            .O(N__7339),
            .I(rTxByteZ0Z_0));
    InMux I__1181 (
            .O(N__7336),
            .I(N__7333));
    LocalMux I__1180 (
            .O(N__7333),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_0 ));
    InMux I__1179 (
            .O(N__7330),
            .I(N__7326));
    InMux I__1178 (
            .O(N__7329),
            .I(N__7323));
    LocalMux I__1177 (
            .O(N__7326),
            .I(N__7319));
    LocalMux I__1176 (
            .O(N__7323),
            .I(N__7316));
    InMux I__1175 (
            .O(N__7322),
            .I(N__7313));
    Span4Mux_h I__1174 (
            .O(N__7319),
            .I(N__7309));
    Span4Mux_v I__1173 (
            .O(N__7316),
            .I(N__7304));
    LocalMux I__1172 (
            .O(N__7313),
            .I(N__7304));
    InMux I__1171 (
            .O(N__7312),
            .I(N__7301));
    Odrv4 I__1170 (
            .O(N__7309),
            .I(rTxByteZ0Z_1));
    Odrv4 I__1169 (
            .O(N__7304),
            .I(rTxByteZ0Z_1));
    LocalMux I__1168 (
            .O(N__7301),
            .I(rTxByteZ0Z_1));
    InMux I__1167 (
            .O(N__7294),
            .I(N__7291));
    LocalMux I__1166 (
            .O(N__7291),
            .I(N__7286));
    InMux I__1165 (
            .O(N__7290),
            .I(N__7283));
    InMux I__1164 (
            .O(N__7289),
            .I(N__7280));
    Span4Mux_h I__1163 (
            .O(N__7286),
            .I(N__7276));
    LocalMux I__1162 (
            .O(N__7283),
            .I(N__7273));
    LocalMux I__1161 (
            .O(N__7280),
            .I(N__7270));
    InMux I__1160 (
            .O(N__7279),
            .I(N__7267));
    Odrv4 I__1159 (
            .O(N__7276),
            .I(rTxByteZ0Z_3));
    Odrv4 I__1158 (
            .O(N__7273),
            .I(rTxByteZ0Z_3));
    Odrv4 I__1157 (
            .O(N__7270),
            .I(rTxByteZ0Z_3));
    LocalMux I__1156 (
            .O(N__7267),
            .I(rTxByteZ0Z_3));
    InMux I__1155 (
            .O(N__7258),
            .I(N__7255));
    LocalMux I__1154 (
            .O(N__7255),
            .I(\DUT.uart_inst0.G_11_i_a4_0_4 ));
    InMux I__1153 (
            .O(N__7252),
            .I(N__7249));
    LocalMux I__1152 (
            .O(N__7249),
            .I(\DUT.uart_inst0.N_4_i_1 ));
    InMux I__1151 (
            .O(N__7246),
            .I(N__7242));
    InMux I__1150 (
            .O(N__7245),
            .I(N__7238));
    LocalMux I__1149 (
            .O(N__7242),
            .I(N__7234));
    InMux I__1148 (
            .O(N__7241),
            .I(N__7231));
    LocalMux I__1147 (
            .O(N__7238),
            .I(N__7228));
    InMux I__1146 (
            .O(N__7237),
            .I(N__7225));
    Span4Mux_v I__1145 (
            .O(N__7234),
            .I(N__7220));
    LocalMux I__1144 (
            .O(N__7231),
            .I(N__7220));
    Span4Mux_h I__1143 (
            .O(N__7228),
            .I(N__7215));
    LocalMux I__1142 (
            .O(N__7225),
            .I(N__7215));
    Span4Mux_h I__1141 (
            .O(N__7220),
            .I(N__7211));
    Span4Mux_v I__1140 (
            .O(N__7215),
            .I(N__7208));
    InMux I__1139 (
            .O(N__7214),
            .I(N__7205));
    Odrv4 I__1138 (
            .O(N__7211),
            .I(\DUT.wRxByte_1 ));
    Odrv4 I__1137 (
            .O(N__7208),
            .I(\DUT.wRxByte_1 ));
    LocalMux I__1136 (
            .O(N__7205),
            .I(\DUT.wRxByte_1 ));
    InMux I__1135 (
            .O(N__7198),
            .I(N__7195));
    LocalMux I__1134 (
            .O(N__7195),
            .I(N__7189));
    InMux I__1133 (
            .O(N__7194),
            .I(N__7186));
    InMux I__1132 (
            .O(N__7193),
            .I(N__7183));
    InMux I__1131 (
            .O(N__7192),
            .I(N__7180));
    Span4Mux_v I__1130 (
            .O(N__7189),
            .I(N__7173));
    LocalMux I__1129 (
            .O(N__7186),
            .I(N__7173));
    LocalMux I__1128 (
            .O(N__7183),
            .I(N__7173));
    LocalMux I__1127 (
            .O(N__7180),
            .I(N__7170));
    Span4Mux_v I__1126 (
            .O(N__7173),
            .I(N__7167));
    Span4Mux_h I__1125 (
            .O(N__7170),
            .I(N__7164));
    Odrv4 I__1124 (
            .O(N__7167),
            .I(\DUT.wRxByte_0 ));
    Odrv4 I__1123 (
            .O(N__7164),
            .I(\DUT.wRxByte_0 ));
    InMux I__1122 (
            .O(N__7159),
            .I(N__7155));
    InMux I__1121 (
            .O(N__7158),
            .I(N__7152));
    LocalMux I__1120 (
            .O(N__7155),
            .I(N__7145));
    LocalMux I__1119 (
            .O(N__7152),
            .I(N__7145));
    InMux I__1118 (
            .O(N__7151),
            .I(N__7142));
    InMux I__1117 (
            .O(N__7150),
            .I(N__7139));
    Span4Mux_v I__1116 (
            .O(N__7145),
            .I(N__7134));
    LocalMux I__1115 (
            .O(N__7142),
            .I(N__7134));
    LocalMux I__1114 (
            .O(N__7139),
            .I(N__7131));
    Span4Mux_v I__1113 (
            .O(N__7134),
            .I(N__7127));
    Span4Mux_v I__1112 (
            .O(N__7131),
            .I(N__7124));
    InMux I__1111 (
            .O(N__7130),
            .I(N__7121));
    Odrv4 I__1110 (
            .O(N__7127),
            .I(\DUT.wRxByte_4 ));
    Odrv4 I__1109 (
            .O(N__7124),
            .I(\DUT.wRxByte_4 ));
    LocalMux I__1108 (
            .O(N__7121),
            .I(\DUT.wRxByte_4 ));
    InMux I__1107 (
            .O(N__7114),
            .I(N__7110));
    InMux I__1106 (
            .O(N__7113),
            .I(N__7107));
    LocalMux I__1105 (
            .O(N__7110),
            .I(N__7100));
    LocalMux I__1104 (
            .O(N__7107),
            .I(N__7100));
    InMux I__1103 (
            .O(N__7106),
            .I(N__7097));
    InMux I__1102 (
            .O(N__7105),
            .I(N__7094));
    Span4Mux_v I__1101 (
            .O(N__7100),
            .I(N__7089));
    LocalMux I__1100 (
            .O(N__7097),
            .I(N__7089));
    LocalMux I__1099 (
            .O(N__7094),
            .I(N__7086));
    Span4Mux_v I__1098 (
            .O(N__7089),
            .I(N__7082));
    Span4Mux_v I__1097 (
            .O(N__7086),
            .I(N__7079));
    InMux I__1096 (
            .O(N__7085),
            .I(N__7076));
    Odrv4 I__1095 (
            .O(N__7082),
            .I(\DUT.wRxByte_5 ));
    Odrv4 I__1094 (
            .O(N__7079),
            .I(\DUT.wRxByte_5 ));
    LocalMux I__1093 (
            .O(N__7076),
            .I(\DUT.wRxByte_5 ));
    InMux I__1092 (
            .O(N__7069),
            .I(N__7065));
    InMux I__1091 (
            .O(N__7068),
            .I(N__7062));
    LocalMux I__1090 (
            .O(N__7065),
            .I(N__7058));
    LocalMux I__1089 (
            .O(N__7062),
            .I(N__7055));
    InMux I__1088 (
            .O(N__7061),
            .I(N__7052));
    Span4Mux_v I__1087 (
            .O(N__7058),
            .I(N__7044));
    Span4Mux_h I__1086 (
            .O(N__7055),
            .I(N__7044));
    LocalMux I__1085 (
            .O(N__7052),
            .I(N__7044));
    InMux I__1084 (
            .O(N__7051),
            .I(N__7041));
    Span4Mux_v I__1083 (
            .O(N__7044),
            .I(N__7037));
    LocalMux I__1082 (
            .O(N__7041),
            .I(N__7034));
    InMux I__1081 (
            .O(N__7040),
            .I(N__7031));
    Odrv4 I__1080 (
            .O(N__7037),
            .I(\DUT.wRxByte_6 ));
    Odrv4 I__1079 (
            .O(N__7034),
            .I(\DUT.wRxByte_6 ));
    LocalMux I__1078 (
            .O(N__7031),
            .I(\DUT.wRxByte_6 ));
    InMux I__1077 (
            .O(N__7024),
            .I(N__7019));
    InMux I__1076 (
            .O(N__7023),
            .I(N__7016));
    InMux I__1075 (
            .O(N__7022),
            .I(N__7013));
    LocalMux I__1074 (
            .O(N__7019),
            .I(N__7007));
    LocalMux I__1073 (
            .O(N__7016),
            .I(N__7007));
    LocalMux I__1072 (
            .O(N__7013),
            .I(N__7004));
    InMux I__1071 (
            .O(N__7012),
            .I(N__7001));
    Span4Mux_v I__1070 (
            .O(N__7007),
            .I(N__6997));
    Span4Mux_h I__1069 (
            .O(N__7004),
            .I(N__6992));
    LocalMux I__1068 (
            .O(N__7001),
            .I(N__6992));
    InMux I__1067 (
            .O(N__7000),
            .I(N__6989));
    Odrv4 I__1066 (
            .O(N__6997),
            .I(\DUT.wRxByte_7 ));
    Odrv4 I__1065 (
            .O(N__6992),
            .I(\DUT.wRxByte_7 ));
    LocalMux I__1064 (
            .O(N__6989),
            .I(\DUT.wRxByte_7 ));
    InMux I__1063 (
            .O(N__6982),
            .I(N__6979));
    LocalMux I__1062 (
            .O(N__6979),
            .I(\DUT.uart_inst0.rx_bits_remaining_2_sqmuxa_0_a2_0_a2_0_a3_1 ));
    CascadeMux I__1061 (
            .O(N__6976),
            .I(\DUT.uart_inst0.rx_countdown_8_i_0_o2_1_2_2_cascade_ ));
    InMux I__1060 (
            .O(N__6973),
            .I(N__6967));
    InMux I__1059 (
            .O(N__6972),
            .I(N__6967));
    LocalMux I__1058 (
            .O(N__6967),
            .I(\DUT.uart_inst0.recv_state_ns_0_i_0_0_o2_0_3 ));
    CascadeMux I__1057 (
            .O(N__6964),
            .I(\DUT.uart_inst0.G_9_1_cascade_ ));
    InMux I__1056 (
            .O(N__6961),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_11 ));
    InMux I__1055 (
            .O(N__6958),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_12 ));
    CascadeMux I__1054 (
            .O(N__6955),
            .I(N__6952));
    InMux I__1053 (
            .O(N__6952),
            .I(N__6949));
    LocalMux I__1052 (
            .O(N__6949),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_14 ));
    InMux I__1051 (
            .O(N__6946),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_13 ));
    InMux I__1050 (
            .O(N__6943),
            .I(N__6940));
    LocalMux I__1049 (
            .O(N__6940),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_15 ));
    InMux I__1048 (
            .O(N__6937),
            .I(N__6933));
    InMux I__1047 (
            .O(N__6936),
            .I(N__6930));
    LocalMux I__1046 (
            .O(N__6933),
            .I(\DUT.uart_inst0.rx_clk_divider_1_15 ));
    LocalMux I__1045 (
            .O(N__6930),
            .I(\DUT.uart_inst0.rx_clk_divider_1_15 ));
    InMux I__1044 (
            .O(N__6925),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_14 ));
    InMux I__1043 (
            .O(N__6922),
            .I(N__6919));
    LocalMux I__1042 (
            .O(N__6919),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_16 ));
    InMux I__1041 (
            .O(N__6916),
            .I(bfn_15_3_0_));
    InMux I__1040 (
            .O(N__6913),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_16 ));
    CascadeMux I__1039 (
            .O(N__6910),
            .I(\DUT.uart_inst0.recv_state_RNO_2Z0Z_4_cascade_ ));
    InMux I__1038 (
            .O(N__6907),
            .I(N__6904));
    LocalMux I__1037 (
            .O(N__6904),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_4 ));
    InMux I__1036 (
            .O(N__6901),
            .I(N__6897));
    InMux I__1035 (
            .O(N__6900),
            .I(N__6894));
    LocalMux I__1034 (
            .O(N__6897),
            .I(\DUT.uart_inst0.rx_clk_divider_1_4 ));
    LocalMux I__1033 (
            .O(N__6894),
            .I(\DUT.uart_inst0.rx_clk_divider_1_4 ));
    InMux I__1032 (
            .O(N__6889),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_3 ));
    CascadeMux I__1031 (
            .O(N__6886),
            .I(N__6883));
    InMux I__1030 (
            .O(N__6883),
            .I(N__6880));
    LocalMux I__1029 (
            .O(N__6880),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_5 ));
    InMux I__1028 (
            .O(N__6877),
            .I(N__6868));
    InMux I__1027 (
            .O(N__6876),
            .I(N__6868));
    InMux I__1026 (
            .O(N__6875),
            .I(N__6868));
    LocalMux I__1025 (
            .O(N__6868),
            .I(\DUT.uart_inst0.rx_clk_divider_1_5 ));
    InMux I__1024 (
            .O(N__6865),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_4 ));
    InMux I__1023 (
            .O(N__6862),
            .I(N__6859));
    LocalMux I__1022 (
            .O(N__6859),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_6 ));
    CascadeMux I__1021 (
            .O(N__6856),
            .I(N__6851));
    CascadeMux I__1020 (
            .O(N__6855),
            .I(N__6848));
    InMux I__1019 (
            .O(N__6854),
            .I(N__6845));
    InMux I__1018 (
            .O(N__6851),
            .I(N__6840));
    InMux I__1017 (
            .O(N__6848),
            .I(N__6840));
    LocalMux I__1016 (
            .O(N__6845),
            .I(\DUT.uart_inst0.rx_clk_divider_1_6 ));
    LocalMux I__1015 (
            .O(N__6840),
            .I(\DUT.uart_inst0.rx_clk_divider_1_6 ));
    InMux I__1014 (
            .O(N__6835),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_5 ));
    InMux I__1013 (
            .O(N__6832),
            .I(N__6829));
    LocalMux I__1012 (
            .O(N__6829),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_7 ));
    InMux I__1011 (
            .O(N__6826),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_6 ));
    InMux I__1010 (
            .O(N__6823),
            .I(bfn_15_2_0_));
    InMux I__1009 (
            .O(N__6820),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_8 ));
    InMux I__1008 (
            .O(N__6817),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_9 ));
    InMux I__1007 (
            .O(N__6814),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_10 ));
    CascadeMux I__1006 (
            .O(N__6811),
            .I(N__6807));
    InMux I__1005 (
            .O(N__6810),
            .I(N__6803));
    InMux I__1004 (
            .O(N__6807),
            .I(N__6797));
    InMux I__1003 (
            .O(N__6806),
            .I(N__6797));
    LocalMux I__1002 (
            .O(N__6803),
            .I(N__6794));
    InMux I__1001 (
            .O(N__6802),
            .I(N__6791));
    LocalMux I__1000 (
            .O(N__6797),
            .I(\DUT.fifo_rx_inst.N_194 ));
    Odrv4 I__999 (
            .O(N__6794),
            .I(\DUT.fifo_rx_inst.N_194 ));
    LocalMux I__998 (
            .O(N__6791),
            .I(\DUT.fifo_rx_inst.N_194 ));
    InMux I__997 (
            .O(N__6784),
            .I(N__6779));
    CascadeMux I__996 (
            .O(N__6783),
            .I(N__6773));
    InMux I__995 (
            .O(N__6782),
            .I(N__6770));
    LocalMux I__994 (
            .O(N__6779),
            .I(N__6767));
    InMux I__993 (
            .O(N__6778),
            .I(N__6764));
    InMux I__992 (
            .O(N__6777),
            .I(N__6757));
    InMux I__991 (
            .O(N__6776),
            .I(N__6757));
    InMux I__990 (
            .O(N__6773),
            .I(N__6757));
    LocalMux I__989 (
            .O(N__6770),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_0 ));
    Odrv4 I__988 (
            .O(N__6767),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_0 ));
    LocalMux I__987 (
            .O(N__6764),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_0 ));
    LocalMux I__986 (
            .O(N__6757),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_0 ));
    InMux I__985 (
            .O(N__6748),
            .I(N__6745));
    LocalMux I__984 (
            .O(N__6745),
            .I(N__6738));
    InMux I__983 (
            .O(N__6744),
            .I(N__6735));
    InMux I__982 (
            .O(N__6743),
            .I(N__6728));
    InMux I__981 (
            .O(N__6742),
            .I(N__6728));
    InMux I__980 (
            .O(N__6741),
            .I(N__6728));
    Odrv4 I__979 (
            .O(N__6738),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_1 ));
    LocalMux I__978 (
            .O(N__6735),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_1 ));
    LocalMux I__977 (
            .O(N__6728),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_1 ));
    InMux I__976 (
            .O(N__6721),
            .I(N__6718));
    LocalMux I__975 (
            .O(N__6718),
            .I(N__6715));
    Span4Mux_v I__974 (
            .O(N__6715),
            .I(N__6712));
    Odrv4 I__973 (
            .O(N__6712),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_5 ));
    InMux I__972 (
            .O(N__6709),
            .I(N__6706));
    LocalMux I__971 (
            .O(N__6706),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_3 ));
    InMux I__970 (
            .O(N__6703),
            .I(N__6700));
    LocalMux I__969 (
            .O(N__6700),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_4 ));
    CEMux I__968 (
            .O(N__6697),
            .I(N__6694));
    LocalMux I__967 (
            .O(N__6694),
            .I(N__6691));
    Span4Mux_v I__966 (
            .O(N__6691),
            .I(N__6686));
    CEMux I__965 (
            .O(N__6690),
            .I(N__6683));
    InMux I__964 (
            .O(N__6689),
            .I(N__6679));
    Span4Mux_h I__963 (
            .O(N__6686),
            .I(N__6674));
    LocalMux I__962 (
            .O(N__6683),
            .I(N__6674));
    CEMux I__961 (
            .O(N__6682),
            .I(N__6671));
    LocalMux I__960 (
            .O(N__6679),
            .I(N__6668));
    Span4Mux_h I__959 (
            .O(N__6674),
            .I(N__6665));
    LocalMux I__958 (
            .O(N__6671),
            .I(N__6660));
    Span4Mux_h I__957 (
            .O(N__6668),
            .I(N__6660));
    Odrv4 I__956 (
            .O(N__6665),
            .I(\DUT.fifo_rx_inst.rFifoData_awe1 ));
    Odrv4 I__955 (
            .O(N__6660),
            .I(\DUT.fifo_rx_inst.rFifoData_awe1 ));
    InMux I__954 (
            .O(N__6655),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_0 ));
    InMux I__953 (
            .O(N__6652),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_1 ));
    CascadeMux I__952 (
            .O(N__6649),
            .I(N__6646));
    InMux I__951 (
            .O(N__6646),
            .I(N__6643));
    LocalMux I__950 (
            .O(N__6643),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_3 ));
    InMux I__949 (
            .O(N__6640),
            .I(N__6636));
    InMux I__948 (
            .O(N__6639),
            .I(N__6633));
    LocalMux I__947 (
            .O(N__6636),
            .I(N__6630));
    LocalMux I__946 (
            .O(N__6633),
            .I(\DUT.uart_inst0.rx_clk_divider_1_3 ));
    Odrv4 I__945 (
            .O(N__6630),
            .I(\DUT.uart_inst0.rx_clk_divider_1_3 ));
    InMux I__944 (
            .O(N__6625),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_2 ));
    CEMux I__943 (
            .O(N__6622),
            .I(N__6619));
    LocalMux I__942 (
            .O(N__6619),
            .I(N__6614));
    CEMux I__941 (
            .O(N__6618),
            .I(N__6610));
    CEMux I__940 (
            .O(N__6617),
            .I(N__6607));
    Span4Mux_h I__939 (
            .O(N__6614),
            .I(N__6604));
    CEMux I__938 (
            .O(N__6613),
            .I(N__6601));
    LocalMux I__937 (
            .O(N__6610),
            .I(N__6598));
    LocalMux I__936 (
            .O(N__6607),
            .I(N__6595));
    Span4Mux_h I__935 (
            .O(N__6604),
            .I(N__6591));
    LocalMux I__934 (
            .O(N__6601),
            .I(N__6588));
    Span4Mux_v I__933 (
            .O(N__6598),
            .I(N__6583));
    Span4Mux_v I__932 (
            .O(N__6595),
            .I(N__6583));
    InMux I__931 (
            .O(N__6594),
            .I(N__6580));
    Odrv4 I__930 (
            .O(N__6591),
            .I(\DUT.fifo_rx_inst.rFifoData_awe2 ));
    Odrv12 I__929 (
            .O(N__6588),
            .I(\DUT.fifo_rx_inst.rFifoData_awe2 ));
    Odrv4 I__928 (
            .O(N__6583),
            .I(\DUT.fifo_rx_inst.rFifoData_awe2 ));
    LocalMux I__927 (
            .O(N__6580),
            .I(\DUT.fifo_rx_inst.rFifoData_awe2 ));
    InMux I__926 (
            .O(N__6571),
            .I(N__6567));
    InMux I__925 (
            .O(N__6570),
            .I(N__6564));
    LocalMux I__924 (
            .O(N__6567),
            .I(\DUT.fifo_rx_inst.rFifoDataro_2 ));
    LocalMux I__923 (
            .O(N__6564),
            .I(\DUT.fifo_rx_inst.rFifoDataro_2 ));
    CEMux I__922 (
            .O(N__6559),
            .I(N__6556));
    LocalMux I__921 (
            .O(N__6556),
            .I(N__6553));
    Span4Mux_h I__920 (
            .O(N__6553),
            .I(N__6549));
    InMux I__919 (
            .O(N__6552),
            .I(N__6546));
    Odrv4 I__918 (
            .O(N__6549),
            .I(\DUT.fifo_tx_inst.rFifoData_awe1 ));
    LocalMux I__917 (
            .O(N__6546),
            .I(\DUT.fifo_tx_inst.rFifoData_awe1 ));
    CascadeMux I__916 (
            .O(N__6541),
            .I(\DUT.fifo_tx_inst.rFifoData_awe3_cascade_ ));
    InMux I__915 (
            .O(N__6538),
            .I(N__6535));
    LocalMux I__914 (
            .O(N__6535),
            .I(\DUT.fifo_tx_inst.un1_i11_i ));
    CascadeMux I__913 (
            .O(N__6532),
            .I(\DUT.fifo_tx_inst.un1_i11_i_cascade_ ));
    InMux I__912 (
            .O(N__6529),
            .I(N__6526));
    LocalMux I__911 (
            .O(N__6526),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_1 ));
    CascadeMux I__910 (
            .O(N__6523),
            .I(N__6520));
    InMux I__909 (
            .O(N__6520),
            .I(N__6517));
    LocalMux I__908 (
            .O(N__6517),
            .I(N__6514));
    Odrv4 I__907 (
            .O(N__6514),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_6 ));
    InMux I__906 (
            .O(N__6511),
            .I(N__6508));
    LocalMux I__905 (
            .O(N__6508),
            .I(N__6505));
    Odrv4 I__904 (
            .O(N__6505),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_7 ));
    CEMux I__903 (
            .O(N__6502),
            .I(N__6497));
    InMux I__902 (
            .O(N__6501),
            .I(N__6494));
    InMux I__901 (
            .O(N__6500),
            .I(N__6491));
    LocalMux I__900 (
            .O(N__6497),
            .I(\DUT.fifo_rx_inst.rFifoData_awe3 ));
    LocalMux I__899 (
            .O(N__6494),
            .I(\DUT.fifo_rx_inst.rFifoData_awe3 ));
    LocalMux I__898 (
            .O(N__6491),
            .I(\DUT.fifo_rx_inst.rFifoData_awe3 ));
    InMux I__897 (
            .O(N__6484),
            .I(N__6480));
    InMux I__896 (
            .O(N__6483),
            .I(N__6477));
    LocalMux I__895 (
            .O(N__6480),
            .I(\DUT.fifo_rx_inst.rFifoDataro_3 ));
    LocalMux I__894 (
            .O(N__6477),
            .I(\DUT.fifo_rx_inst.rFifoDataro_3 ));
    InMux I__893 (
            .O(N__6472),
            .I(N__6469));
    LocalMux I__892 (
            .O(N__6469),
            .I(N__6465));
    InMux I__891 (
            .O(N__6468),
            .I(N__6462));
    Span4Mux_s2_v I__890 (
            .O(N__6465),
            .I(N__6459));
    LocalMux I__889 (
            .O(N__6462),
            .I(\DUT.uart_inst0.recv_stateZ0Z_4 ));
    Odrv4 I__888 (
            .O(N__6459),
            .I(\DUT.uart_inst0.recv_stateZ0Z_4 ));
    CEMux I__887 (
            .O(N__6454),
            .I(N__6451));
    LocalMux I__886 (
            .O(N__6451),
            .I(N__6447));
    CEMux I__885 (
            .O(N__6450),
            .I(N__6444));
    Span4Mux_h I__884 (
            .O(N__6447),
            .I(N__6441));
    LocalMux I__883 (
            .O(N__6444),
            .I(N__6438));
    Odrv4 I__882 (
            .O(N__6441),
            .I(\fifo_inst.ftdi_output_inst.rFifoState_0_1 ));
    Odrv4 I__881 (
            .O(N__6438),
            .I(\fifo_inst.ftdi_output_inst.rFifoState_0_1 ));
    InMux I__880 (
            .O(N__6433),
            .I(N__6430));
    LocalMux I__879 (
            .O(N__6430),
            .I(N__6427));
    Odrv12 I__878 (
            .O(N__6427),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_0 ));
    CascadeMux I__877 (
            .O(N__6424),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ));
    CascadeMux I__876 (
            .O(N__6421),
            .I(N__6418));
    InMux I__875 (
            .O(N__6418),
            .I(N__6415));
    LocalMux I__874 (
            .O(N__6415),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_0 ));
    InMux I__873 (
            .O(N__6412),
            .I(N__6409));
    LocalMux I__872 (
            .O(N__6409),
            .I(N__6406));
    Span4Mux_h I__871 (
            .O(N__6406),
            .I(N__6403));
    Odrv4 I__870 (
            .O(N__6403),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_1 ));
    InMux I__869 (
            .O(N__6400),
            .I(N__6397));
    LocalMux I__868 (
            .O(N__6397),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_0 ));
    InMux I__867 (
            .O(N__6394),
            .I(N__6391));
    LocalMux I__866 (
            .O(N__6391),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_1 ));
    InMux I__865 (
            .O(N__6388),
            .I(N__6382));
    InMux I__864 (
            .O(N__6387),
            .I(N__6382));
    LocalMux I__863 (
            .O(N__6382),
            .I(N__6379));
    Odrv4 I__862 (
            .O(N__6379),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_0 ));
    CascadeMux I__861 (
            .O(N__6376),
            .I(N__6372));
    CascadeMux I__860 (
            .O(N__6375),
            .I(N__6369));
    InMux I__859 (
            .O(N__6372),
            .I(N__6362));
    InMux I__858 (
            .O(N__6369),
            .I(N__6362));
    InMux I__857 (
            .O(N__6368),
            .I(N__6354));
    InMux I__856 (
            .O(N__6367),
            .I(N__6351));
    LocalMux I__855 (
            .O(N__6362),
            .I(N__6348));
    InMux I__854 (
            .O(N__6361),
            .I(N__6337));
    InMux I__853 (
            .O(N__6360),
            .I(N__6337));
    InMux I__852 (
            .O(N__6359),
            .I(N__6337));
    InMux I__851 (
            .O(N__6358),
            .I(N__6337));
    InMux I__850 (
            .O(N__6357),
            .I(N__6337));
    LocalMux I__849 (
            .O(N__6354),
            .I(\DUT.uart_inst0.rx_clk_divider_1_i_3 ));
    LocalMux I__848 (
            .O(N__6351),
            .I(\DUT.uart_inst0.rx_clk_divider_1_i_3 ));
    Odrv4 I__847 (
            .O(N__6348),
            .I(\DUT.uart_inst0.rx_clk_divider_1_i_3 ));
    LocalMux I__846 (
            .O(N__6337),
            .I(\DUT.uart_inst0.rx_clk_divider_1_i_3 ));
    CascadeMux I__845 (
            .O(N__6328),
            .I(N__6321));
    CascadeMux I__844 (
            .O(N__6327),
            .I(N__6318));
    InMux I__843 (
            .O(N__6326),
            .I(N__6313));
    InMux I__842 (
            .O(N__6325),
            .I(N__6308));
    InMux I__841 (
            .O(N__6324),
            .I(N__6308));
    InMux I__840 (
            .O(N__6321),
            .I(N__6299));
    InMux I__839 (
            .O(N__6318),
            .I(N__6299));
    InMux I__838 (
            .O(N__6317),
            .I(N__6299));
    InMux I__837 (
            .O(N__6316),
            .I(N__6299));
    LocalMux I__836 (
            .O(N__6313),
            .I(\DUT.uart_inst0.N_275 ));
    LocalMux I__835 (
            .O(N__6308),
            .I(\DUT.uart_inst0.N_275 ));
    LocalMux I__834 (
            .O(N__6299),
            .I(\DUT.uart_inst0.N_275 ));
    CascadeMux I__833 (
            .O(N__6292),
            .I(\DUT.uart_inst0.N_196_cascade_ ));
    CascadeMux I__832 (
            .O(N__6289),
            .I(\DUT.uart_inst0.N_33_cascade_ ));
    CEMux I__831 (
            .O(N__6286),
            .I(N__6283));
    LocalMux I__830 (
            .O(N__6283),
            .I(N__6280));
    Span4Mux_s3_v I__829 (
            .O(N__6280),
            .I(N__6277));
    Odrv4 I__828 (
            .O(N__6277),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_3_0_c_RNIP8IZ0Z482 ));
    InMux I__827 (
            .O(N__6274),
            .I(N__6271));
    LocalMux I__826 (
            .O(N__6271),
            .I(\DUT.uart_inst0.rx_bits_remaining_RNO_0Z0Z_1 ));
    CascadeMux I__825 (
            .O(N__6268),
            .I(N__6264));
    InMux I__824 (
            .O(N__6267),
            .I(N__6261));
    InMux I__823 (
            .O(N__6264),
            .I(N__6258));
    LocalMux I__822 (
            .O(N__6261),
            .I(\DUT.uart_inst0.g0_8_1 ));
    LocalMux I__821 (
            .O(N__6258),
            .I(\DUT.uart_inst0.g0_8_1 ));
    CEMux I__820 (
            .O(N__6253),
            .I(N__6250));
    LocalMux I__819 (
            .O(N__6250),
            .I(P1A2_c_0_0));
    CascadeMux I__818 (
            .O(N__6247),
            .I(\DUT.uart_inst0.rx_clk_divider_5_i_a2_11_5_cascade_ ));
    InMux I__817 (
            .O(N__6244),
            .I(N__6241));
    LocalMux I__816 (
            .O(N__6241),
            .I(\DUT.uart_inst0.N_221 ));
    CascadeMux I__815 (
            .O(N__6238),
            .I(N__6235));
    InMux I__814 (
            .O(N__6235),
            .I(N__6232));
    LocalMux I__813 (
            .O(N__6232),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_0_0_c_RNOZ0 ));
    CascadeMux I__812 (
            .O(N__6229),
            .I(N__6226));
    InMux I__811 (
            .O(N__6226),
            .I(N__6223));
    LocalMux I__810 (
            .O(N__6223),
            .I(\DUT.uart_inst0.rx_clk_divider_RNIP8N2B_0Z0Z_0 ));
    InMux I__809 (
            .O(N__6220),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_0 ));
    CascadeMux I__808 (
            .O(N__6217),
            .I(N__6214));
    InMux I__807 (
            .O(N__6214),
            .I(N__6211));
    LocalMux I__806 (
            .O(N__6211),
            .I(\DUT.uart_inst0.rx_clk_divider_RNIP8N2B_1Z0Z_0 ));
    InMux I__805 (
            .O(N__6208),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_1 ));
    InMux I__804 (
            .O(N__6205),
            .I(N__6202));
    LocalMux I__803 (
            .O(N__6202),
            .I(N__6199));
    Odrv4 I__802 (
            .O(N__6199),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    CascadeMux I__801 (
            .O(N__6196),
            .I(N__6193));
    InMux I__800 (
            .O(N__6193),
            .I(N__6190));
    LocalMux I__799 (
            .O(N__6190),
            .I(\DUT.uart_inst0.rx_clk_divider_RNIP8N2BZ0Z_0 ));
    InMux I__798 (
            .O(N__6187),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_2 ));
    InMux I__797 (
            .O(N__6184),
            .I(N__6181));
    LocalMux I__796 (
            .O(N__6181),
            .I(\DUT.uart_inst0.rx_clk_divider_RNIP8N2B_2Z0Z_0 ));
    InMux I__795 (
            .O(N__6178),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_3 ));
    InMux I__794 (
            .O(N__6175),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_4 ));
    CascadeMux I__793 (
            .O(N__6172),
            .I(\DUT.uart_inst0.rx_countdown_3_5_cascade_ ));
    InMux I__792 (
            .O(N__6169),
            .I(N__6166));
    LocalMux I__791 (
            .O(N__6166),
            .I(\DUT.uart_inst0.g3_4 ));
    InMux I__790 (
            .O(N__6163),
            .I(N__6160));
    LocalMux I__789 (
            .O(N__6160),
            .I(\DUT.uart_inst0.rx_clk_divider_5_i_a2_1_3 ));
    CascadeMux I__788 (
            .O(N__6157),
            .I(\DUT.uart_inst0.N_222_cascade_ ));
    CascadeMux I__787 (
            .O(N__6154),
            .I(\DUT.uart_inst0.rx_clk_divider_5_i_a2_11_0_5_cascade_ ));
    InMux I__786 (
            .O(N__6151),
            .I(N__6147));
    InMux I__785 (
            .O(N__6150),
            .I(N__6144));
    LocalMux I__784 (
            .O(N__6147),
            .I(\DUT.uart_inst0.rx_clk_divider_5_i_a2_11_5 ));
    LocalMux I__783 (
            .O(N__6144),
            .I(\DUT.uart_inst0.rx_clk_divider_5_i_a2_11_5 ));
    InMux I__782 (
            .O(N__6139),
            .I(N__6136));
    LocalMux I__781 (
            .O(N__6136),
            .I(N__6133));
    Odrv4 I__780 (
            .O(N__6133),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_2 ));
    InMux I__779 (
            .O(N__6130),
            .I(N__6127));
    LocalMux I__778 (
            .O(N__6127),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_3 ));
    InMux I__777 (
            .O(N__6124),
            .I(N__6121));
    LocalMux I__776 (
            .O(N__6121),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_4 ));
    CEMux I__775 (
            .O(N__6118),
            .I(N__6115));
    LocalMux I__774 (
            .O(N__6115),
            .I(N__6110));
    CEMux I__773 (
            .O(N__6114),
            .I(N__6107));
    CEMux I__772 (
            .O(N__6113),
            .I(N__6104));
    Span4Mux_h I__771 (
            .O(N__6110),
            .I(N__6097));
    LocalMux I__770 (
            .O(N__6107),
            .I(N__6097));
    LocalMux I__769 (
            .O(N__6104),
            .I(N__6094));
    CEMux I__768 (
            .O(N__6103),
            .I(N__6091));
    InMux I__767 (
            .O(N__6102),
            .I(N__6088));
    Span4Mux_h I__766 (
            .O(N__6097),
            .I(N__6085));
    Sp12to4 I__765 (
            .O(N__6094),
            .I(N__6078));
    LocalMux I__764 (
            .O(N__6091),
            .I(N__6078));
    LocalMux I__763 (
            .O(N__6088),
            .I(N__6078));
    Odrv4 I__762 (
            .O(N__6085),
            .I(\DUT.fifo_rx_inst.rFifoData_awe0 ));
    Odrv12 I__761 (
            .O(N__6078),
            .I(\DUT.fifo_rx_inst.rFifoData_awe0 ));
    InMux I__760 (
            .O(N__6073),
            .I(N__6070));
    LocalMux I__759 (
            .O(N__6070),
            .I(N__6067));
    Odrv4 I__758 (
            .O(N__6067),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_2 ));
    InMux I__757 (
            .O(N__6064),
            .I(N__6061));
    LocalMux I__756 (
            .O(N__6061),
            .I(N__6058));
    Odrv4 I__755 (
            .O(N__6058),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_5 ));
    CascadeMux I__754 (
            .O(N__6055),
            .I(\DUT.fifo_rx_inst.N_194_cascade_ ));
    InMux I__753 (
            .O(N__6052),
            .I(N__6049));
    LocalMux I__752 (
            .O(N__6049),
            .I(N__6046));
    Odrv4 I__751 (
            .O(N__6046),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_2 ));
    InMux I__750 (
            .O(N__6043),
            .I(N__6040));
    LocalMux I__749 (
            .O(N__6040),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_2 ));
    CascadeMux I__748 (
            .O(N__6037),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2_cascade_ ));
    InMux I__747 (
            .O(N__6034),
            .I(N__6031));
    LocalMux I__746 (
            .O(N__6031),
            .I(N__6028));
    Odrv4 I__745 (
            .O(N__6028),
            .I(\DUT.rFifoDatarx_0_2 ));
    CascadeMux I__744 (
            .O(N__6025),
            .I(\DUT.rFifoDataror_0_0_cascade_ ));
    InMux I__743 (
            .O(N__6022),
            .I(N__6019));
    LocalMux I__742 (
            .O(N__6019),
            .I(\DUT.rFifoDataror_1 ));
    InMux I__741 (
            .O(N__6016),
            .I(N__6002));
    InMux I__740 (
            .O(N__6015),
            .I(N__6002));
    InMux I__739 (
            .O(N__6014),
            .I(N__6002));
    InMux I__738 (
            .O(N__6013),
            .I(N__5991));
    InMux I__737 (
            .O(N__6012),
            .I(N__5991));
    InMux I__736 (
            .O(N__6011),
            .I(N__5991));
    InMux I__735 (
            .O(N__6010),
            .I(N__5991));
    InMux I__734 (
            .O(N__6009),
            .I(N__5991));
    LocalMux I__733 (
            .O(N__6002),
            .I(N__5986));
    LocalMux I__732 (
            .O(N__5991),
            .I(N__5986));
    Odrv4 I__731 (
            .O(N__5986),
            .I(\DUT.uart_inst0.N_257 ));
    InMux I__730 (
            .O(N__5983),
            .I(N__5980));
    LocalMux I__729 (
            .O(N__5980),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_3 ));
    InMux I__728 (
            .O(N__5977),
            .I(N__5974));
    LocalMux I__727 (
            .O(N__5974),
            .I(N__5971));
    Odrv4 I__726 (
            .O(N__5971),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_3 ));
    CascadeMux I__725 (
            .O(N__5968),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ));
    InMux I__724 (
            .O(N__5965),
            .I(N__5962));
    LocalMux I__723 (
            .O(N__5962),
            .I(N__5959));
    Odrv4 I__722 (
            .O(N__5959),
            .I(\DUT.rFifoDatarx_3 ));
    CascadeMux I__721 (
            .O(N__5956),
            .I(N__5950));
    InMux I__720 (
            .O(N__5955),
            .I(N__5938));
    InMux I__719 (
            .O(N__5954),
            .I(N__5933));
    InMux I__718 (
            .O(N__5953),
            .I(N__5933));
    InMux I__717 (
            .O(N__5950),
            .I(N__5930));
    InMux I__716 (
            .O(N__5949),
            .I(N__5925));
    InMux I__715 (
            .O(N__5948),
            .I(N__5925));
    InMux I__714 (
            .O(N__5947),
            .I(N__5920));
    InMux I__713 (
            .O(N__5946),
            .I(N__5920));
    InMux I__712 (
            .O(N__5945),
            .I(N__5915));
    InMux I__711 (
            .O(N__5944),
            .I(N__5915));
    InMux I__710 (
            .O(N__5943),
            .I(N__5908));
    InMux I__709 (
            .O(N__5942),
            .I(N__5908));
    InMux I__708 (
            .O(N__5941),
            .I(N__5908));
    LocalMux I__707 (
            .O(N__5938),
            .I(N__5903));
    LocalMux I__706 (
            .O(N__5933),
            .I(N__5903));
    LocalMux I__705 (
            .O(N__5930),
            .I(N__5900));
    LocalMux I__704 (
            .O(N__5925),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__703 (
            .O(N__5920),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__702 (
            .O(N__5915),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__701 (
            .O(N__5908),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    Odrv4 I__700 (
            .O(N__5903),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    Odrv4 I__699 (
            .O(N__5900),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    CascadeMux I__698 (
            .O(N__5887),
            .I(N__5882));
    CascadeMux I__697 (
            .O(N__5886),
            .I(N__5871));
    CascadeMux I__696 (
            .O(N__5885),
            .I(N__5866));
    InMux I__695 (
            .O(N__5882),
            .I(N__5862));
    CascadeMux I__694 (
            .O(N__5881),
            .I(N__5858));
    CascadeMux I__693 (
            .O(N__5880),
            .I(N__5855));
    CascadeMux I__692 (
            .O(N__5879),
            .I(N__5848));
    CascadeMux I__691 (
            .O(N__5878),
            .I(N__5844));
    CascadeMux I__690 (
            .O(N__5877),
            .I(N__5841));
    CascadeMux I__689 (
            .O(N__5876),
            .I(N__5838));
    InMux I__688 (
            .O(N__5875),
            .I(N__5831));
    InMux I__687 (
            .O(N__5874),
            .I(N__5831));
    InMux I__686 (
            .O(N__5871),
            .I(N__5831));
    InMux I__685 (
            .O(N__5870),
            .I(N__5822));
    InMux I__684 (
            .O(N__5869),
            .I(N__5822));
    InMux I__683 (
            .O(N__5866),
            .I(N__5822));
    InMux I__682 (
            .O(N__5865),
            .I(N__5822));
    LocalMux I__681 (
            .O(N__5862),
            .I(N__5819));
    InMux I__680 (
            .O(N__5861),
            .I(N__5814));
    InMux I__679 (
            .O(N__5858),
            .I(N__5814));
    InMux I__678 (
            .O(N__5855),
            .I(N__5811));
    InMux I__677 (
            .O(N__5854),
            .I(N__5800));
    InMux I__676 (
            .O(N__5853),
            .I(N__5800));
    InMux I__675 (
            .O(N__5852),
            .I(N__5800));
    InMux I__674 (
            .O(N__5851),
            .I(N__5800));
    InMux I__673 (
            .O(N__5848),
            .I(N__5800));
    InMux I__672 (
            .O(N__5847),
            .I(N__5793));
    InMux I__671 (
            .O(N__5844),
            .I(N__5793));
    InMux I__670 (
            .O(N__5841),
            .I(N__5793));
    InMux I__669 (
            .O(N__5838),
            .I(N__5790));
    LocalMux I__668 (
            .O(N__5831),
            .I(N__5787));
    LocalMux I__667 (
            .O(N__5822),
            .I(N__5784));
    Odrv4 I__666 (
            .O(N__5819),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__665 (
            .O(N__5814),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__664 (
            .O(N__5811),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__663 (
            .O(N__5800),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__662 (
            .O(N__5793),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__661 (
            .O(N__5790),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    Odrv4 I__660 (
            .O(N__5787),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    Odrv4 I__659 (
            .O(N__5784),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    InMux I__658 (
            .O(N__5767),
            .I(N__5764));
    LocalMux I__657 (
            .O(N__5764),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4 ));
    InMux I__656 (
            .O(N__5761),
            .I(N__5758));
    LocalMux I__655 (
            .O(N__5758),
            .I(wRxFifoData_3));
    InMux I__654 (
            .O(N__5755),
            .I(N__5752));
    LocalMux I__653 (
            .O(N__5752),
            .I(N__5749));
    Span4Mux_h I__652 (
            .O(N__5749),
            .I(N__5746));
    Odrv4 I__651 (
            .O(N__5746),
            .I(\DUT.rFifoDatarx_0_5 ));
    CascadeMux I__650 (
            .O(N__5743),
            .I(N__5740));
    InMux I__649 (
            .O(N__5740),
            .I(N__5737));
    LocalMux I__648 (
            .O(N__5737),
            .I(wRxFifoData_5));
    InMux I__647 (
            .O(N__5734),
            .I(N__5731));
    LocalMux I__646 (
            .O(N__5731),
            .I(\DUT.rFifoDatarx_0_7 ));
    CascadeMux I__645 (
            .O(N__5728),
            .I(N__5725));
    InMux I__644 (
            .O(N__5725),
            .I(N__5722));
    LocalMux I__643 (
            .O(N__5722),
            .I(wRxFifoData_7));
    CEMux I__642 (
            .O(N__5719),
            .I(N__5715));
    CEMux I__641 (
            .O(N__5718),
            .I(N__5712));
    LocalMux I__640 (
            .O(N__5715),
            .I(N__5709));
    LocalMux I__639 (
            .O(N__5712),
            .I(N__5706));
    Odrv4 I__638 (
            .O(N__5709),
            .I(un1_oRxFlag_0_i_0));
    Odrv4 I__637 (
            .O(N__5706),
            .I(un1_oRxFlag_0_i_0));
    CascadeMux I__636 (
            .O(N__5701),
            .I(\DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1_cascade_ ));
    InMux I__635 (
            .O(N__5698),
            .I(N__5695));
    LocalMux I__634 (
            .O(N__5695),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_1 ));
    InMux I__633 (
            .O(N__5692),
            .I(N__5689));
    LocalMux I__632 (
            .O(N__5689),
            .I(N__5686));
    Odrv4 I__631 (
            .O(N__5686),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1 ));
    InMux I__630 (
            .O(N__5683),
            .I(N__5680));
    LocalMux I__629 (
            .O(N__5680),
            .I(\DUT.rFifoDatarx_0_1 ));
    InMux I__628 (
            .O(N__5677),
            .I(N__5674));
    LocalMux I__627 (
            .O(N__5674),
            .I(\DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1 ));
    InMux I__626 (
            .O(N__5671),
            .I(N__5665));
    InMux I__625 (
            .O(N__5670),
            .I(N__5665));
    LocalMux I__624 (
            .O(N__5665),
            .I(N__5658));
    InMux I__623 (
            .O(N__5664),
            .I(N__5653));
    InMux I__622 (
            .O(N__5663),
            .I(N__5653));
    InMux I__621 (
            .O(N__5662),
            .I(N__5650));
    InMux I__620 (
            .O(N__5661),
            .I(N__5647));
    Span4Mux_v I__619 (
            .O(N__5658),
            .I(N__5642));
    LocalMux I__618 (
            .O(N__5653),
            .I(N__5642));
    LocalMux I__617 (
            .O(N__5650),
            .I(\DUT.wRcvd ));
    LocalMux I__616 (
            .O(N__5647),
            .I(\DUT.wRcvd ));
    Odrv4 I__615 (
            .O(N__5642),
            .I(\DUT.wRcvd ));
    InMux I__614 (
            .O(N__5635),
            .I(N__5629));
    InMux I__613 (
            .O(N__5634),
            .I(N__5629));
    LocalMux I__612 (
            .O(N__5629),
            .I(N__5625));
    InMux I__611 (
            .O(N__5628),
            .I(N__5618));
    Span4Mux_v I__610 (
            .O(N__5625),
            .I(N__5615));
    InMux I__609 (
            .O(N__5624),
            .I(N__5610));
    InMux I__608 (
            .O(N__5623),
            .I(N__5610));
    InMux I__607 (
            .O(N__5622),
            .I(N__5605));
    InMux I__606 (
            .O(N__5621),
            .I(N__5605));
    LocalMux I__605 (
            .O(N__5618),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ));
    Odrv4 I__604 (
            .O(N__5615),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ));
    LocalMux I__603 (
            .O(N__5610),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ));
    LocalMux I__602 (
            .O(N__5605),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ));
    CascadeMux I__601 (
            .O(N__5596),
            .I(N__5592));
    InMux I__600 (
            .O(N__5595),
            .I(N__5586));
    InMux I__599 (
            .O(N__5592),
            .I(N__5583));
    InMux I__598 (
            .O(N__5591),
            .I(N__5580));
    InMux I__597 (
            .O(N__5590),
            .I(N__5575));
    InMux I__596 (
            .O(N__5589),
            .I(N__5575));
    LocalMux I__595 (
            .O(N__5586),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_1 ));
    LocalMux I__594 (
            .O(N__5583),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_1 ));
    LocalMux I__593 (
            .O(N__5580),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_1 ));
    LocalMux I__592 (
            .O(N__5575),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_1 ));
    InMux I__591 (
            .O(N__5566),
            .I(N__5556));
    InMux I__590 (
            .O(N__5565),
            .I(N__5556));
    InMux I__589 (
            .O(N__5564),
            .I(N__5556));
    CascadeMux I__588 (
            .O(N__5563),
            .I(N__5552));
    LocalMux I__587 (
            .O(N__5556),
            .I(N__5549));
    CascadeMux I__586 (
            .O(N__5555),
            .I(N__5546));
    InMux I__585 (
            .O(N__5552),
            .I(N__5543));
    Span4Mux_v I__584 (
            .O(N__5549),
            .I(N__5540));
    InMux I__583 (
            .O(N__5546),
            .I(N__5537));
    LocalMux I__582 (
            .O(N__5543),
            .I(\DUT.fifo_rx_inst.N_148 ));
    Odrv4 I__581 (
            .O(N__5540),
            .I(\DUT.fifo_rx_inst.N_148 ));
    LocalMux I__580 (
            .O(N__5537),
            .I(\DUT.fifo_rx_inst.N_148 ));
    InMux I__579 (
            .O(N__5530),
            .I(N__5527));
    LocalMux I__578 (
            .O(N__5527),
            .I(N__5524));
    Span4Mux_v I__577 (
            .O(N__5524),
            .I(N__5521));
    Sp12to4 I__576 (
            .O(N__5521),
            .I(N__5518));
    Span12Mux_h I__575 (
            .O(N__5518),
            .I(N__5515));
    Span12Mux_v I__574 (
            .O(N__5515),
            .I(N__5512));
    Odrv12 I__573 (
            .O(N__5512),
            .I(ioFifoData_in_7));
    InMux I__572 (
            .O(N__5509),
            .I(N__5506));
    LocalMux I__571 (
            .O(N__5506),
            .I(N__5503));
    Span4Mux_h I__570 (
            .O(N__5503),
            .I(N__5500));
    Span4Mux_v I__569 (
            .O(N__5500),
            .I(N__5497));
    Odrv4 I__568 (
            .O(N__5497),
            .I(ioFifoData_in_1));
    InMux I__567 (
            .O(N__5494),
            .I(N__5491));
    LocalMux I__566 (
            .O(N__5491),
            .I(N__5488));
    Span4Mux_h I__565 (
            .O(N__5488),
            .I(N__5485));
    Span4Mux_h I__564 (
            .O(N__5485),
            .I(N__5482));
    Span4Mux_v I__563 (
            .O(N__5482),
            .I(N__5479));
    Odrv4 I__562 (
            .O(N__5479),
            .I(ioFifoData_in_3));
    InMux I__561 (
            .O(N__5476),
            .I(N__5473));
    LocalMux I__560 (
            .O(N__5473),
            .I(N__5470));
    Span4Mux_v I__559 (
            .O(N__5470),
            .I(N__5467));
    Span4Mux_h I__558 (
            .O(N__5467),
            .I(N__5464));
    Odrv4 I__557 (
            .O(N__5464),
            .I(ioFifoData_in_5));
    InMux I__556 (
            .O(N__5461),
            .I(N__5458));
    LocalMux I__555 (
            .O(N__5458),
            .I(N__5455));
    Span4Mux_v I__554 (
            .O(N__5455),
            .I(N__5452));
    Span4Mux_h I__553 (
            .O(N__5452),
            .I(N__5449));
    Span4Mux_h I__552 (
            .O(N__5449),
            .I(N__5446));
    Odrv4 I__551 (
            .O(N__5446),
            .I(ioFifoData_in_2));
    CascadeMux I__550 (
            .O(N__5443),
            .I(N__5440));
    InMux I__549 (
            .O(N__5440),
            .I(N__5437));
    LocalMux I__548 (
            .O(N__5437),
            .I(wRxFifoData_1));
    CascadeMux I__547 (
            .O(N__5434),
            .I(N__5431));
    InMux I__546 (
            .O(N__5431),
            .I(N__5428));
    LocalMux I__545 (
            .O(N__5428),
            .I(N__5425));
    Odrv4 I__544 (
            .O(N__5425),
            .I(wRxFifoData_2));
    CascadeMux I__543 (
            .O(N__5422),
            .I(\DUT.uart_inst0.g0_0_5_cascade_ ));
    CascadeMux I__542 (
            .O(N__5419),
            .I(\DUT.uart_inst0.g0_6_cascade_ ));
    InMux I__541 (
            .O(N__5416),
            .I(N__5413));
    LocalMux I__540 (
            .O(N__5413),
            .I(N__5410));
    Odrv4 I__539 (
            .O(N__5410),
            .I(\DUT.uart_inst0.g0_1_0 ));
    CascadeMux I__538 (
            .O(N__5407),
            .I(\DUT.uart_inst0.g3_0_cascade_ ));
    InMux I__537 (
            .O(N__5404),
            .I(N__5401));
    LocalMux I__536 (
            .O(N__5401),
            .I(\DUT.uart_inst0.g0_0_4 ));
    InMux I__535 (
            .O(N__5398),
            .I(N__5395));
    LocalMux I__534 (
            .O(N__5395),
            .I(N__5392));
    Odrv4 I__533 (
            .O(N__5392),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_4 ));
    IoInMux I__532 (
            .O(N__5389),
            .I(N__5386));
    LocalMux I__531 (
            .O(N__5386),
            .I(wPllLocked_i));
    CascadeMux I__530 (
            .O(N__5383),
            .I(\DUT.uart_inst0.N_275_cascade_ ));
    CascadeMux I__529 (
            .O(N__5380),
            .I(\DUT.fifo_rx_inst.rReadPtr_RNIDU4H2Z0Z_0_cascade_ ));
    InMux I__528 (
            .O(N__5377),
            .I(N__5374));
    LocalMux I__527 (
            .O(N__5374),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_6 ));
    InMux I__526 (
            .O(N__5371),
            .I(N__5368));
    LocalMux I__525 (
            .O(N__5368),
            .I(N__5365));
    Odrv4 I__524 (
            .O(N__5365),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6 ));
    InMux I__523 (
            .O(N__5362),
            .I(N__5359));
    LocalMux I__522 (
            .O(N__5359),
            .I(\DUT.fifo_rx_inst.rReadPtr_RNIDU4H2Z0Z_0 ));
    CascadeMux I__521 (
            .O(N__5356),
            .I(N__5353));
    InMux I__520 (
            .O(N__5353),
            .I(N__5350));
    LocalMux I__519 (
            .O(N__5350),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_4 ));
    InMux I__518 (
            .O(N__5347),
            .I(N__5344));
    LocalMux I__517 (
            .O(N__5344),
            .I(N__5341));
    Odrv4 I__516 (
            .O(N__5341),
            .I(\DUT.rFifoDatarx_0_4 ));
    InMux I__515 (
            .O(N__5338),
            .I(N__5335));
    LocalMux I__514 (
            .O(N__5335),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_5 ));
    CascadeMux I__513 (
            .O(N__5332),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ));
    InMux I__512 (
            .O(N__5329),
            .I(N__5326));
    LocalMux I__511 (
            .O(N__5326),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_5 ));
    InMux I__510 (
            .O(N__5323),
            .I(N__5320));
    LocalMux I__509 (
            .O(N__5320),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_6 ));
    InMux I__508 (
            .O(N__5317),
            .I(N__5313));
    InMux I__507 (
            .O(N__5316),
            .I(N__5310));
    LocalMux I__506 (
            .O(N__5313),
            .I(N__5305));
    LocalMux I__505 (
            .O(N__5310),
            .I(N__5305));
    Odrv4 I__504 (
            .O(N__5305),
            .I(\DUT.fifo_rx_inst.rFifoDataro_0 ));
    InMux I__503 (
            .O(N__5302),
            .I(N__5298));
    InMux I__502 (
            .O(N__5301),
            .I(N__5295));
    LocalMux I__501 (
            .O(N__5298),
            .I(\DUT.fifo_rx_inst.rFifoDataro_1 ));
    LocalMux I__500 (
            .O(N__5295),
            .I(\DUT.fifo_rx_inst.rFifoDataro_1 ));
    InMux I__499 (
            .O(N__5290),
            .I(N__5287));
    LocalMux I__498 (
            .O(N__5287),
            .I(N__5284));
    Odrv4 I__497 (
            .O(N__5284),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_0 ));
    InMux I__496 (
            .O(N__5281),
            .I(N__5278));
    LocalMux I__495 (
            .O(N__5278),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_6 ));
    InMux I__494 (
            .O(N__5275),
            .I(N__5272));
    LocalMux I__493 (
            .O(N__5272),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_7 ));
    InMux I__492 (
            .O(N__5269),
            .I(N__5266));
    LocalMux I__491 (
            .O(N__5266),
            .I(N__5263));
    Sp12to4 I__490 (
            .O(N__5263),
            .I(N__5260));
    Odrv12 I__489 (
            .O(N__5260),
            .I(ioFifoData_in_0));
    InMux I__488 (
            .O(N__5257),
            .I(N__5254));
    LocalMux I__487 (
            .O(N__5254),
            .I(N__5251));
    Span4Mux_h I__486 (
            .O(N__5251),
            .I(N__5248));
    Span4Mux_h I__485 (
            .O(N__5248),
            .I(N__5245));
    Span4Mux_v I__484 (
            .O(N__5245),
            .I(N__5242));
    Odrv4 I__483 (
            .O(N__5242),
            .I(ioFifoData_in_4));
    CascadeMux I__482 (
            .O(N__5239),
            .I(N__5236));
    InMux I__481 (
            .O(N__5236),
            .I(N__5233));
    LocalMux I__480 (
            .O(N__5233),
            .I(wRxFifoData_0));
    InMux I__479 (
            .O(N__5230),
            .I(N__5227));
    LocalMux I__478 (
            .O(N__5227),
            .I(\DUT.rFifoDatarx_0 ));
    CascadeMux I__477 (
            .O(N__5224),
            .I(N__5221));
    InMux I__476 (
            .O(N__5221),
            .I(N__5218));
    LocalMux I__475 (
            .O(N__5218),
            .I(wRxFifoData_4));
    CascadeMux I__474 (
            .O(N__5215),
            .I(N__5212));
    InMux I__473 (
            .O(N__5212),
            .I(N__5209));
    LocalMux I__472 (
            .O(N__5209),
            .I(wRxFifoData_6));
    InMux I__471 (
            .O(N__5206),
            .I(N__5203));
    LocalMux I__470 (
            .O(N__5203),
            .I(\DUT.rFifoDatarx_6 ));
    InMux I__469 (
            .O(N__5200),
            .I(N__5197));
    LocalMux I__468 (
            .O(N__5197),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_7 ));
    CascadeMux I__467 (
            .O(N__5194),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7_cascade_ ));
    InMux I__466 (
            .O(N__5191),
            .I(N__5188));
    LocalMux I__465 (
            .O(N__5188),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_7 ));
    InMux I__464 (
            .O(N__5185),
            .I(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0 ));
    InMux I__463 (
            .O(N__5182),
            .I(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1 ));
    CascadeMux I__462 (
            .O(N__5179),
            .I(un1_oRxFlag_0_i_cascade_));
    InMux I__461 (
            .O(N__5176),
            .I(N__5173));
    LocalMux I__460 (
            .O(N__5173),
            .I(\DUT.fifo_rx_inst.rFifoCount_RNITA8H2Z0Z_1 ));
    CascadeMux I__459 (
            .O(N__5170),
            .I(rFifoCount_RNIHH0D1_0_cascade_));
    InMux I__458 (
            .O(N__5167),
            .I(N__5164));
    LocalMux I__457 (
            .O(N__5164),
            .I(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0 ));
    InMux I__456 (
            .O(N__5161),
            .I(N__5158));
    LocalMux I__455 (
            .O(N__5158),
            .I(N__5155));
    Span4Mux_v I__454 (
            .O(N__5155),
            .I(N__5152));
    Sp12to4 I__453 (
            .O(N__5152),
            .I(N__5149));
    Span12Mux_h I__452 (
            .O(N__5149),
            .I(N__5146));
    Span12Mux_v I__451 (
            .O(N__5146),
            .I(N__5143));
    Odrv12 I__450 (
            .O(N__5143),
            .I(ioFifoData_in_6));
    CascadeMux I__449 (
            .O(N__5140),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ));
    CascadeMux I__448 (
            .O(N__5137),
            .I(N__5134));
    InMux I__447 (
            .O(N__5134),
            .I(N__5131));
    LocalMux I__446 (
            .O(N__5131),
            .I(N__5128));
    Odrv4 I__445 (
            .O(N__5128),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_0 ));
    InMux I__444 (
            .O(N__5125),
            .I(N__5122));
    LocalMux I__443 (
            .O(N__5122),
            .I(N__5119));
    Odrv4 I__442 (
            .O(N__5119),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_1 ));
    InMux I__441 (
            .O(N__5116),
            .I(N__5113));
    LocalMux I__440 (
            .O(N__5113),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_1 ));
    InMux I__439 (
            .O(N__5110),
            .I(N__5107));
    LocalMux I__438 (
            .O(N__5107),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_0 ));
    InMux I__437 (
            .O(N__5104),
            .I(N__5101));
    LocalMux I__436 (
            .O(N__5101),
            .I(N__5098));
    Odrv4 I__435 (
            .O(N__5098),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_0 ));
    InMux I__434 (
            .O(N__5095),
            .I(N__5092));
    LocalMux I__433 (
            .O(N__5092),
            .I(\PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO ));
    IoInMux I__432 (
            .O(N__5089),
            .I(N__5086));
    LocalMux I__431 (
            .O(N__5086),
            .I(N__5083));
    Span12Mux_s9_v I__430 (
            .O(N__5083),
            .I(N__5080));
    Span12Mux_v I__429 (
            .O(N__5080),
            .I(N__5077));
    Odrv12 I__428 (
            .O(N__5077),
            .I(BTN_N_c));
    defparam IN_MUX_bfv_21_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_9_0_));
    defparam IN_MUX_bfv_21_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_10_0_ (
            .carryinitin(\DUT.uart_inst0.tx_clk_divider_cry_7 ),
            .carryinitout(bfn_21_10_0_));
    defparam IN_MUX_bfv_14_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_3_0_));
    defparam IN_MUX_bfv_15_1_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_1_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_1_0_));
    defparam IN_MUX_bfv_15_2_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_2_0_ (
            .carryinitin(\DUT.uart_inst0.rx_clk_divider_1_cry_7 ),
            .carryinitout(bfn_15_2_0_));
    defparam IN_MUX_bfv_15_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_3_0_ (
            .carryinitin(\DUT.uart_inst0.rx_clk_divider_1_cry_15 ),
            .carryinitout(bfn_15_3_0_));
    defparam IN_MUX_bfv_16_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_11_0_));
    defparam IN_MUX_bfv_12_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_4_0_));
    ICE_GB wPllLocked_i_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__5389),
            .GLOBALBUFFEROUTPUT(wPllLocked_i_g));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB \top_pll_inst.top_pll_inst_RNISDA2  (
            .USERSIGNALTOGLOBALBUFFER(N__10639),
            .GLOBALBUFFEROUTPUT(wPllLocked_g));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0 .C_ON=1'b0;
    defparam \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0 .SEQ_MODE=4'b0000;
    defparam \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5095),
            .lcout(wPllLocked),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_10_5_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_10_5_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_10_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_10_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7330),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12807),
            .ce(N__10080),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_10_6_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_10_6_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_10_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_10_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7372),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12801),
            .ce(N__7414),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_10_7_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_10_7_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_10_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_10_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7582),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12793),
            .ce(N__10071),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_LC_10_8_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_LC_10_8_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_LC_10_8_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_0_LC_10_8_0  (
            .in0(_gnd_net_),
            .in1(N__6102),
            .in2(_gnd_net_),
            .in3(N__5317),
            .lcout(\DUT.fifo_rx_inst.rFifoDataro_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12788),
            .ce(),
            .sr(N__11116));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_10_9_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_10_9_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_10_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_10_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7591),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12782),
            .ce(N__7412),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_11_6_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_11_6_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_11_6_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_11_6_5  (
            .in0(_gnd_net_),
            .in1(N__7241),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12794),
            .ce(N__6697),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_1_LC_11_7_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_1_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_1_LC_11_7_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_1_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(N__5302),
            .in2(_gnd_net_),
            .in3(N__6689),
            .lcout(\DUT.fifo_rx_inst.rFifoDataro_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12789),
            .ce(),
            .sr(N__11117));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_11_8_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_11_8_0 .LUT_INIT=16'b0011001101000111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_11_8_0  (
            .in0(N__5110),
            .in1(N__5954),
            .in2(N__5137),
            .in3(N__5874),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI5EJ22_0_LC_11_8_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI5EJ22_0_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI5EJ22_0_LC_11_8_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI5EJ22_0_LC_11_8_1  (
            .in0(N__5875),
            .in1(N__5290),
            .in2(N__5140),
            .in3(N__5104),
            .lcout(\DUT.rFifoDatarx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_11_8_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_11_8_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_11_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7192),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12783),
            .ce(N__6113),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_11_8_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_11_8_3 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_11_8_3  (
            .in0(N__5953),
            .in1(N__5125),
            .in2(N__5886),
            .in3(N__5116),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_11_8_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_11_8_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_11_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7246),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12783),
            .ce(N__6113),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_11_9_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_11_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8461),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12778),
            .ce(N__6690),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_11_9_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_11_9_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_11_9_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_11_9_2  (
            .in0(N__7024),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12778),
            .ce(N__6690),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_11_9_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_11_9_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_11_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7194),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12778),
            .ce(N__6690),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_11_9_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_11_9_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_11_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7068),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12778),
            .ce(N__6690),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_11_10_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_11_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7198),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12775),
            .ce(N__6618),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_LC_12_4_0 .C_ON=1'b1;
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_LC_12_4_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_LC_12_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_LC_12_4_0  (
            .in0(_gnd_net_),
            .in1(N__5167),
            .in2(N__10417),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_4_0_),
            .carryout(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_1_LC_12_4_1 .C_ON=1'b1;
    defparam \DUT.fifo_rx_inst.rFifoCount_1_LC_12_4_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoCount_1_LC_12_4_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_1_LC_12_4_1  (
            .in0(_gnd_net_),
            .in1(N__5176),
            .in2(N__5596),
            .in3(N__5185),
            .lcout(\DUT.fifo_rx_inst.rFifoCountZ0Z_1 ),
            .ltout(),
            .carryin(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0 ),
            .carryout(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1 ),
            .clk(N__12800),
            .ce(),
            .sr(N__11124));
    defparam \DUT.fifo_rx_inst.rFifoCount_2_LC_12_4_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_2_LC_12_4_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoCount_2_LC_12_4_2 .LUT_INIT=16'b0011011011001001;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_2_LC_12_4_2  (
            .in0(N__5662),
            .in1(N__5628),
            .in2(N__5563),
            .in3(N__5182),
            .lcout(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12800),
            .ce(),
            .sr(N__11124));
    defparam \DUT.uart_inst0.un1_oRxFlag_0_i_LC_12_5_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.un1_oRxFlag_0_i_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.un1_oRxFlag_0_i_LC_12_5_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.uart_inst0.un1_oRxFlag_0_i_LC_12_5_0  (
            .in0(_gnd_net_),
            .in1(N__10322),
            .in2(_gnd_net_),
            .in3(N__10233),
            .lcout(),
            .ltout(un1_oRxFlag_0_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rTxByte_esr_ctle_7_LC_12_5_1.C_ON=1'b0;
    defparam rTxByte_esr_ctle_7_LC_12_5_1.SEQ_MODE=4'b0000;
    defparam rTxByte_esr_ctle_7_LC_12_5_1.LUT_INIT=16'b1111101011111010;
    LogicCell40 rTxByte_esr_ctle_7_LC_12_5_1 (
            .in0(N__11146),
            .in1(_gnd_net_),
            .in2(N__5179),
            .in3(_gnd_net_),
            .lcout(un1_oRxFlag_0_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNITA8H2_1_LC_12_5_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNITA8H2_1_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNITA8H2_1_LC_12_5_3 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNITA8H2_1_LC_12_5_3  (
            .in0(N__5664),
            .in1(_gnd_net_),
            .in2(N__5555),
            .in3(N__5595),
            .lcout(\DUT.fifo_rx_inst.rFifoCount_RNITA8H2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_LC_12_5_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_LC_12_5_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_LC_12_5_4  (
            .in0(N__10404),
            .in1(N__5591),
            .in2(_gnd_net_),
            .in3(N__5622),
            .lcout(rFifoCount_RNIHH0D1_0),
            .ltout(rFifoCount_RNIHH0D1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_12_5_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_12_5_5 .LUT_INIT=16'b0000000011110011;
    LogicCell40 \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_12_5_5  (
            .in0(N__10412),
            .in1(N__10451),
            .in2(N__5170),
            .in3(N__10428),
            .lcout(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIDQ741_2_LC_12_5_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIDQ741_2_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIDQ741_2_LC_12_5_6 .LUT_INIT=16'b1101110110011001;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNIDQ741_2_LC_12_5_6  (
            .in0(N__10450),
            .in1(N__5663),
            .in2(_gnd_net_),
            .in3(N__5621),
            .lcout(\DUT.fifo_rx_inst.N_206 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_6_LC_12_6_3 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_6_LC_12_6_3 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_6_LC_12_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rRxData_esr_6_LC_12_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5161),
            .lcout(wRxFifoData_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12787),
            .ce(N__6454),
            .sr(N__11115));
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_0_LC_12_6_4 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_0_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_0_LC_12_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rRxData_esr_0_LC_12_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5269),
            .lcout(wRxFifoData_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12787),
            .ce(N__6454),
            .sr(N__11115));
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_4_LC_12_6_6 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_4_LC_12_6_6 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_4_LC_12_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rRxData_esr_4_LC_12_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5257),
            .lcout(wRxFifoData_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12787),
            .ce(N__6454),
            .sr(N__11115));
    defparam rTxByte_esr_0_LC_12_7_0.C_ON=1'b0;
    defparam rTxByte_esr_0_LC_12_7_0.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_0_LC_12_7_0.LUT_INIT=16'b1110101011000000;
    LogicCell40 rTxByte_esr_0_LC_12_7_0 (
            .in0(N__6014),
            .in1(N__10342),
            .in2(N__5239),
            .in3(N__5230),
            .lcout(rTxByteZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12781),
            .ce(N__5718),
            .sr(N__11112));
    defparam rTxByte_esr_4_LC_12_7_1.C_ON=1'b0;
    defparam rTxByte_esr_4_LC_12_7_1.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_4_LC_12_7_1.LUT_INIT=16'b1110110010100000;
    LogicCell40 rTxByte_esr_4_LC_12_7_1 (
            .in0(N__10341),
            .in1(N__6015),
            .in2(N__5224),
            .in3(N__5347),
            .lcout(rTxByteZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12781),
            .ce(N__5718),
            .sr(N__11112));
    defparam rTxByte_esr_6_LC_12_7_2.C_ON=1'b0;
    defparam rTxByte_esr_6_LC_12_7_2.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_6_LC_12_7_2.LUT_INIT=16'b1111100010001000;
    LogicCell40 rTxByte_esr_6_LC_12_7_2 (
            .in0(N__6016),
            .in1(N__5206),
            .in2(N__5215),
            .in3(N__10343),
            .lcout(rTxByteZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12781),
            .ce(N__5718),
            .sr(N__11112));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIT6K22_6_LC_12_8_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIT6K22_6_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIT6K22_6_LC_12_8_1 .LUT_INIT=16'b1010000011011101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIT6K22_6_LC_12_8_1  (
            .in0(N__5869),
            .in1(N__5281),
            .in2(N__6523),
            .in3(N__5371),
            .lcout(\DUT.rFifoDatarx_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_12_8_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_12_8_3 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_12_8_3  (
            .in0(N__5955),
            .in1(N__5200),
            .in2(N__5885),
            .in3(N__5191),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI1BK22_7_LC_12_8_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI1BK22_7_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI1BK22_7_LC_12_8_4 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI1BK22_7_LC_12_8_4  (
            .in0(N__5275),
            .in1(N__6511),
            .in2(N__5194),
            .in3(N__5870),
            .lcout(\DUT.rFifoDatarx_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_12_8_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_12_8_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_12_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_12_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7022),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12777),
            .ce(N__6103),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNI0AQO1_LC_12_8_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNI0AQO1_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNI0AQO1_LC_12_8_6 .LUT_INIT=16'b1111111100110101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_0_RNI0AQO1_LC_12_8_6  (
            .in0(N__5316),
            .in1(N__5301),
            .in2(N__5956),
            .in3(N__5865),
            .lcout(\DUT.rFifoDataror_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_12_9_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_12_9_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_12_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7193),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12774),
            .ce(N__6502),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_12_9_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_12_9_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_12_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7245),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12774),
            .ce(N__6502),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_12_9_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_12_9_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_12_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8449),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12774),
            .ce(N__6502),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_12_9_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_12_9_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_12_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_12_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8510),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12774),
            .ce(N__6502),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_12_9_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_12_9_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_12_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7151),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12774),
            .ce(N__6502),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_12_9_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_12_9_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_12_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_12_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7106),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12774),
            .ce(N__6502),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_12_9_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_12_9_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_12_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_12_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7061),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12774),
            .ce(N__6502),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_12_9_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_12_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_12_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7023),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12774),
            .ce(N__6502),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rReadPtr_RNIDU4H2_0_LC_12_10_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rReadPtr_RNIDU4H2_0_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rReadPtr_RNIDU4H2_0_LC_12_10_0 .LUT_INIT=16'b0000111110001111;
    LogicCell40 \DUT.fifo_rx_inst.rReadPtr_RNIDU4H2_0_LC_12_10_0  (
            .in0(N__5853),
            .in1(N__5943),
            .in2(N__12440),
            .in3(N__5564),
            .lcout(\DUT.fifo_rx_inst.rReadPtr_RNIDU4H2Z0Z_0 ),
            .ltout(\DUT.fifo_rx_inst.rReadPtr_RNIDU4H2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rReadPtr_1_LC_12_10_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rReadPtr_1_LC_12_10_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rReadPtr_1_LC_12_10_1 .LUT_INIT=16'b0000100100001100;
    LogicCell40 \DUT.fifo_rx_inst.rReadPtr_1_LC_12_10_1  (
            .in0(N__5566),
            .in1(N__5854),
            .in2(N__5380),
            .in3(N__5949),
            .lcout(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12772),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_12_10_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_12_10_3 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_12_10_3  (
            .in0(N__5941),
            .in1(N__5377),
            .in2(N__5876),
            .in3(N__5323),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rReadPtr_0_LC_12_10_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rReadPtr_0_LC_12_10_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rReadPtr_0_LC_12_10_4 .LUT_INIT=16'b0010001000010001;
    LogicCell40 \DUT.fifo_rx_inst.rReadPtr_0_LC_12_10_4  (
            .in0(N__5948),
            .in1(N__5362),
            .in2(_gnd_net_),
            .in3(N__5565),
            .lcout(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12772),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNILUJ22_4_LC_12_10_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNILUJ22_4_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNILUJ22_4_LC_12_10_5 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNILUJ22_4_LC_12_10_5  (
            .in0(N__5398),
            .in1(N__5852),
            .in2(N__5356),
            .in3(N__5767),
            .lcout(\DUT.rFifoDatarx_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_12_10_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_12_10_6 .LUT_INIT=16'b0000001111110101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_12_10_6  (
            .in0(N__5329),
            .in1(N__6721),
            .in2(N__5879),
            .in3(N__5942),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIP2K22_5_LC_12_10_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIP2K22_5_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIP2K22_5_LC_12_10_7 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIP2K22_5_LC_12_10_7  (
            .in0(N__5338),
            .in1(N__6064),
            .in2(N__5332),
            .in3(N__5851),
            .lcout(\DUT.rFifoDatarx_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_12_11_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_12_11_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_12_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7113),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12770),
            .ce(N__6118),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_12_11_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_12_11_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_12_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7069),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12770),
            .ce(N__6118),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_12_12_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_12_12_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_12_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8514),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12769),
            .ce(N__6622),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_12_12_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_12_12_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_12_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7159),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12769),
            .ce(N__6622),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.wPllLocked_i_LC_12_30_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.wPllLocked_i_LC_12_30_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.wPllLocked_i_LC_12_30_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \DUT.uart_inst0.wPllLocked_i_LC_12_30_3  (
            .in0(N__12439),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(wPllLocked_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIHF7P_0_3_LC_13_1_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIHF7P_0_3_LC_13_1_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIHF7P_0_3_LC_13_1_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIHF7P_0_3_LC_13_1_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6640),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_i_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_2_0_LC_13_2_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_2_0_LC_13_2_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_2_0_LC_13_2_0 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_2_0_LC_13_2_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6328),
            .in3(N__6361),
            .lcout(\DUT.uart_inst0.rx_clk_divider_RNIP8N2B_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_0_0_LC_13_2_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_0_0_LC_13_2_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_0_0_LC_13_2_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_0_0_LC_13_2_1  (
            .in0(N__6358),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6316),
            .lcout(\DUT.uart_inst0.rx_clk_divider_RNIP8N2B_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_0_LC_13_2_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_0_LC_13_2_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_0_LC_13_2_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_0_LC_13_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6327),
            .in3(N__6360),
            .lcout(\DUT.uart_inst0.rx_clk_divider_RNIP8N2BZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNI8PF9A_0_LC_13_2_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI8PF9A_0_LC_13_2_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI8PF9A_0_LC_13_2_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNI8PF9A_0_LC_13_2_3  (
            .in0(N__8220),
            .in1(N__6163),
            .in2(N__8260),
            .in3(N__6150),
            .lcout(\DUT.uart_inst0.N_275 ),
            .ltout(\DUT.uart_inst0.N_275_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_0_c_RNO_LC_13_2_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_0_c_RNO_LC_13_2_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_0_c_RNO_LC_13_2_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_0_0_c_RNO_LC_13_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5383),
            .in3(N__6357),
            .lcout(\DUT.uart_inst0.rx_countdown_3_cry_0_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_1_0_LC_13_2_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_1_0_LC_13_2_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_1_0_LC_13_2_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIP8N2B_1_0_LC_13_2_5  (
            .in0(N__6359),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6317),
            .lcout(\DUT.uart_inst0.rx_clk_divider_RNIP8N2B_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_0_LC_13_3_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_0_LC_13_3_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_0_LC_13_3_0 .LUT_INIT=16'b1111110111011101;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_0_LC_13_3_0  (
            .in0(N__12421),
            .in1(N__5661),
            .in2(N__9856),
            .in3(N__8279),
            .lcout(\DUT.uart_inst0.g0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_2_LC_13_3_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_2_LC_13_3_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_2_LC_13_3_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_1_2_LC_13_3_1  (
            .in0(N__9640),
            .in1(N__9429),
            .in2(N__9504),
            .in3(N__9716),
            .lcout(),
            .ltout(\DUT.uart_inst0.g0_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_2_LC_13_3_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_2_LC_13_3_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_bits_remaining_2_LC_13_3_2 .LUT_INIT=16'b0101110011001100;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_2_LC_13_3_2  (
            .in0(N__8728),
            .in1(N__8702),
            .in2(N__5422),
            .in3(N__5404),
            .lcout(\DUT.uart_inst0.rx_bits_remainingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12814),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_1_6_LC_13_3_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_1_6_LC_13_3_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_1_6_LC_13_3_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_1_6_LC_13_3_3  (
            .in0(N__9639),
            .in1(N__9428),
            .in2(N__9503),
            .in3(N__9715),
            .lcout(),
            .ltout(\DUT.uart_inst0.g0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_6_LC_13_3_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_6_LC_13_3_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_6_LC_13_3_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \DUT.uart_inst0.recv_state_6_LC_13_3_4  (
            .in0(N__9560),
            .in1(N__9784),
            .in2(N__5419),
            .in3(N__8050),
            .lcout(\DUT.wRcvd ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12814),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_1_0_LC_13_3_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_1_0_LC_13_3_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_1_0_LC_13_3_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_1_0_LC_13_3_5  (
            .in0(_gnd_net_),
            .in1(N__6472),
            .in2(_gnd_net_),
            .in3(N__8032),
            .lcout(),
            .ltout(\DUT.uart_inst0.g3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_0_LC_13_3_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_0_LC_13_3_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_0_LC_13_3_6 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \DUT.uart_inst0.recv_state_0_LC_13_3_6  (
            .in0(N__9561),
            .in1(N__5416),
            .in2(N__5407),
            .in3(N__6169),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12814),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_2_LC_13_3_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_2_LC_13_3_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_2_LC_13_3_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_0_2_LC_13_3_7  (
            .in0(N__8308),
            .in1(N__9559),
            .in2(N__10626),
            .in3(N__8031),
            .lcout(\DUT.uart_inst0.g0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_13_4_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_13_4_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_13_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_13_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7290),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12808),
            .ce(N__10079),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNISS2R41_2_LC_13_4_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNISS2R41_2_LC_13_4_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNISS2R41_2_LC_13_4_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \DUT.uart_inst0.recv_state_RNISS2R41_2_LC_13_4_6  (
            .in0(N__8524),
            .in1(N__8027),
            .in2(N__9499),
            .in3(N__9416),
            .lcout(\DUT.uart_inst0.g0_8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rRxRead_esr_LC_13_5_1.C_ON=1'b0;
    defparam rRxRead_esr_LC_13_5_1.SEQ_MODE=4'b1000;
    defparam rRxRead_esr_LC_13_5_1.LUT_INIT=16'b1111111111101110;
    LogicCell40 rRxRead_esr_LC_13_5_1 (
            .in0(N__5624),
            .in1(N__10408),
            .in2(_gnd_net_),
            .in3(N__5590),
            .lcout(rRxReadZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12802),
            .ce(N__6253),
            .sr(N__11125));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIIL8L1_0_LC_13_5_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIIL8L1_0_LC_13_5_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIIL8L1_0_LC_13_5_6 .LUT_INIT=16'b0011001100110111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNIIL8L1_0_LC_13_5_6  (
            .in0(N__5589),
            .in1(N__10452),
            .in2(N__10413),
            .in3(N__5623),
            .lcout(\DUT.fifo_rx_inst.N_148 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_7_LC_13_6_0 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_7_LC_13_6_0 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_7_LC_13_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rRxData_esr_7_LC_13_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5530),
            .lcout(wRxFifoData_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12795),
            .ce(N__6450),
            .sr(N__11123));
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_1_LC_13_6_2 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_1_LC_13_6_2 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_1_LC_13_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rRxData_esr_1_LC_13_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5509),
            .lcout(wRxFifoData_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12795),
            .ce(N__6450),
            .sr(N__11123));
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_3_LC_13_6_3 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_3_LC_13_6_3 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_3_LC_13_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rRxData_esr_3_LC_13_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5494),
            .lcout(wRxFifoData_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12795),
            .ce(N__6450),
            .sr(N__11123));
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_5_LC_13_6_5 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_5_LC_13_6_5 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_5_LC_13_6_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \fifo_inst.ftdi_output_inst.rRxData_esr_5_LC_13_6_5  (
            .in0(N__5476),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(wRxFifoData_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12795),
            .ce(N__6450),
            .sr(N__11123));
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_2_LC_13_6_7 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_2_LC_13_6_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rRxData_esr_2_LC_13_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rRxData_esr_2_LC_13_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5461),
            .lcout(wRxFifoData_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12795),
            .ce(N__6450),
            .sr(N__11123));
    defparam rTxByte_esr_1_LC_13_7_1.C_ON=1'b0;
    defparam rTxByte_esr_1_LC_13_7_1.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_1_LC_13_7_1.LUT_INIT=16'b1110110010100000;
    LogicCell40 rTxByte_esr_1_LC_13_7_1 (
            .in0(N__10334),
            .in1(N__6009),
            .in2(N__5443),
            .in3(N__5683),
            .lcout(rTxByteZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12790),
            .ce(N__5719),
            .sr(N__11118));
    defparam rTxByte_esr_2_LC_13_7_2.C_ON=1'b0;
    defparam rTxByte_esr_2_LC_13_7_2.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_2_LC_13_7_2.LUT_INIT=16'b1110101011000000;
    LogicCell40 rTxByte_esr_2_LC_13_7_2 (
            .in0(N__6010),
            .in1(N__10336),
            .in2(N__5434),
            .in3(N__6034),
            .lcout(rTxByteZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12790),
            .ce(N__5719),
            .sr(N__11118));
    defparam rTxByte_esr_3_LC_13_7_4.C_ON=1'b0;
    defparam rTxByte_esr_3_LC_13_7_4.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_3_LC_13_7_4.LUT_INIT=16'b1110101011000000;
    LogicCell40 rTxByte_esr_3_LC_13_7_4 (
            .in0(N__6011),
            .in1(N__5761),
            .in2(N__10347),
            .in3(N__5965),
            .lcout(rTxByteZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12790),
            .ce(N__5719),
            .sr(N__11118));
    defparam rTxByte_esr_5_LC_13_7_5.C_ON=1'b0;
    defparam rTxByte_esr_5_LC_13_7_5.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_5_LC_13_7_5.LUT_INIT=16'b1110110010100000;
    LogicCell40 rTxByte_esr_5_LC_13_7_5 (
            .in0(N__10335),
            .in1(N__5755),
            .in2(N__5743),
            .in3(N__6012),
            .lcout(rTxByteZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12790),
            .ce(N__5719),
            .sr(N__11118));
    defparam rTxByte_esr_7_LC_13_7_7.C_ON=1'b0;
    defparam rTxByte_esr_7_LC_13_7_7.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_7_LC_13_7_7.LUT_INIT=16'b1110101011000000;
    LogicCell40 rTxByte_esr_7_LC_13_7_7 (
            .in0(N__5734),
            .in1(N__10340),
            .in2(N__5728),
            .in3(N__6013),
            .lcout(rTxByteZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12790),
            .ce(N__5719),
            .sr(N__11118));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1_1_LC_13_8_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1_1_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1_1_LC_13_8_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1_1_LC_13_8_0  (
            .in0(N__12424),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6500),
            .lcout(\DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1 ),
            .ltout(\DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_0_LC_13_8_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_0_LC_13_8_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rWritePtr_0_LC_13_8_1 .LUT_INIT=16'b0000101000000101;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_0_LC_13_8_1  (
            .in0(N__6777),
            .in1(_gnd_net_),
            .in2(N__5701),
            .in3(N__6806),
            .lcout(\DUT.fifo_rx_inst.rWritePtrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12784),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI9IJ22_1_LC_13_8_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI9IJ22_1_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI9IJ22_1_LC_13_8_2 .LUT_INIT=16'b1010000011001111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNI9IJ22_1_LC_13_8_2  (
            .in0(N__6529),
            .in1(N__5698),
            .in2(N__5887),
            .in3(N__5692),
            .lcout(\DUT.rFifoDatarx_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_2_1_LC_13_8_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_2_1_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_2_1_LC_13_8_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI96D91_2_1_LC_13_8_3  (
            .in0(N__6741),
            .in1(N__5670),
            .in2(N__6783),
            .in3(N__5635),
            .lcout(\DUT.fifo_rx_inst.rFifoData_awe3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_1_LC_13_8_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_1_LC_13_8_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rWritePtr_1_LC_13_8_4 .LUT_INIT=16'b0000000011000110;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_1_LC_13_8_4  (
            .in0(N__6782),
            .in1(N__6743),
            .in2(N__6811),
            .in3(N__5677),
            .lcout(\DUT.fifo_rx_inst.rWritePtrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12784),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_13_8_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_13_8_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_13_8_5  (
            .in0(_gnd_net_),
            .in1(N__5671),
            .in2(_gnd_net_),
            .in3(N__5634),
            .lcout(\DUT.fifo_rx_inst.N_194 ),
            .ltout(\DUT.fifo_rx_inst.N_194_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_13_8_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_13_8_6 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_13_8_6  (
            .in0(_gnd_net_),
            .in1(N__6776),
            .in2(N__6055),
            .in3(N__6742),
            .lcout(\DUT.fifo_rx_inst.rFifoData_awe0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_13_9_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_13_9_2 .LUT_INIT=16'b0000010111110011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_13_9_2  (
            .in0(N__6052),
            .in1(N__6139),
            .in2(N__5881),
            .in3(N__5947),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIDMJ22_2_LC_13_9_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIDMJ22_2_LC_13_9_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIDMJ22_2_LC_13_9_3 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIDMJ22_2_LC_13_9_3  (
            .in0(N__6043),
            .in1(N__6073),
            .in2(N__6037),
            .in3(N__5861),
            .lcout(\DUT.rFifoDatarx_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_13_9_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_13_9_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_13_9_4  (
            .in0(N__6802),
            .in1(N__6778),
            .in2(_gnd_net_),
            .in3(N__6744),
            .lcout(\DUT.fifo_rx_inst.rFifoData_awe2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_13_9_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_13_9_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_13_9_5 .LUT_INIT=16'b0001111110111111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_13_9_5  (
            .in0(N__5946),
            .in1(N__6570),
            .in2(N__5880),
            .in3(N__6483),
            .lcout(),
            .ltout(\DUT.rFifoDataror_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rTxByte_6_0_a2_0_LC_13_9_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rTxByte_6_0_a2_0_LC_13_9_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rTxByte_6_0_a2_0_LC_13_9_6 .LUT_INIT=16'b0000010101010101;
    LogicCell40 \DUT.uart_inst0.rTxByte_6_0_a2_0_LC_13_9_6  (
            .in0(N__10333),
            .in1(_gnd_net_),
            .in2(N__6025),
            .in3(N__6022),
            .lcout(\DUT.uart_inst0.N_257 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_13_10_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_13_10_0 .LUT_INIT=16'b0101000101011011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_13_10_0  (
            .in0(N__5945),
            .in1(N__6130),
            .in2(N__5878),
            .in3(N__6709),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIHQJ22_3_LC_13_10_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIHQJ22_3_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIHQJ22_3_LC_13_10_1 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__RNIHQJ22_3_LC_13_10_1  (
            .in0(N__5983),
            .in1(N__5977),
            .in2(N__5968),
            .in3(N__5847),
            .lcout(\DUT.rFifoDatarx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_13_10_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_13_10_6 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_13_10_6  (
            .in0(N__5944),
            .in1(N__6703),
            .in2(N__5877),
            .in3(N__6124),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_13_11_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_13_11_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_13_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8459),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12773),
            .ce(N__6114),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_13_11_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_13_11_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_13_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8515),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12773),
            .ce(N__6114),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_13_11_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_13_11_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_13_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_13_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7158),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12773),
            .ce(N__6114),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_13_12_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_13_12_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_13_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_13_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8460),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12771),
            .ce(N__6613),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_13_12_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_13_12_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_13_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7114),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12771),
            .ce(N__6613),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_3_LC_14_1_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_3_LC_14_1_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_3_LC_14_1_0 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_3_LC_14_1_0  (
            .in0(N__6639),
            .in1(N__9349),
            .in2(_gnd_net_),
            .in3(N__6326),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12826),
            .ce(N__12340),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_15_LC_14_1_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_15_LC_14_1_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_15_LC_14_1_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_15_LC_14_1_1  (
            .in0(_gnd_net_),
            .in1(N__9352),
            .in2(_gnd_net_),
            .in3(N__6937),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12826),
            .ce(N__12340),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_0_LC_14_1_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_0_LC_14_1_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_0_LC_14_1_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_0_LC_14_1_2  (
            .in0(N__9351),
            .in1(N__9771),
            .in2(_gnd_net_),
            .in3(N__9575),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12826),
            .ce(N__12340),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_LC_14_1_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_LC_14_1_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_3_LC_14_1_3 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_LC_14_1_3  (
            .in0(N__9772),
            .in1(N__9354),
            .in2(_gnd_net_),
            .in3(N__9435),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12826),
            .ce(N__12340),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_4_LC_14_1_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_4_LC_14_1_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_4_LC_14_1_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_4_LC_14_1_4  (
            .in0(_gnd_net_),
            .in1(N__9348),
            .in2(_gnd_net_),
            .in3(N__6901),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12826),
            .ce(N__12340),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_7_LC_14_1_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_7_LC_14_1_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_7_LC_14_1_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_7_LC_14_1_5  (
            .in0(_gnd_net_),
            .in1(N__8095),
            .in2(_gnd_net_),
            .in3(N__9353),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12826),
            .ce(N__12340),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_6_LC_14_1_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_6_LC_14_1_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_6_LC_14_1_6 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_6_LC_14_1_6  (
            .in0(N__9350),
            .in1(N__6244),
            .in2(_gnd_net_),
            .in3(N__6854),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12826),
            .ce(N__12340),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_LC_14_1_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_LC_14_1_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_out_LC_14_1_7 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \DUT.uart_inst0.tx_out_LC_14_1_7  (
            .in0(N__11441),
            .in1(N__10867),
            .in2(N__9046),
            .in3(N__8764),
            .lcout(P1A7_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12826),
            .ce(N__12340),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIQ3QE2_14_LC_14_2_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIQ3QE2_14_LC_14_2_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIQ3QE2_14_LC_14_2_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIQ3QE2_14_LC_14_2_0  (
            .in0(N__6875),
            .in1(N__8195),
            .in2(N__6855),
            .in3(N__8234),
            .lcout(\DUT.uart_inst0.rx_clk_divider_5_i_a2_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_14_LC_14_2_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_14_LC_14_2_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_14_LC_14_2_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_14_LC_14_2_1  (
            .in0(N__8196),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9363),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12822),
            .ce(N__12344),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_5_LC_14_2_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_5_LC_14_2_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_5_LC_14_2_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNO_0_5_LC_14_2_2  (
            .in0(N__6368),
            .in1(N__8182),
            .in2(N__6856),
            .in3(N__6151),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_222_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_5_LC_14_2_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_5_LC_14_2_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_5_LC_14_2_3 .LUT_INIT=16'b1111111111110011;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_5_LC_14_2_3  (
            .in0(_gnd_net_),
            .in1(N__9362),
            .in2(N__6157),
            .in3(N__6877),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12822),
            .ce(N__12344),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNI2VEI1_2_LC_14_2_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI2VEI1_2_LC_14_2_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI2VEI1_2_LC_14_2_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNI2VEI1_2_LC_14_2_4  (
            .in0(_gnd_net_),
            .in1(N__7968),
            .in2(_gnd_net_),
            .in3(N__6900),
            .lcout(),
            .ltout(\DUT.uart_inst0.rx_clk_divider_5_i_a2_11_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIQEH13_10_LC_14_2_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIQEH13_10_LC_14_2_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIQEH13_10_LC_14_2_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIQEH13_10_LC_14_2_5  (
            .in0(N__8343),
            .in1(N__6936),
            .in2(N__6154),
            .in3(N__8361),
            .lcout(\DUT.uart_inst0.rx_clk_divider_5_i_a2_11_5 ),
            .ltout(\DUT.uart_inst0.rx_clk_divider_5_i_a2_11_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_6_LC_14_2_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_6_LC_14_2_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNO_0_6_LC_14_2_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNO_0_6_LC_14_2_6  (
            .in0(N__6876),
            .in1(N__8181),
            .in2(N__6247),
            .in3(N__6367),
            .lcout(\DUT.uart_inst0.N_221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_16_LC_14_2_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_16_LC_14_2_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_16_LC_14_2_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_16_LC_14_2_7  (
            .in0(N__8235),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9364),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12822),
            .ce(N__12344),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_0_c_LC_14_3_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_0_c_LC_14_3_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_0_c_LC_14_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_0_0_c_LC_14_3_0  (
            .in0(_gnd_net_),
            .in1(N__6387),
            .in2(N__6238),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_3_0_),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_0_c_RNIPQVSB_LC_14_3_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_0_c_RNIPQVSB_LC_14_3_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_0_c_RNIPQVSB_LC_14_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_0_0_c_RNIPQVSB_LC_14_3_1  (
            .in0(_gnd_net_),
            .in1(N__7984),
            .in2(N__6229),
            .in3(N__6220),
            .lcout(\DUT.uart_inst0.rx_countdown_3_1 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_countdown_3_cry_0 ),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_0_c_RNIRV51C_LC_14_3_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_0_c_RNIRV51C_LC_14_3_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_0_c_RNIRV51C_LC_14_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_1_0_c_RNIRV51C_LC_14_3_2  (
            .in0(_gnd_net_),
            .in1(N__8374),
            .in2(N__6217),
            .in3(N__6208),
            .lcout(\DUT.uart_inst0.rx_countdown_3_2 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_countdown_3_cry_1 ),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_2_0_c_RNIT4CLB_LC_14_3_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_2_0_c_RNIT4CLB_LC_14_3_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_2_0_c_RNIT4CLB_LC_14_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_2_0_c_RNIT4CLB_LC_14_3_3  (
            .in0(_gnd_net_),
            .in1(N__6205),
            .in2(N__6196),
            .in3(N__6187),
            .lcout(\DUT.uart_inst0.rx_countdown_3_3 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_countdown_3_cry_2 ),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_0_c_RNIV9IPB_LC_14_3_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_0_c_RNIV9IPB_LC_14_3_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_0_c_RNIV9IPB_LC_14_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_3_0_c_RNIV9IPB_LC_14_3_4  (
            .in0(_gnd_net_),
            .in1(N__6184),
            .in2(N__9664),
            .in3(N__6178),
            .lcout(\DUT.uart_inst0.rx_countdown_3_4 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_countdown_3_cry_3 ),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_4_0_c_RNI1FOTB_LC_14_3_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_4_0_c_RNI1FOTB_LC_14_3_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_4_0_c_RNI1FOTB_LC_14_3_5 .LUT_INIT=16'b1001010101101010;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_4_0_c_RNI1FOTB_LC_14_3_5  (
            .in0(N__8062),
            .in1(N__6324),
            .in2(N__6375),
            .in3(N__6175),
            .lcout(\DUT.uart_inst0.rx_countdown_3_5 ),
            .ltout(\DUT.uart_inst0.rx_countdown_3_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_2_0_LC_14_3_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_2_0_LC_14_3_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_2_0_LC_14_3_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_2_0_LC_14_3_6  (
            .in0(N__9486),
            .in1(N__9421),
            .in2(N__6172),
            .in3(N__9714),
            .lcout(\DUT.uart_inst0.g3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNITI4IB_0_LC_14_3_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNITI4IB_0_LC_14_3_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNITI4IB_0_LC_14_3_7 .LUT_INIT=16'b0101101010101010;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNITI4IB_0_LC_14_3_7  (
            .in0(N__6388),
            .in1(_gnd_net_),
            .in2(N__6376),
            .in3(N__6325),
            .lcout(\DUT.uart_inst0.rx_countdown_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_3_LC_14_4_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_3_LC_14_4_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_3_LC_14_4_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_0_3_LC_14_4_2  (
            .in0(N__8662),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8605),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_196_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_3_LC_14_4_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_3_LC_14_4_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_bits_remaining_3_LC_14_4_3 .LUT_INIT=16'b1110111011101011;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_3_LC_14_4_3  (
            .in0(N__9237),
            .in1(N__8631),
            .in2(N__6292),
            .in3(N__8701),
            .lcout(\DUT.uart_inst0.rx_bits_remainingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12815),
            .ce(N__6286),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_1_LC_14_4_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_1_LC_14_4_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_1_1_LC_14_4_4 .LUT_INIT=16'b1111111101100110;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_1_1_LC_14_4_4  (
            .in0(N__8660),
            .in1(N__8604),
            .in2(_gnd_net_),
            .in3(N__9235),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_33_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_1_LC_14_4_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_1_LC_14_4_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_0_1_LC_14_4_5 .LUT_INIT=16'b0000000001000001;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_0_1_LC_14_4_5  (
            .in0(N__9712),
            .in1(N__8661),
            .in2(N__6289),
            .in3(N__9627),
            .lcout(\DUT.uart_inst0.rx_bits_remaining_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_0_c_RNIP8I482_LC_14_4_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_0_c_RNIP8I482_LC_14_4_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_0_c_RNIP8I482_LC_14_4_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_3_0_c_RNIP8I482_LC_14_4_6  (
            .in0(N__9626),
            .in1(N__9552),
            .in2(N__6268),
            .in3(N__9713),
            .lcout(\DUT.uart_inst0.rx_countdown_3_cry_3_0_c_RNIP8IZ0Z482 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_0_LC_14_4_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_0_LC_14_4_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_bits_remaining_0_LC_14_4_7 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_0_LC_14_4_7  (
            .in0(N__9236),
            .in1(_gnd_net_),
            .in2(N__8613),
            .in3(_gnd_net_),
            .lcout(\DUT.uart_inst0.rx_bits_remainingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12815),
            .ce(N__6286),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_1_LC_14_5_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_1_LC_14_5_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_bits_remaining_1_LC_14_5_1 .LUT_INIT=16'b1011010011110000;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_1_LC_14_5_1  (
            .in0(N__9576),
            .in1(N__6274),
            .in2(N__8672),
            .in3(N__6267),
            .lcout(\DUT.uart_inst0.rx_bits_remainingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12809),
            .ce(),
            .sr(_gnd_net_));
    defparam rRxRead_esr_RNO_LC_14_5_2.C_ON=1'b0;
    defparam rRxRead_esr_RNO_LC_14_5_2.SEQ_MODE=4'b0000;
    defparam rRxRead_esr_RNO_LC_14_5_2.LUT_INIT=16'b1111111101010101;
    LogicCell40 rRxRead_esr_RNO_LC_14_5_2 (
            .in0(N__10321),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11148),
            .lcout(P1A2_c_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_4_LC_14_5_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_4_LC_14_5_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_4_LC_14_5_6 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \DUT.uart_inst0.recv_state_4_LC_14_5_6  (
            .in0(N__6468),
            .in1(N__9759),
            .in2(N__10640),
            .in3(N__7252),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12809),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIDTQ4_1_LC_14_5_7 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIDTQ4_1_LC_14_5_7 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIDTQ4_1_LC_14_5_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_RNIDTQ4_1_LC_14_5_7  (
            .in0(N__11147),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10369),
            .lcout(\fifo_inst.ftdi_output_inst.rFifoState_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_14_6_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_14_6_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_14_6_0 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_14_6_0  (
            .in0(N__6400),
            .in1(N__11674),
            .in2(N__6421),
            .in3(N__11536),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_14_6_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_14_6_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_14_6_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_14_6_1  (
            .in0(N__11675),
            .in1(N__6433),
            .in2(N__6424),
            .in3(N__7336),
            .lcout(\DUT.rFifoDatarx_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_14_6_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_14_6_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_14_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_14_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7371),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12803),
            .ce(N__10078),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_14_6_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_14_6_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_14_6_3 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_14_6_3  (
            .in0(N__11535),
            .in1(N__6394),
            .in2(N__11680),
            .in3(N__6412),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_14_7_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_14_7_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_14_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_14_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7360),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12796),
            .ce(N__6559),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_14_7_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_14_7_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_14_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_14_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7312),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12796),
            .ce(N__6559),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_14_7_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_14_7_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_14_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_14_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10141),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12796),
            .ce(N__6559),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_14_7_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_14_7_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_14_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_14_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7279),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12796),
            .ce(N__6559),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_14_7_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_14_7_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_14_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_14_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7516),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12796),
            .ce(N__6559),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_14_7_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_14_7_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_14_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_14_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7438),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12796),
            .ce(N__6559),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_14_7_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_14_7_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_14_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_14_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7583),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12796),
            .ce(N__6559),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_14_7_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_14_7_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_14_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_14_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10102),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12796),
            .ce(N__6559),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_14_8_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_14_8_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_14_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7237),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12791),
            .ce(N__6617),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_14_8_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_14_8_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_14_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_14_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7051),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12791),
            .ce(N__6617),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_14_8_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_14_8_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_14_8_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_14_8_7  (
            .in0(N__7012),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12791),
            .ce(N__6617),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_3_LC_14_9_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_3_LC_14_9_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_3_LC_14_9_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_3_LC_14_9_0  (
            .in0(_gnd_net_),
            .in1(N__6484),
            .in2(_gnd_net_),
            .in3(N__6501),
            .lcout(\DUT.fifo_rx_inst.rFifoDataro_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12785),
            .ce(),
            .sr(N__11113));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_LC_14_9_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_LC_14_9_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_LC_14_9_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_0_LC_14_9_2  (
            .in0(_gnd_net_),
            .in1(N__7717),
            .in2(_gnd_net_),
            .in3(N__10027),
            .lcout(\DUT.fifo_tx_inst.rFifoDataro_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12785),
            .ce(),
            .sr(N__11113));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_1_LC_14_9_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_1_LC_14_9_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_1_LC_14_9_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_1_LC_14_9_3  (
            .in0(_gnd_net_),
            .in1(N__7704),
            .in2(_gnd_net_),
            .in3(N__6552),
            .lcout(\DUT.fifo_tx_inst.rFifoDataro_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12785),
            .ce(),
            .sr(N__11113));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_3_LC_14_9_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_3_LC_14_9_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_3_LC_14_9_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_3_LC_14_9_5  (
            .in0(_gnd_net_),
            .in1(N__7393),
            .in2(_gnd_net_),
            .in3(N__7729),
            .lcout(\DUT.fifo_tx_inst.rFifoDataro_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12785),
            .ce(),
            .sr(N__11113));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_LC_14_9_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_LC_14_9_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_LC_14_9_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_2_LC_14_9_6  (
            .in0(_gnd_net_),
            .in1(N__6571),
            .in2(_gnd_net_),
            .in3(N__6594),
            .lcout(\DUT.fifo_rx_inst.rFifoDataro_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12785),
            .ce(),
            .sr(N__11113));
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_0_1_LC_14_10_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_0_1_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_0_1_LC_14_10_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_0_1_LC_14_10_1  (
            .in0(N__7646),
            .in1(N__7612),
            .in2(_gnd_net_),
            .in3(N__8982),
            .lcout(\DUT.fifo_tx_inst.rFifoData_awe1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_1_1_LC_14_10_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_1_1_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_1_1_LC_14_10_2 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_1_1_LC_14_10_2  (
            .in0(N__8983),
            .in1(_gnd_net_),
            .in2(N__7618),
            .in3(N__7647),
            .lcout(\DUT.fifo_tx_inst.rFifoData_awe0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_1_LC_14_10_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_1_LC_14_10_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rWritePtr_1_LC_14_10_3 .LUT_INIT=16'b0010001000010010;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_1_LC_14_10_3  (
            .in0(N__7617),
            .in1(N__6538),
            .in2(N__7654),
            .in3(N__8985),
            .lcout(\DUT.fifo_tx_inst.rWritePtrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12779),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNI8BKM_2_LC_14_10_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNI8BKM_2_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNI8BKM_2_LC_14_10_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNI8BKM_2_LC_14_10_4  (
            .in0(N__7611),
            .in1(N__10222),
            .in2(N__7653),
            .in3(N__9919),
            .lcout(\DUT.fifo_tx_inst.rFifoData_awe3 ),
            .ltout(\DUT.fifo_tx_inst.rFifoData_awe3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNI4PUO_2_LC_14_10_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNI4PUO_2_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNI4PUO_2_LC_14_10_5 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNI4PUO_2_LC_14_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6541),
            .in3(N__12428),
            .lcout(\DUT.fifo_tx_inst.un1_i11_i ),
            .ltout(\DUT.fifo_tx_inst.un1_i11_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_0_LC_14_10_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_0_LC_14_10_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rWritePtr_0_LC_14_10_6 .LUT_INIT=16'b0000101000000101;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_0_LC_14_10_6  (
            .in0(N__8984),
            .in1(_gnd_net_),
            .in2(N__6532),
            .in3(N__7648),
            .lcout(\DUT.fifo_tx_inst.rWritePtrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12779),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_14_10_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_14_10_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_14_10_7  (
            .in0(N__6810),
            .in1(N__6784),
            .in2(_gnd_net_),
            .in3(N__6748),
            .lcout(\DUT.fifo_rx_inst.rFifoData_awe1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_14_11_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_14_11_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_14_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_14_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7105),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12776),
            .ce(N__6682),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_14_11_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_14_11_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_14_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_14_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8506),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12776),
            .ce(N__6682),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_14_11_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_14_11_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_14_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_14_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7150),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12776),
            .ce(N__6682),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_14_23_2.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_14_23_2.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_14_23_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_14_23_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_15_1_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_15_1_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_15_1_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_15_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8115),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_15_1_0_),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNID95P_1_LC_15_1_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_RNID95P_1_LC_15_1_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNID95P_1_LC_15_1_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNID95P_1_LC_15_1_1  (
            .in0(_gnd_net_),
            .in1(N__12944),
            .in2(N__8071),
            .in3(N__6655),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_1 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_0 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIFC6P_2_LC_15_1_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIFC6P_2_LC_15_1_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIFC6P_2_LC_15_1_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIFC6P_2_LC_15_1_2  (
            .in0(_gnd_net_),
            .in1(N__12953),
            .in2(N__7957),
            .in3(N__6652),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_2 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_1 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIHF7P_3_LC_15_1_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIHF7P_3_LC_15_1_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIHF7P_3_LC_15_1_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIHF7P_3_LC_15_1_3  (
            .in0(_gnd_net_),
            .in1(N__12945),
            .in2(N__6649),
            .in3(N__6625),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_3 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_2 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIJI8P_4_LC_15_1_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIJI8P_4_LC_15_1_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIJI8P_4_LC_15_1_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIJI8P_4_LC_15_1_4  (
            .in0(_gnd_net_),
            .in1(N__6907),
            .in2(N__12996),
            .in3(N__6889),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_4 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_3 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNILL9P_5_LC_15_1_5 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_RNILL9P_5_LC_15_1_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNILL9P_5_LC_15_1_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNILL9P_5_LC_15_1_5  (
            .in0(_gnd_net_),
            .in1(N__12949),
            .in2(N__6886),
            .in3(N__6865),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_5 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_4 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNINOAP_6_LC_15_1_6 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_RNINOAP_6_LC_15_1_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNINOAP_6_LC_15_1_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNINOAP_6_LC_15_1_6  (
            .in0(_gnd_net_),
            .in1(N__6862),
            .in2(N__12997),
            .in3(N__6835),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_6 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_5 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIPRBP_7_LC_15_1_7 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIPRBP_7_LC_15_1_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIPRBP_7_LC_15_1_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIPRBP_7_LC_15_1_7  (
            .in0(_gnd_net_),
            .in1(N__6832),
            .in2(N__12998),
            .in3(N__6826),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_7 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_6 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIRUCP_8_LC_15_2_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIRUCP_8_LC_15_2_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIRUCP_8_LC_15_2_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIRUCP_8_LC_15_2_0  (
            .in0(_gnd_net_),
            .in1(N__7759),
            .in2(N__13078),
            .in3(N__6823),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_8 ),
            .ltout(),
            .carryin(bfn_15_2_0_),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIT1EP_9_LC_15_2_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIT1EP_9_LC_15_2_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIT1EP_9_LC_15_2_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIT1EP_9_LC_15_2_1  (
            .in0(_gnd_net_),
            .in1(N__8152),
            .in2(N__13075),
            .in3(N__6820),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_9 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_8 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNI6KQI_10_LC_15_2_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI6KQI_10_LC_15_2_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI6KQI_10_LC_15_2_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNI6KQI_10_LC_15_2_2  (
            .in0(_gnd_net_),
            .in1(N__8332),
            .in2(N__13076),
            .in3(N__6817),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_10 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_9 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIFEUD_11_LC_15_2_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIFEUD_11_LC_15_2_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIFEUD_11_LC_15_2_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIFEUD_11_LC_15_2_3  (
            .in0(_gnd_net_),
            .in1(N__8137),
            .in2(N__13072),
            .in3(N__6814),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_11 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_10 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIHHVD_12_LC_15_2_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIHHVD_12_LC_15_2_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIHHVD_12_LC_15_2_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIHHVD_12_LC_15_2_4  (
            .in0(_gnd_net_),
            .in1(N__8122),
            .in2(N__13077),
            .in3(N__6961),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_12 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_11 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIJK0E_13_LC_15_2_5 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIJK0E_13_LC_15_2_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIJK0E_13_LC_15_2_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIJK0E_13_LC_15_2_5  (
            .in0(_gnd_net_),
            .in1(N__8314),
            .in2(N__13073),
            .in3(N__6958),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_13 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_12 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNILN1E_14_LC_15_2_6 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_RNILN1E_14_LC_15_2_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNILN1E_14_LC_15_2_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNILN1E_14_LC_15_2_6  (
            .in0(_gnd_net_),
            .in1(N__13055),
            .in2(N__6955),
            .in3(N__6946),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_14 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_13 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNINQ2E_15_LC_15_2_7 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_RNINQ2E_15_LC_15_2_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNINQ2E_15_LC_15_2_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNINQ2E_15_LC_15_2_7  (
            .in0(_gnd_net_),
            .in1(N__6943),
            .in2(N__13074),
            .in3(N__6925),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_15 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_14 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIPT3E_16_LC_15_3_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIPT3E_16_LC_15_3_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIPT3E_16_LC_15_3_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIPT3E_16_LC_15_3_0  (
            .in0(_gnd_net_),
            .in1(N__6922),
            .in2(N__13071),
            .in3(N__6916),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_16 ),
            .ltout(),
            .carryin(bfn_15_3_0_),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIR05E_17_LC_15_3_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIR05E_17_LC_15_3_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIR05E_17_LC_15_3_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIR05E_17_LC_15_3_1  (
            .in0(_gnd_net_),
            .in1(N__8350),
            .in2(_gnd_net_),
            .in3(N__6913),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_15_3_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_15_3_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_15_3_2 .LUT_INIT=16'b0100010101000100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_15_3_2  (
            .in0(N__8026),
            .in1(N__8556),
            .in2(N__9869),
            .in3(N__9241),
            .lcout(\DUT.uart_inst0.g0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_2_4_LC_15_3_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_2_4_LC_15_3_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_2_4_LC_15_3_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_2_4_LC_15_3_3  (
            .in0(N__9746),
            .in1(N__8022),
            .in2(N__9430),
            .in3(N__9705),
            .lcout(),
            .ltout(\DUT.uart_inst0.recv_state_RNO_2Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_1_4_LC_15_3_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_1_4_LC_15_3_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_1_4_LC_15_3_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_1_4_LC_15_3_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6910),
            .in3(N__9625),
            .lcout(\DUT.uart_inst0.G_11_i_a4_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_2_2_LC_15_3_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_2_2_LC_15_3_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_2_2_LC_15_3_5 .LUT_INIT=16'b0100010100000000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_2_2_LC_15_3_5  (
            .in0(N__9747),
            .in1(N__9860),
            .in2(N__8284),
            .in3(N__9487),
            .lcout(\DUT.uart_inst0.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNI1K9CC_2_LC_15_3_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNI1K9CC_2_LC_15_3_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNI1K9CC_2_LC_15_3_6 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNI1K9CC_2_LC_15_3_6  (
            .in0(_gnd_net_),
            .in1(N__10638),
            .in2(N__8039),
            .in3(N__8555),
            .lcout(\DUT.uart_inst0.rx_bits_remaining_2_sqmuxa_0_a2_0_a2_0_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_15_3_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_15_3_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_15_3_7 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_15_3_7  (
            .in0(N__9551),
            .in1(_gnd_net_),
            .in2(N__9431),
            .in3(N__9706),
            .lcout(\DUT.uart_inst0.g0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNIM4BC72_2_LC_15_4_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNIM4BC72_2_LC_15_4_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNIM4BC72_2_LC_15_4_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \DUT.uart_inst0.recv_state_RNIM4BC72_2_LC_15_4_0  (
            .in0(N__9628),
            .in1(N__6982),
            .in2(N__9571),
            .in3(N__6972),
            .lcout(\DUT.uart_inst0.rx_bits_remaining_2_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_5_LC_15_4_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_5_LC_15_4_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_5_LC_15_4_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_5_LC_15_4_1  (
            .in0(N__8030),
            .in1(N__9556),
            .in2(_gnd_net_),
            .in3(N__9630),
            .lcout(),
            .ltout(\DUT.uart_inst0.rx_countdown_8_i_0_o2_1_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_5_LC_15_4_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_5_LC_15_4_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_5_LC_15_4_2 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \DUT.uart_inst0.recv_state_5_LC_15_4_2  (
            .in0(N__8719),
            .in1(N__10633),
            .in2(N__6976),
            .in3(N__6973),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12818),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_0_c_RNINE4G31_LC_15_4_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_0_c_RNINE4G31_LC_15_4_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_0_c_RNINE4G31_LC_15_4_3 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_1_0_c_RNINE4G31_LC_15_4_3  (
            .in0(_gnd_net_),
            .in1(N__9417),
            .in2(N__9497),
            .in3(N__9707),
            .lcout(\DUT.uart_inst0.recv_state_ns_0_i_0_0_o2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_0_c_RNIHVHJ31_LC_15_4_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_0_c_RNIHVHJ31_LC_15_4_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_0_c_RNIHVHJ31_LC_15_4_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_1_0_c_RNIHVHJ31_LC_15_4_4  (
            .in0(N__9419),
            .in1(N__9479),
            .in2(_gnd_net_),
            .in3(N__8029),
            .lcout(),
            .ltout(\DUT.uart_inst0.G_9_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_0_c_RNIEB1T62_LC_15_4_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_0_c_RNIEB1T62_LC_15_4_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_0_c_RNIEB1T62_LC_15_4_5 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_3_0_c_RNIEB1T62_LC_15_4_5  (
            .in0(N__9558),
            .in1(N__9629),
            .in2(N__6964),
            .in3(N__9711),
            .lcout(\DUT.uart_inst0.N_193 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_2_1_LC_15_4_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_2_1_LC_15_4_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_2_1_LC_15_4_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_2_1_LC_15_4_6  (
            .in0(N__9418),
            .in1(N__9316),
            .in2(N__9720),
            .in3(N__8028),
            .lcout(\DUT.uart_inst0.recv_state_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_4_LC_15_4_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_4_LC_15_4_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_4_LC_15_4_7 .LUT_INIT=16'b0100010100000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_4_LC_15_4_7  (
            .in0(N__9557),
            .in1(N__9420),
            .in2(N__9498),
            .in3(N__7258),
            .lcout(\DUT.uart_inst0.N_4_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_1_LC_15_5_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_1_LC_15_5_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_1_LC_15_5_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.uart_inst0.rx_data_1_LC_15_5_1  (
            .in0(N__8430),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.wRxByte_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12816),
            .ce(N__8418),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_0_LC_15_5_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_0_LC_15_5_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_0_LC_15_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_0_LC_15_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7214),
            .lcout(\DUT.wRxByte_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12816),
            .ce(N__8418),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_3_LC_15_5_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_3_LC_15_5_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_3_LC_15_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_3_LC_15_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7130),
            .lcout(\DUT.wRxByte_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12816),
            .ce(N__8418),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_4_LC_15_5_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_4_LC_15_5_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_4_LC_15_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_4_LC_15_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7085),
            .lcout(\DUT.wRxByte_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12816),
            .ce(N__8418),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_5_LC_15_5_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_5_LC_15_5_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_5_LC_15_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_5_LC_15_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7040),
            .lcout(\DUT.wRxByte_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12816),
            .ce(N__8418),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_6_LC_15_5_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_6_LC_15_5_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_6_LC_15_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_6_LC_15_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7000),
            .lcout(\DUT.wRxByte_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12816),
            .ce(N__8418),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_7_LC_15_5_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_7_LC_15_5_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_7_LC_15_5_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.uart_inst0.rx_data_7_LC_15_5_7  (
            .in0(N__9855),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.wRxByte_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12816),
            .ce(N__8418),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_15_6_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_15_6_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_15_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_15_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7329),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12810),
            .ce(N__7413),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_15_6_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_15_6_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_15_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_15_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10158),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12810),
            .ce(N__7413),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_15_6_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_15_6_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_15_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_15_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7294),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12810),
            .ce(N__7413),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_15_6_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_15_6_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_15_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_15_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7528),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12810),
            .ce(N__7413),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_15_6_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_15_6_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_15_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_15_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7456),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12810),
            .ce(N__7413),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_15_6_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_15_6_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_15_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_15_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10120),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12810),
            .ce(N__7413),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_15_7_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_15_7_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_15_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_15_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7370),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12804),
            .ce(N__7948),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_15_7_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_15_7_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_15_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_15_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7322),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12804),
            .ce(N__7948),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_15_7_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_15_7_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_15_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_15_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10151),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12804),
            .ce(N__7948),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_15_7_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_15_7_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_15_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_15_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7289),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12804),
            .ce(N__7948),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_15_7_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_15_7_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_15_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_15_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7526),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12804),
            .ce(N__7948),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_15_7_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_15_7_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_15_7_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_15_7_5  (
            .in0(N__7448),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12804),
            .ce(N__7948),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_15_7_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_15_7_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_15_7_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_15_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7590),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12804),
            .ce(N__7948),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_15_7_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_15_7_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_15_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_15_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10112),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12804),
            .ce(N__7948),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_15_8_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_15_8_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_15_8_0 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_15_8_0  (
            .in0(N__11540),
            .in1(N__7555),
            .in2(N__7492),
            .in3(N__11661),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_15_8_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_15_8_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_15_8_1  (
            .in0(N__11666),
            .in1(N__7549),
            .in2(N__7540),
            .in3(N__7537),
            .lcout(\DUT.rFifoDatarx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_15_8_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_15_8_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_15_8_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_15_8_2  (
            .in0(N__7527),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12797),
            .ce(N__10061),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_15_8_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_15_8_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_15_8_3 .LUT_INIT=16'b0000010111110011;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_15_8_3  (
            .in0(N__7483),
            .in1(N__7420),
            .in2(N__11678),
            .in3(N__11541),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_15_8_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_15_8_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_15_8_4 .LUT_INIT=16'b1010110000001111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_15_8_4  (
            .in0(N__7477),
            .in1(N__7468),
            .in2(N__7459),
            .in3(N__11665),
            .lcout(\DUT.rFifoDatarx_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_15_8_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_15_8_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_15_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_15_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7455),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12797),
            .ce(N__10061),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_15_8_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_15_8_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_15_8_6 .LUT_INIT=16'b0101010100100111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_15_8_6  (
            .in0(N__11539),
            .in1(N__7753),
            .in2(N__7747),
            .in3(N__11660),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_15_9_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_15_9_0 .LUT_INIT=16'b0100111101111111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_15_9_0  (
            .in0(N__7728),
            .in1(N__11522),
            .in2(N__11676),
            .in3(N__7930),
            .lcout(\DUT.rFifoDataror_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_RNI86BE_LC_15_9_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_RNI86BE_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_RNI86BE_LC_15_9_1 .LUT_INIT=16'b1111111100011011;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_0_RNI86BE_LC_15_9_1  (
            .in0(N__11523),
            .in1(N__7716),
            .in2(N__7705),
            .in3(N__11651),
            .lcout(),
            .ltout(\DUT.rFifoDataror_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNIQOK61_0_LC_15_9_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNIQOK61_0_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNIQOK61_0_LC_15_9_2 .LUT_INIT=16'b0000000000111111;
    LogicCell40 \DUT.uart_inst0.tx_state_RNIQOK61_0_LC_15_9_2  (
            .in0(_gnd_net_),
            .in1(N__7690),
            .in2(N__7684),
            .in3(N__11434),
            .lcout(\DUT.uart_inst0.N_145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_15_9_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_15_9_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_15_9_6 .LUT_INIT=16'b1000100011110101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_15_9_6  (
            .in0(N__11652),
            .in1(N__7681),
            .in2(N__7672),
            .in3(N__7660),
            .lcout(\DUT.rFifoDatarx_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNI7FOF_2_LC_15_10_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNI7FOF_2_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNI7FOF_2_LC_15_10_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNI7FOF_2_LC_15_10_0  (
            .in0(_gnd_net_),
            .in1(N__10217),
            .in2(_gnd_net_),
            .in3(N__9910),
            .lcout(\DUT.fifo_tx_inst.N_79 ),
            .ltout(\DUT.fifo_tx_inst.N_79_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_1_LC_15_10_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_1_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_1_LC_15_10_1 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_RNI8BKM_1_LC_15_10_1  (
            .in0(_gnd_net_),
            .in1(N__7652),
            .in2(N__7621),
            .in3(N__7616),
            .lcout(\DUT.fifo_tx_inst.rFifoData_awe2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIFFVH_4_LC_15_10_5 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIFFVH_4_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIFFVH_4_LC_15_10_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_RNIFFVH_4_LC_15_10_5  (
            .in0(_gnd_net_),
            .in1(N__7895),
            .in2(_gnd_net_),
            .in3(N__7913),
            .lcout(\fifo_inst.ftdi_output_inst.N_68_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_0_LC_15_11_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_0_LC_15_11_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoCount_0_LC_15_11_0 .LUT_INIT=16'b1001100110100101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_0_LC_15_11_0  (
            .in0(N__10001),
            .in1(N__9940),
            .in2(N__8989),
            .in3(N__11754),
            .lcout(\DUT.fifo_tx_inst.rFifoCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12780),
            .ce(),
            .sr(N__11111));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_LC_15_11_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_LC_15_11_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_LC_15_11_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_2_LC_15_11_2  (
            .in0(_gnd_net_),
            .in1(N__7941),
            .in2(_gnd_net_),
            .in3(N__7929),
            .lcout(\DUT.fifo_tx_inst.rFifoDataro_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12780),
            .ce(),
            .sr(N__11111));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_3_LC_15_11_3 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_3_LC_15_11_3 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_3_LC_15_11_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_3_LC_15_11_3  (
            .in0(N__11044),
            .in1(N__11241),
            .in2(_gnd_net_),
            .in3(N__10975),
            .lcout(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12780),
            .ce(),
            .sr(N__11111));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_4_LC_15_11_4 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_4_LC_15_11_4 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_4_LC_15_11_4 .LUT_INIT=16'b1111111100001010;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_4_LC_15_11_4  (
            .in0(N__7915),
            .in1(_gnd_net_),
            .in2(N__7900),
            .in3(N__7881),
            .lcout(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12780),
            .ce(),
            .sr(N__11111));
    defparam \fifo_inst.ftdi_output_inst.rWrDelay_LC_15_11_5 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rWrDelay_LC_15_11_5 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rWrDelay_LC_15_11_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \fifo_inst.ftdi_output_inst.rWrDelay_LC_15_11_5  (
            .in0(_gnd_net_),
            .in1(N__7896),
            .in2(_gnd_net_),
            .in3(N__7914),
            .lcout(\fifo_inst.ftdi_output_inst.rWrDelayZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12780),
            .ce(),
            .sr(N__11111));
    defparam \fifo_inst.ftdi_output_inst.oTx_n_LC_15_11_6 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.oTx_n_LC_15_11_6 .SEQ_MODE=4'b1001;
    defparam \fifo_inst.ftdi_output_inst.oTx_n_LC_15_11_6 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \fifo_inst.ftdi_output_inst.oTx_n_LC_15_11_6  (
            .in0(N__11171),
            .in1(N__7847),
            .in2(_gnd_net_),
            .in3(N__7882),
            .lcout(P1A4_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12780),
            .ce(),
            .sr(N__11111));
    defparam \fifo_inst.ftdi_output_inst.rTxBusReady_LC_15_11_7 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rTxBusReady_LC_15_11_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rTxBusReady_LC_15_11_7 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \fifo_inst.ftdi_output_inst.rTxBusReady_LC_15_11_7  (
            .in0(N__7784),
            .in1(N__8995),
            .in2(_gnd_net_),
            .in3(N__11170),
            .lcout(rTxBusReady),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12780),
            .ce(),
            .sr(N__11111));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIO0PE2_11_LC_16_1_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIO0PE2_11_LC_16_1_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIO0PE2_11_LC_16_1_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIO0PE2_11_LC_16_1_0  (
            .in0(N__7767),
            .in1(N__8130),
            .in2(N__8166),
            .in3(N__8145),
            .lcout(\DUT.uart_inst0.rx_clk_divider_5_i_a2_12_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_8_LC_16_1_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_8_LC_16_1_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_8_LC_16_1_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_8_LC_16_1_1  (
            .in0(N__9319),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7768),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12832),
            .ce(N__12345),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_9_LC_16_1_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_9_LC_16_1_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_9_LC_16_1_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_9_LC_16_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8167),
            .in3(N__9318),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12832),
            .ce(N__12345),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_11_LC_16_1_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_11_LC_16_1_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_11_LC_16_1_3 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_11_LC_16_1_3  (
            .in0(N__8146),
            .in1(_gnd_net_),
            .in2(N__9346),
            .in3(_gnd_net_),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12832),
            .ce(N__12345),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_12_LC_16_1_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_12_LC_16_1_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_12_LC_16_1_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_12_LC_16_1_4  (
            .in0(_gnd_net_),
            .in1(N__9317),
            .in2(_gnd_net_),
            .in3(N__8131),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12832),
            .ce(N__12345),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_0_LC_16_1_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_0_LC_16_1_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_0_LC_16_1_5 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_0_LC_16_1_5  (
            .in0(N__9320),
            .in1(N__8114),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12832),
            .ce(N__12345),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIS5BA2_0_LC_16_1_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIS5BA2_0_LC_16_1_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIS5BA2_0_LC_16_1_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIS5BA2_0_LC_16_1_6  (
            .in0(N__8325),
            .in1(N__8079),
            .in2(N__8116),
            .in3(N__8091),
            .lcout(\DUT.uart_inst0.rx_clk_divider_5_i_a2_12_4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_LC_16_1_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_1_LC_16_1_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_LC_16_1_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_LC_16_1_7  (
            .in0(N__8080),
            .in1(_gnd_net_),
            .in2(N__9347),
            .in3(_gnd_net_),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12832),
            .ce(N__12345),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_5_LC_16_2_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_5_LC_16_2_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_5_LC_16_2_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_5_LC_16_2_1  (
            .in0(N__9311),
            .in1(N__9761),
            .in2(_gnd_net_),
            .in3(N__9651),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12829),
            .ce(N__12346),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_1_LC_16_2_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_1_LC_16_2_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_1_LC_16_2_2 .LUT_INIT=16'b0111011100110011;
    LogicCell40 \DUT.uart_inst0.rx_countdown_1_LC_16_2_2  (
            .in0(N__9760),
            .in1(N__9313),
            .in2(_gnd_net_),
            .in3(N__8046),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12829),
            .ce(N__12346),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_2_LC_16_2_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_2_LC_16_2_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_2_LC_16_2_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_2_LC_16_2_3  (
            .in0(_gnd_net_),
            .in1(N__9310),
            .in2(_gnd_net_),
            .in3(N__7972),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12829),
            .ce(N__12346),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_2_LC_16_2_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_2_LC_16_2_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_2_LC_16_2_4 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_2_LC_16_2_4  (
            .in0(N__8395),
            .in1(N__8389),
            .in2(N__8383),
            .in3(N__9652),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12829),
            .ce(N__12346),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_17_LC_16_2_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_17_LC_16_2_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_17_LC_16_2_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_17_LC_16_2_5  (
            .in0(_gnd_net_),
            .in1(N__9309),
            .in2(_gnd_net_),
            .in3(N__8362),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12829),
            .ce(N__12346),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_10_LC_16_2_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_10_LC_16_2_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_10_LC_16_2_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_10_LC_16_2_6  (
            .in0(_gnd_net_),
            .in1(N__9312),
            .in2(_gnd_net_),
            .in3(N__8344),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12829),
            .ce(N__12346),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_13_LC_16_2_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_13_LC_16_2_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_13_LC_16_2_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_13_LC_16_2_7  (
            .in0(_gnd_net_),
            .in1(N__9308),
            .in2(_gnd_net_),
            .in3(N__8326),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12829),
            .ce(N__12346),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_3_2_LC_16_3_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_3_2_LC_16_3_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_3_2_LC_16_3_0 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_3_2_LC_16_3_0  (
            .in0(N__9862),
            .in1(N__8554),
            .in2(_gnd_net_),
            .in3(N__9222),
            .lcout(\DUT.uart_inst0.N_199_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ioFifoData_iobuf_RNO_0_LC_16_3_1.C_ON=1'b0;
    defparam ioFifoData_iobuf_RNO_0_LC_16_3_1.SEQ_MODE=4'b0000;
    defparam ioFifoData_iobuf_RNO_0_LC_16_3_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 ioFifoData_iobuf_RNO_0_LC_16_3_1 (
            .in0(N__11266),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_1239_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNI237O_0_LC_16_3_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNI237O_0_LC_16_3_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNI237O_0_LC_16_3_3 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \DUT.uart_inst0.recv_state_RNI237O_0_LC_16_3_3  (
            .in0(_gnd_net_),
            .in1(N__9861),
            .in2(_gnd_net_),
            .in3(N__8280),
            .lcout(\DUT.uart_inst0.N_149 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_3_LC_16_3_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_3_LC_16_3_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_3_LC_16_3_4 .LUT_INIT=16'b1010000011000000;
    LogicCell40 \DUT.uart_inst0.recv_state_3_LC_16_3_4  (
            .in0(N__9802),
            .in1(N__8713),
            .in2(N__10642),
            .in3(N__8569),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12827),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNI2S9L5_0_LC_16_3_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI2S9L5_0_LC_16_3_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI2S9L5_0_LC_16_3_5 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNI2S9L5_0_LC_16_3_5  (
            .in0(N__8256),
            .in1(N__8236),
            .in2(N__8221),
            .in3(N__8197),
            .lcout(\DUT.uart_inst0.rx_clk_divider_5_i_a2_12_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_2_2_LC_16_3_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_2_2_LC_16_3_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNO_2_2_LC_16_3_7 .LUT_INIT=16'b1011101110111110;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNO_2_2_LC_16_3_7  (
            .in0(N__9223),
            .in1(N__8706),
            .in2(N__8617),
            .in3(N__8674),
            .lcout(\DUT.uart_inst0.N_31_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_1_5_LC_16_4_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_1_5_LC_16_4_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_1_5_LC_16_4_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_1_5_LC_16_4_1  (
            .in0(N__9882),
            .in1(N__9801),
            .in2(_gnd_net_),
            .in3(N__9220),
            .lcout(\DUT.uart_inst0.N_203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_3_LC_16_4_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_3_LC_16_4_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_3_LC_16_4_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_3_LC_16_4_2  (
            .in0(N__8552),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8581),
            .lcout(\DUT.uart_inst0.recv_state_ns_0_i_0_0_a3_0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIUJI11_3_LC_16_4_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIUJI11_3_LC_16_4_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIUJI11_3_LC_16_4_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNIUJI11_3_LC_16_4_3  (
            .in0(N__8707),
            .in1(N__8673),
            .in2(N__8635),
            .in3(N__8609),
            .lcout(\DUT.uart_inst0.N_215_4 ),
            .ltout(\DUT.uart_inst0.N_215_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_2_LC_16_4_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_2_LC_16_4_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_2_LC_16_4_4 .LUT_INIT=16'b0000110010101110;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_2_LC_16_4_4  (
            .in0(N__9221),
            .in1(N__8557),
            .in2(N__8575),
            .in3(N__9881),
            .lcout(),
            .ltout(\DUT.uart_inst0.recv_state_srsts_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_2_LC_16_4_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_2_LC_16_4_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_2_LC_16_4_5 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \DUT.uart_inst0.recv_state_2_LC_16_4_5  (
            .in0(N__10634),
            .in1(N__8553),
            .in2(N__8572),
            .in3(N__8568),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12823),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNIBTG71_2_LC_16_4_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNIBTG71_2_LC_16_4_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNIBTG71_2_LC_16_4_7 .LUT_INIT=16'b1000101010001000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNIBTG71_2_LC_16_4_7  (
            .in0(N__12423),
            .in1(N__8551),
            .in2(N__9883),
            .in3(N__9219),
            .lcout(\DUT.uart_inst0.g0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_2_LC_16_5_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_2_LC_16_5_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_2_LC_16_5_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_2_LC_16_5_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8482),
            .lcout(\DUT.wRxByte_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12819),
            .ce(N__8419),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_16_6_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_16_6_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_16_6_0 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_16_6_0  (
            .in0(N__8875),
            .in1(N__11659),
            .in2(N__8869),
            .in3(N__8824),
            .lcout(\DUT.rFifoDatarx_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_16_6_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_16_6_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_16_6_1 .LUT_INIT=16'b1010000011011101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_16_6_1  (
            .in0(N__11658),
            .in1(N__8860),
            .in2(N__8854),
            .in3(N__8845),
            .lcout(\DUT.rFifoDatarx_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_16_6_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_16_6_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_16_6_5 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_16_6_5  (
            .in0(N__11537),
            .in1(N__8836),
            .in2(N__11677),
            .in3(N__10126),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_16_6_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_16_6_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_16_6_6 .LUT_INIT=16'b0001000111001111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_16_6_6  (
            .in0(N__8818),
            .in1(N__11656),
            .in2(N__8806),
            .in3(N__11538),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_16_6_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_16_6_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_16_6_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_16_6_7  (
            .in0(N__11657),
            .in1(N__8791),
            .in2(N__8785),
            .in3(N__8782),
            .lcout(\DUT.rFifoDatarx_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_0_LC_16_7_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_0_LC_16_7_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_0_LC_16_7_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \DUT.uart_inst0.tx_data_0_LC_16_7_0  (
            .in0(N__8776),
            .in1(N__9148),
            .in2(N__8743),
            .in3(N__11436),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12811),
            .ce(N__9102),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_RNO_0_LC_16_7_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_RNO_0_LC_16_7_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_out_RNO_0_LC_16_7_2 .LUT_INIT=16'b1111101011111110;
    LogicCell40 \DUT.uart_inst0.tx_out_RNO_0_LC_16_7_2  (
            .in0(N__8902),
            .in1(N__8908),
            .in2(N__9007),
            .in3(N__10859),
            .lcout(\DUT.uart_inst0.tx_out_6_iv_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_1_LC_16_7_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_1_LC_16_7_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_1_LC_16_7_4 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \DUT.uart_inst0.tx_data_1_LC_16_7_4  (
            .in0(N__8959),
            .in1(N__8749),
            .in2(N__11443),
            .in3(N__9149),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12811),
            .ce(N__9102),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_2_LC_16_7_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_2_LC_16_7_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_2_LC_16_7_5 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \DUT.uart_inst0.tx_data_2_LC_16_7_5  (
            .in0(N__11435),
            .in1(N__8734),
            .in2(N__9154),
            .in3(N__8947),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12811),
            .ce(N__9102),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_3_LC_16_7_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_3_LC_16_7_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_3_LC_16_7_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \DUT.uart_inst0.tx_data_3_LC_16_7_6  (
            .in0(N__8953),
            .in1(N__9153),
            .in2(N__9172),
            .in3(N__11437),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12811),
            .ce(N__9102),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_16_8_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_16_8_0 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_16_8_0  (
            .in0(N__11542),
            .in1(N__8938),
            .in2(N__11679),
            .in3(N__10087),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_16_8_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_16_8_1 .LUT_INIT=16'b1100101100001011;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_16_8_1  (
            .in0(N__8926),
            .in1(N__11670),
            .in2(N__8917),
            .in3(N__8914),
            .lcout(\DUT.rFifoDatarx_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNINQKO8_0_0_LC_16_8_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNINQKO8_0_0_LC_16_8_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNINQKO8_0_0_LC_16_8_4 .LUT_INIT=16'b0001000000110000;
    LogicCell40 \DUT.uart_inst0.tx_state_RNINQKO8_0_0_LC_16_8_4  (
            .in0(N__11433),
            .in1(N__11461),
            .in2(N__12441),
            .in3(N__10852),
            .lcout(\DUT.uart_inst0.N_22_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_RNO_1_LC_16_8_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_RNO_1_LC_16_8_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_out_RNO_1_LC_16_8_5 .LUT_INIT=16'b0100010001000000;
    LogicCell40 \DUT.uart_inst0.tx_out_RNO_1_LC_16_8_5  (
            .in0(N__11821),
            .in1(N__11432),
            .in2(N__9081),
            .in3(N__10769),
            .lcout(\DUT.uart_inst0.tx_out_6_iv_0_a3_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_RNO_3_LC_16_8_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_RNO_3_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_out_RNO_3_LC_16_8_6 .LUT_INIT=16'b1000000010001100;
    LogicCell40 \DUT.uart_inst0.tx_out_RNO_3_LC_16_8_6  (
            .in0(N__10770),
            .in1(N__9053),
            .in2(N__11442),
            .in3(N__11746),
            .lcout(\DUT.uart_inst0.N_101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_5_LC_16_9_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_5_LC_16_9_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_5_LC_16_9_0 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \DUT.uart_inst0.tx_data_5_LC_16_9_0  (
            .in0(N__11406),
            .in1(N__8896),
            .in2(N__8884),
            .in3(N__9137),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12798),
            .ce(N__9109),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_6_LC_16_9_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_6_LC_16_9_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_6_LC_16_9_1 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \DUT.uart_inst0.tx_data_6_LC_16_9_1  (
            .in0(N__9138),
            .in1(N__8890),
            .in2(N__9118),
            .in3(N__11408),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12798),
            .ce(N__9109),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_4_LC_16_9_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_4_LC_16_9_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_4_LC_16_9_5 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \DUT.uart_inst0.tx_data_4_LC_16_9_5  (
            .in0(N__9136),
            .in1(N__9187),
            .in2(N__9181),
            .in3(N__11407),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12798),
            .ce(N__9109),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_7_LC_16_9_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_7_LC_16_9_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_7_LC_16_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \DUT.uart_inst0.tx_data_7_LC_16_9_6  (
            .in0(_gnd_net_),
            .in1(N__9160),
            .in2(_gnd_net_),
            .in3(N__9135),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12798),
            .ce(N__9109),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNI0AJL_0_LC_16_10_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNI0AJL_0_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNI0AJL_0_LC_16_10_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNI0AJL_0_LC_16_10_0  (
            .in0(_gnd_net_),
            .in1(N__10218),
            .in2(_gnd_net_),
            .in3(N__11832),
            .lcout(\DUT.fifo_tx_inst.N_83 ),
            .ltout(\DUT.fifo_tx_inst.N_83_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNISSQ21_1_LC_16_10_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNISSQ21_1_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNISSQ21_1_LC_16_10_1 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNISSQ21_1_LC_16_10_1  (
            .in0(N__11749),
            .in1(_gnd_net_),
            .in2(N__9085),
            .in3(N__9963),
            .lcout(\DUT.fifo_tx_inst.rFifoCount_RNISSQ21Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_RNO_2_LC_16_10_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_RNO_2_LC_16_10_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_out_RNO_2_LC_16_10_2 .LUT_INIT=16'b1000000011000000;
    LogicCell40 \DUT.uart_inst0.tx_out_RNO_2_LC_16_10_2  (
            .in0(N__9082),
            .in1(N__11801),
            .in2(N__9064),
            .in3(N__11370),
            .lcout(\DUT.uart_inst0.N_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNI7AJQ_0_0_LC_16_10_3 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNI7AJQ_0_0_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNI7AJQ_0_0_LC_16_10_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_RNI7AJQ_0_0_LC_16_10_3  (
            .in0(N__11054),
            .in1(N__11250),
            .in2(_gnd_net_),
            .in3(N__10939),
            .lcout(\fifo_inst.ftdi_output_inst.rFifoStatec_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIN9O8_0_LC_16_10_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIN9O8_0_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIN9O8_0_LC_16_10_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNIN9O8_0_LC_16_10_4  (
            .in0(N__9906),
            .in1(N__9961),
            .in2(_gnd_net_),
            .in3(N__9993),
            .lcout(\DUT.N_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIME2J_0_LC_16_10_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIME2J_0_LC_16_10_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIME2J_0_LC_16_10_6 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNIME2J_0_LC_16_10_6  (
            .in0(N__9962),
            .in1(N__9994),
            .in2(N__9915),
            .in3(N__11747),
            .lcout(\DUT.fifo_tx_inst.rReadPtr11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_16_10_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_16_10_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_16_10_7 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_16_10_7  (
            .in0(N__11748),
            .in1(N__8981),
            .in2(N__10002),
            .in3(N__9938),
            .lcout(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_16_11_0 .C_ON=1'b1;
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_16_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_16_11_0  (
            .in0(_gnd_net_),
            .in1(N__10009),
            .in2(N__10003),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_11_0_),
            .carryout(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_1_LC_16_11_1 .C_ON=1'b1;
    defparam \DUT.fifo_tx_inst.rFifoCount_1_LC_16_11_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoCount_1_LC_16_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_1_LC_16_11_1  (
            .in0(_gnd_net_),
            .in1(N__9964),
            .in2(N__9973),
            .in3(N__9943),
            .lcout(\DUT.fifo_tx_inst.rFifoCountZ0Z_1 ),
            .ltout(),
            .carryin(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0 ),
            .carryout(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1 ),
            .clk(N__12786),
            .ce(),
            .sr(N__11114));
    defparam \DUT.fifo_tx_inst.rFifoCount_2_LC_16_11_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_2_LC_16_11_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoCount_2_LC_16_11_2 .LUT_INIT=16'b0110010110011010;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_2_LC_16_11_2  (
            .in0(N__9914),
            .in1(N__9939),
            .in2(N__11755),
            .in3(N__9922),
            .lcout(\DUT.fifo_tx_inst.rFifoCountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12786),
            .ce(),
            .sr(N__11114));
    defparam \DUT.uart_inst0.recv_state_RNO_0_6_LC_17_2_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_6_LC_17_2_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_6_LC_17_2_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_6_LC_17_2_7  (
            .in0(N__9870),
            .in1(N__12422),
            .in2(_gnd_net_),
            .in3(N__9800),
            .lcout(\DUT.uart_inst0.g0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_4_LC_17_3_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_4_LC_17_3_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_4_LC_17_3_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_4_LC_17_3_3  (
            .in0(N__9770),
            .in1(N__9314),
            .in2(_gnd_net_),
            .in3(N__9721),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12830),
            .ce(N__12353),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_1_1_LC_17_4_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_1_1_LC_17_4_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_1_1_LC_17_4_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_1_1_LC_17_4_1  (
            .in0(_gnd_net_),
            .in1(N__9650),
            .in2(_gnd_net_),
            .in3(N__9586),
            .lcout(),
            .ltout(\DUT.uart_inst0.G_10_i_a4_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_1_LC_17_4_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_1_LC_17_4_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_1_LC_17_4_2 .LUT_INIT=16'b0101000000010000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_1_LC_17_4_2  (
            .in0(N__9577),
            .in1(N__9505),
            .in2(N__9439),
            .in3(N__9436),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_4_i_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_1_LC_17_4_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_1_LC_17_4_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_1_LC_17_4_3 .LUT_INIT=16'b0000100000001010;
    LogicCell40 \DUT.uart_inst0.recv_state_1_LC_17_4_3  (
            .in0(N__10641),
            .in1(N__9234),
            .in2(N__9367),
            .in3(N__9315),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12828),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_0_LC_17_5_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_0_LC_17_5_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoCount_0_LC_17_5_0 .LUT_INIT=16'b1010101001011001;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_0_LC_17_5_0  (
            .in0(N__10403),
            .in1(N__10456),
            .in2(N__10252),
            .in3(N__10432),
            .lcout(\DUT.fifo_rx_inst.rFifoCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12824),
            .ce(),
            .sr(N__11130));
    defparam \fifo_inst.ftdi_output_inst.oRxFlag_LC_17_5_2 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.oRxFlag_LC_17_5_2 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.oRxFlag_LC_17_5_2 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \fifo_inst.ftdi_output_inst.oRxFlag_LC_17_5_2  (
            .in0(N__10790),
            .in1(N__10367),
            .in2(_gnd_net_),
            .in3(N__10302),
            .lcout(P1A2_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12824),
            .ce(),
            .sr(N__11130));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_2_LC_17_5_4 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_2_LC_17_5_4 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_2_LC_17_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_2_LC_17_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10368),
            .lcout(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12824),
            .ce(),
            .sr(N__11130));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_1_LC_17_5_6 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_1_LC_17_5_6 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_1_LC_17_5_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_1_LC_17_5_6  (
            .in0(_gnd_net_),
            .in1(N__11059),
            .in2(_gnd_net_),
            .in3(N__10970),
            .lcout(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12824),
            .ce(),
            .sr(N__11130));
    defparam rTxWrite_LC_17_6_0.C_ON=1'b0;
    defparam rTxWrite_LC_17_6_0.SEQ_MODE=4'b1000;
    defparam rTxWrite_LC_17_6_0.LUT_INIT=16'b1111111111001100;
    LogicCell40 rTxWrite_LC_17_6_0 (
            .in0(_gnd_net_),
            .in1(N__10301),
            .in2(_gnd_net_),
            .in3(N__10251),
            .lcout(rTxWriteZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12820),
            .ce(),
            .sr(N__11129));
    defparam \fifo_inst.ftdi_output_inst.oRx_n_LC_17_6_1 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.oRx_n_LC_17_6_1 .SEQ_MODE=4'b1001;
    defparam \fifo_inst.ftdi_output_inst.oRx_n_LC_17_6_1 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \fifo_inst.ftdi_output_inst.oRx_n_LC_17_6_1  (
            .in0(N__10791),
            .in1(N__10175),
            .in2(_gnd_net_),
            .in3(N__10906),
            .lcout(P1A3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12820),
            .ce(),
            .sr(N__11129));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_17_7_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_17_7_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_17_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_17_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10159),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12817),
            .ce(N__10081),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_17_7_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_17_7_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_17_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_17_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10116),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12817),
            .ce(N__10081),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_17_8_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_17_8_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_17_8_0 .LUT_INIT=16'b0000000011111110;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_17_8_0  (
            .in0(N__10660),
            .in1(N__10695),
            .in2(N__10683),
            .in3(N__10495),
            .lcout(\DUT.uart_inst0.un1_tx_bits_remaining_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_2_LC_17_8_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_2_LC_17_8_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_bits_remaining_2_LC_17_8_1 .LUT_INIT=16'b1010101010101001;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_2_LC_17_8_1  (
            .in0(N__10696),
            .in1(N__10682),
            .in2(N__10501),
            .in3(N__10663),
            .lcout(\DUT.uart_inst0.tx_bits_remainingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12812),
            .ce(),
            .sr(N__11845));
    defparam \DUT.uart_inst0.tx_bits_remaining_1_LC_17_8_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_1_LC_17_8_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_bits_remaining_1_LC_17_8_2 .LUT_INIT=16'b1111000010100101;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_1_LC_17_8_2  (
            .in0(N__10662),
            .in1(_gnd_net_),
            .in2(N__10684),
            .in3(N__10497),
            .lcout(\DUT.uart_inst0.tx_bits_remainingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12812),
            .ce(),
            .sr(N__11845));
    defparam \DUT.uart_inst0.tx_bits_remaining_0_LC_17_8_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_0_LC_17_8_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_bits_remaining_0_LC_17_8_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_0_LC_17_8_3  (
            .in0(N__10496),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10661),
            .lcout(\DUT.uart_inst0.tx_bits_remainingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12812),
            .ce(),
            .sr(N__11845));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_3_LC_17_8_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_3_LC_17_8_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_3_LC_17_8_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_3_LC_17_8_5  (
            .in0(N__10694),
            .in1(N__10675),
            .in2(N__10471),
            .in3(N__10659),
            .lcout(\DUT.uart_inst0.N_142 ),
            .ltout(\DUT.uart_inst0.N_142_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNIJ5C81_1_LC_17_8_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNIJ5C81_1_LC_17_8_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNIJ5C81_1_LC_17_8_6 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \DUT.uart_inst0.tx_state_RNIJ5C81_1_LC_17_8_6  (
            .in0(_gnd_net_),
            .in1(N__11804),
            .in2(N__10645),
            .in3(N__11391),
            .lcout(\DUT.uart_inst0.N_144 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNI6Q5N3_1_LC_17_8_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNI6Q5N3_1_LC_17_8_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNI6Q5N3_1_LC_17_8_7 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \DUT.uart_inst0.tx_state_RNI6Q5N3_1_LC_17_8_7  (
            .in0(N__11392),
            .in1(N__10726),
            .in2(N__11818),
            .in3(N__10771),
            .lcout(\DUT.uart_inst0.N_146 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNI3MLP6_3_LC_17_9_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNI3MLP6_3_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNI3MLP6_3_LC_17_9_0 .LUT_INIT=16'b0101111100001010;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNI3MLP6_3_LC_17_9_0  (
            .in0(N__12244),
            .in1(_gnd_net_),
            .in2(N__10888),
            .in3(N__10721),
            .lcout(\DUT.uart_inst0.N_84 ),
            .ltout(\DUT.uart_inst0.N_84_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNINQKO8_0_LC_17_9_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNINQKO8_0_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNINQKO8_0_LC_17_9_1 .LUT_INIT=16'b1111110111011101;
    LogicCell40 \DUT.uart_inst0.tx_state_RNINQKO8_0_LC_17_9_1  (
            .in0(N__10625),
            .in1(N__11459),
            .in2(N__10504),
            .in3(N__11395),
            .lcout(\DUT.uart_inst0.N_22 ),
            .ltout(\DUT.uart_inst0.N_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_3_LC_17_9_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_3_LC_17_9_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_bits_remaining_3_LC_17_9_2 .LUT_INIT=16'b0111110111010111;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_3_LC_17_9_2  (
            .in0(N__10897),
            .in1(N__10470),
            .in2(N__10480),
            .in3(N__10477),
            .lcout(\DUT.uart_inst0.tx_bits_remainingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12805),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNICODU_0_LC_17_9_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNICODU_0_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNICODU_0_LC_17_9_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DUT.uart_inst0.tx_state_RNICODU_0_LC_17_9_3  (
            .in0(N__10768),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11394),
            .lcout(\DUT.uart_inst0.N_143 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNO_0_0_LC_17_9_4 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNO_0_0_LC_17_9_4 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNO_0_0_LC_17_9_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_RNO_0_0_LC_17_9_4  (
            .in0(N__11254),
            .in1(N__11055),
            .in2(_gnd_net_),
            .in3(N__10946),
            .lcout(),
            .ltout(\fifo_inst.ftdi_output_inst.N_78_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_0_LC_17_9_5 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_0_LC_17_9_5 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_0_LC_17_9_5 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_0_LC_17_9_5  (
            .in0(N__10795),
            .in1(N__12433),
            .in2(N__10774),
            .in3(N__11182),
            .lcout(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12805),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNIIAMI1_1_LC_17_9_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNIIAMI1_1_LC_17_9_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNIIAMI1_1_LC_17_9_6 .LUT_INIT=16'b1111101111110001;
    LogicCell40 \DUT.uart_inst0.tx_state_RNIIAMI1_1_LC_17_9_6  (
            .in0(N__11393),
            .in1(N__11712),
            .in2(N__11819),
            .in3(N__10767),
            .lcout(\DUT.uart_inst0.N_74 ),
            .ltout(\DUT.uart_inst0.N_74_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNILHU57_1_LC_17_9_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNILHU57_1_LC_17_9_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNILHU57_1_LC_17_9_7 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \DUT.uart_inst0.tx_state_RNILHU57_1_LC_17_9_7  (
            .in0(N__10747),
            .in1(N__10883),
            .in2(N__10741),
            .in3(N__12243),
            .lcout(\DUT.uart_inst0.tx_countdown_7s2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNIFE3O7_0_LC_17_10_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNIFE3O7_0_LC_17_10_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNIFE3O7_0_LC_17_10_0 .LUT_INIT=16'b1011000000010000;
    LogicCell40 \DUT.uart_inst0.tx_state_RNIFE3O7_0_LC_17_10_0  (
            .in0(N__12224),
            .in1(N__10725),
            .in2(N__10738),
            .in3(N__10887),
            .lcout(\DUT.uart_inst0.N_30_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNI45HK1_2_LC_17_10_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNI45HK1_2_LC_17_10_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNI45HK1_2_LC_17_10_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNI45HK1_2_LC_17_10_3  (
            .in0(N__12133),
            .in1(N__12006),
            .in2(N__12049),
            .in3(N__11976),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_state_ns_i_i_o2_0_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNIJKPE2_3_LC_17_10_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNIJKPE2_3_LC_17_10_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNIJKPE2_3_LC_17_10_4 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNIJKPE2_3_LC_17_10_4  (
            .in0(N__11874),
            .in1(_gnd_net_),
            .in2(N__10729),
            .in3(N__12079),
            .lcout(\DUT.uart_inst0.N_75 ),
            .ltout(\DUT.uart_inst0.N_75_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNIBVOQB_0_LC_17_10_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNIBVOQB_0_LC_17_10_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNIBVOQB_0_LC_17_10_5 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \DUT.uart_inst0.tx_state_RNIBVOQB_0_LC_17_10_5  (
            .in0(N__11371),
            .in1(N__12223),
            .in2(N__10705),
            .in3(N__10702),
            .lcout(\DUT.uart_inst0.tx_countdown_7_sm0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNI34HK1_2_LC_17_10_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNI34HK1_2_LC_17_10_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNI34HK1_2_LC_17_10_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNI34HK1_2_LC_17_10_6  (
            .in0(N__11975),
            .in1(N__12132),
            .in2(N__12010),
            .in3(N__12078),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_state_ns_i_i_o2_a0_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNIJKPE2_0_3_LC_17_10_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNIJKPE2_0_3_LC_17_10_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNIJKPE2_0_3_LC_17_10_7 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNIJKPE2_0_3_LC_17_10_7  (
            .in0(N__12042),
            .in1(_gnd_net_),
            .in2(N__10891),
            .in3(N__11873),
            .lcout(\DUT.uart_inst0.N_69_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_2_LC_17_11_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_2_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_2_LC_17_11_0 .LUT_INIT=16'b0001111000001111;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_0_2_LC_17_11_0  (
            .in0(N__12084),
            .in1(N__12046),
            .in2(N__12139),
            .in3(N__12245),
            .lcout(\DUT.uart_inst0.tx_countdown_7_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_17_11_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_17_11_1 .LUT_INIT=16'b1111000011100001;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_17_11_1  (
            .in0(N__12045),
            .in1(N__12135),
            .in2(N__11884),
            .in3(N__12083),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_countdown_30_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_17_11_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_17_11_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_17_11_2 .LUT_INIT=16'b0001000100001111;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_17_11_2  (
            .in0(N__11882),
            .in1(N__12246),
            .in2(N__10870),
            .in3(N__11917),
            .lcout(\DUT.uart_inst0.tx_countdown_7_ns_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_1_LC_17_11_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_1_LC_17_11_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_state_1_LC_17_11_5 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \DUT.uart_inst0.tx_state_1_LC_17_11_5  (
            .in0(N__10827),
            .in1(N__10860),
            .in2(_gnd_net_),
            .in3(N__11802),
            .lcout(\DUT.tx_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12792),
            .ce(),
            .sr(N__11119));
    defparam \DUT.uart_inst0.tx_state_0_LC_17_11_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_0_LC_17_11_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_state_0_LC_17_11_7 .LUT_INIT=16'b0000000001010100;
    LogicCell40 \DUT.uart_inst0.tx_state_0_LC_17_11_7  (
            .in0(N__10828),
            .in1(N__11753),
            .in2(N__11427),
            .in3(N__11803),
            .lcout(\DUT.tx_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12792),
            .ce(),
            .sr(N__11119));
    defparam ioFifoData_iobuf_RNO_3_LC_18_1_7.C_ON=1'b0;
    defparam ioFifoData_iobuf_RNO_3_LC_18_1_7.SEQ_MODE=4'b0000;
    defparam ioFifoData_iobuf_RNO_3_LC_18_1_7.LUT_INIT=16'b0101010101010101;
    LogicCell40 ioFifoData_iobuf_RNO_3_LC_18_1_7 (
            .in0(N__11275),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_1242_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam ioFifoData_iobuf_RNO_1_LC_18_3_3.C_ON=1'b0;
    defparam ioFifoData_iobuf_RNO_1_LC_18_3_3.SEQ_MODE=4'b0000;
    defparam ioFifoData_iobuf_RNO_1_LC_18_3_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 ioFifoData_iobuf_RNO_1_LC_18_3_3 (
            .in0(N__11281),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(N_1240_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rTxBusReady_rep1_i_ess_LC_18_4_0 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rTxBusReady_rep1_i_ess_LC_18_4_0 .SEQ_MODE=4'b1001;
    defparam \fifo_inst.ftdi_output_inst.rTxBusReady_rep1_i_ess_LC_18_4_0 .LUT_INIT=16'b1111010111111111;
    LogicCell40 \fifo_inst.ftdi_output_inst.rTxBusReady_rep1_i_ess_LC_18_4_0  (
            .in0(N__10972),
            .in1(_gnd_net_),
            .in2(N__11249),
            .in3(N__11041),
            .lcout(rTxBusReady_rep1_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12831),
            .ce(N__11065),
            .sr(N__11134));
    defparam \fifo_inst.ftdi_output_inst.rTxBusReady_rep3_i_ess_LC_18_4_1 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rTxBusReady_rep3_i_ess_LC_18_4_1 .SEQ_MODE=4'b1001;
    defparam \fifo_inst.ftdi_output_inst.rTxBusReady_rep3_i_ess_LC_18_4_1 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \fifo_inst.ftdi_output_inst.rTxBusReady_rep3_i_ess_LC_18_4_1  (
            .in0(N__11043),
            .in1(N__11240),
            .in2(_gnd_net_),
            .in3(N__10974),
            .lcout(rTxBusReady_rep3_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12831),
            .ce(N__11065),
            .sr(N__11134));
    defparam \fifo_inst.ftdi_output_inst.rTxBusReady_rep0_i_ess_LC_18_4_3 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rTxBusReady_rep0_i_ess_LC_18_4_3 .SEQ_MODE=4'b1001;
    defparam \fifo_inst.ftdi_output_inst.rTxBusReady_rep0_i_ess_LC_18_4_3 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \fifo_inst.ftdi_output_inst.rTxBusReady_rep0_i_ess_LC_18_4_3  (
            .in0(N__11040),
            .in1(N__11235),
            .in2(_gnd_net_),
            .in3(N__10971),
            .lcout(rTxBusReady_rep0_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12831),
            .ce(N__11065),
            .sr(N__11134));
    defparam \fifo_inst.ftdi_output_inst.rTxBusReady_rep2_i_ess_LC_18_4_5 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rTxBusReady_rep2_i_ess_LC_18_4_5 .SEQ_MODE=4'b1001;
    defparam \fifo_inst.ftdi_output_inst.rTxBusReady_rep2_i_ess_LC_18_4_5 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \fifo_inst.ftdi_output_inst.rTxBusReady_rep2_i_ess_LC_18_4_5  (
            .in0(N__11042),
            .in1(N__11239),
            .in2(_gnd_net_),
            .in3(N__10973),
            .lcout(rTxBusReady_rep2_i_ess),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12831),
            .ce(N__11065),
            .sr(N__11134));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIMPIC1_0_LC_18_5_1 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIMPIC1_0_LC_18_5_1 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIMPIC1_0_LC_18_5_1 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_RNIMPIC1_0_LC_18_5_1  (
            .in0(N__11039),
            .in1(N__10969),
            .in2(N__11248),
            .in3(N__11181),
            .lcout(),
            .ltout(\fifo_inst.ftdi_output_inst.un1_oTx_n_1_sqmuxa_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNII7TE1_0_LC_18_5_2 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNII7TE1_0_LC_18_5_2 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNII7TE1_0_LC_18_5_2 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_RNII7TE1_0_LC_18_5_2  (
            .in0(N__11149),
            .in1(_gnd_net_),
            .in2(N__11068),
            .in3(_gnd_net_),
            .lcout(\fifo_inst.ftdi_output_inst.un1_oTx_n_1_sqmuxa_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIR68B_0_LC_18_6_7 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIR68B_0_LC_18_6_7 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIR68B_0_LC_18_6_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_RNIR68B_0_LC_18_6_7  (
            .in0(_gnd_net_),
            .in1(N__11038),
            .in2(_gnd_net_),
            .in3(N__10956),
            .lcout(\fifo_inst.ftdi_output_inst.N_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNICU6U_1_LC_18_8_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNICU6U_1_LC_18_8_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNICU6U_1_LC_18_8_2 .LUT_INIT=16'b1111111110111011;
    LogicCell40 \DUT.uart_inst0.tx_state_RNICU6U_1_LC_18_8_2  (
            .in0(N__11808),
            .in1(N__11711),
            .in2(_gnd_net_),
            .in3(N__11428),
            .lcout(\DUT.uart_inst0.N_77 ),
            .ltout(\DUT.uart_inst0.N_77_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNI8CH01_1_LC_18_8_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNI8CH01_1_LC_18_8_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNI8CH01_1_LC_18_8_3 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \DUT.uart_inst0.tx_state_RNI8CH01_1_LC_18_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10900),
            .in3(N__12432),
            .lcout(\DUT.uart_inst0.tx_state_RNI8CH01Z0Z_1 ),
            .ltout(\DUT.uart_inst0.tx_state_RNI8CH01Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNI8CH01_0_1_LC_18_8_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNI8CH01_0_1_LC_18_8_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNI8CH01_0_1_LC_18_8_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \DUT.uart_inst0.tx_state_RNI8CH01_0_1_LC_18_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11848),
            .in3(_gnd_net_),
            .lcout(\DUT.uart_inst0.N_59_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.rTransmit_LC_18_9_2 .C_ON=1'b0;
    defparam \DUT.rTransmit_LC_18_9_2 .SEQ_MODE=4'b1000;
    defparam \DUT.rTransmit_LC_18_9_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \DUT.rTransmit_LC_18_9_2  (
            .in0(N__11423),
            .in1(N__11839),
            .in2(N__11820),
            .in3(N__12437),
            .lcout(\DUT.rTransmitZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12813),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rReadPtr_1_LC_18_9_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rReadPtr_1_LC_18_9_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rReadPtr_1_LC_18_9_4 .LUT_INIT=16'b0000000001101100;
    LogicCell40 \DUT.fifo_tx_inst.rReadPtr_1_LC_18_9_4  (
            .in0(N__11563),
            .in1(N__11603),
            .in2(N__11534),
            .in3(N__11569),
            .lcout(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12813),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rReadPtr_RNILV421_0_LC_18_9_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rReadPtr_RNILV421_0_LC_18_9_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rReadPtr_RNILV421_0_LC_18_9_5 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \DUT.fifo_tx_inst.rReadPtr_RNILV421_0_LC_18_9_5  (
            .in0(N__11602),
            .in1(N__11507),
            .in2(N__12442),
            .in3(N__11561),
            .lcout(\DUT.fifo_tx_inst.un1_i11_2_i ),
            .ltout(\DUT.fifo_tx_inst.un1_i11_2_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rReadPtr_0_LC_18_9_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rReadPtr_0_LC_18_9_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rReadPtr_0_LC_18_9_6 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \DUT.fifo_tx_inst.rReadPtr_0_LC_18_9_6  (
            .in0(N__11562),
            .in1(_gnd_net_),
            .in2(N__11545),
            .in3(N__11511),
            .lcout(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12813),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_2_LC_18_9_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_2_LC_18_9_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_2_LC_18_9_7 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_1_2_LC_18_9_7  (
            .in0(N__11953),
            .in1(N__11460),
            .in2(_gnd_net_),
            .in3(N__11422),
            .lcout(\DUT.uart_inst0.N_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_0_LC_18_10_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_0_LC_18_10_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_0_LC_18_10_2 .LUT_INIT=16'b0000101001000000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_0_LC_18_10_2  (
            .in0(N__12085),
            .in1(N__12281),
            .in2(N__12250),
            .in3(N__11920),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12806),
            .ce(N__12375),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_4_LC_18_10_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_4_LC_18_10_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_4_LC_18_10_3 .LUT_INIT=16'b0001101101000100;
    LogicCell40 \DUT.uart_inst0.tx_countdown_4_LC_18_10_3  (
            .in0(N__11918),
            .in1(N__12109),
            .in2(N__12247),
            .in3(N__11980),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12806),
            .ce(N__12375),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_2_LC_18_10_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_2_LC_18_10_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_2_LC_18_10_4 .LUT_INIT=16'b0001000101111111;
    LogicCell40 \DUT.uart_inst0.tx_countdown_2_LC_18_10_4  (
            .in0(N__11296),
            .in1(N__12230),
            .in2(N__11290),
            .in3(N__11921),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12806),
            .ce(N__12375),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_5_LC_18_10_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_5_LC_18_10_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_5_LC_18_10_5 .LUT_INIT=16'b0001101101000100;
    LogicCell40 \DUT.uart_inst0.tx_countdown_5_LC_18_10_5  (
            .in0(N__11919),
            .in1(N__12091),
            .in2(N__12248),
            .in3(N__12009),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12806),
            .ce(N__12375),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNIUUGK1_2_LC_18_11_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNIUUGK1_2_LC_18_11_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNIUUGK1_2_LC_18_11_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNIUUGK1_2_LC_18_11_0  (
            .in0(N__12044),
            .in1(N__12134),
            .in2(N__11883),
            .in3(N__12081),
            .lcout(\DUT.uart_inst0.tx_countdown_0_c4 ),
            .ltout(\DUT.uart_inst0.tx_countdown_0_c4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_4_LC_18_11_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_4_LC_18_11_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_4_LC_18_11_1 .LUT_INIT=16'b0000111100101110;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_0_4_LC_18_11_1  (
            .in0(N__11978),
            .in1(N__12157),
            .in2(N__12112),
            .in3(N__11942),
            .lcout(\DUT.uart_inst0.tx_countdown_7_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_1_LC_18_11_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_1_LC_18_11_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_1_LC_18_11_2 .LUT_INIT=16'b0000010011111110;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_0_1_LC_18_11_2  (
            .in0(N__11943),
            .in1(N__12047),
            .in2(N__12163),
            .in3(N__12082),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_countdown_7_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_1_LC_18_11_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_1_LC_18_11_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_1_LC_18_11_3 .LUT_INIT=16'b0010001001011010;
    LogicCell40 \DUT.uart_inst0.tx_countdown_1_LC_18_11_3  (
            .in0(N__12048),
            .in1(N__12249),
            .in2(N__12103),
            .in3(N__11925),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12799),
            .ce(N__12376),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_5_LC_18_11_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_5_LC_18_11_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_5_LC_18_11_4 .LUT_INIT=16'b0100010001001110;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_0_5_LC_18_11_4  (
            .in0(N__12158),
            .in1(N__12008),
            .in2(N__12100),
            .in3(N__11979),
            .lcout(\DUT.uart_inst0.tx_countdown_7_ns_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_3_2_LC_18_11_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_3_2_LC_18_11_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_3_2_LC_18_11_5 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_3_2_LC_18_11_5  (
            .in0(N__12080),
            .in1(N__11875),
            .in2(_gnd_net_),
            .in3(N__12043),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_countdown_7_m1_0_o2_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_2_2_LC_18_11_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_2_2_LC_18_11_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_2_2_LC_18_11_6 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_2_2_LC_18_11_6  (
            .in0(_gnd_net_),
            .in1(N__12007),
            .in2(N__11983),
            .in3(N__11977),
            .lcout(\DUT.uart_inst0.N_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_3_LC_18_11_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_3_LC_18_11_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_3_LC_18_11_7 .LUT_INIT=16'b1100000011111110;
    LogicCell40 \DUT.uart_inst0.tx_countdown_3_LC_18_11_7  (
            .in0(N__12162),
            .in1(N__11944),
            .in2(N__11926),
            .in3(N__11890),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12799),
            .ce(N__12376),
            .sr(_gnd_net_));
    defparam ioFifoData_iobuf_RNO_2_LC_20_2_6.C_ON=1'b0;
    defparam ioFifoData_iobuf_RNO_2_LC_20_2_6.SEQ_MODE=4'b0000;
    defparam ioFifoData_iobuf_RNO_2_LC_20_2_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 ioFifoData_iobuf_RNO_2_LC_20_2_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12478),
            .lcout(N_1241_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_RNIA7A5_4_LC_20_9_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNIA7A5_4_LC_20_9_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNIA7A5_4_LC_20_9_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNIA7A5_4_LC_20_9_2  (
            .in0(N__12525),
            .in1(N__12543),
            .in2(N__12511),
            .in3(N__12558),
            .lcout(\DUT.uart_inst0.un1_tx_clk_divider_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_RNIHKCN_13_LC_20_10_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNIHKCN_13_LC_20_10_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNIHKCN_13_LC_20_10_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNIHKCN_13_LC_20_10_1  (
            .in0(_gnd_net_),
            .in1(N__13089),
            .in2(_gnd_net_),
            .in3(N__13107),
            .lcout(),
            .ltout(\DUT.uart_inst0.un1_tx_clk_divider_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_RNITC2S1_0_LC_20_10_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNITC2S1_0_LC_20_10_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNITC2S1_0_LC_20_10_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNITC2S1_0_LC_20_10_2  (
            .in0(N__12454),
            .in1(N__12295),
            .in2(N__12448),
            .in3(N__12289),
            .lcout(\DUT.uart_inst0.un1_tx_clk_divider_0 ),
            .ltout(\DUT.uart_inst0.un1_tx_clk_divider_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNI5PJS2_1_LC_20_10_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNI5PJS2_1_LC_20_10_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNI5PJS2_1_LC_20_10_3 .LUT_INIT=16'b1111010111111111;
    LogicCell40 \DUT.uart_inst0.tx_state_RNI5PJS2_1_LC_20_10_3  (
            .in0(N__12283),
            .in1(_gnd_net_),
            .in2(N__12445),
            .in3(N__12438),
            .lcout(\DUT.uart_inst0.N_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_RNIQM95_0_LC_20_10_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNIQM95_0_LC_20_10_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNIQM95_0_LC_20_10_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNIQM95_0_LC_20_10_6  (
            .in0(N__12848),
            .in1(N__12612),
            .in2(N__12580),
            .in3(N__12594),
            .lcout(\DUT.uart_inst0.un1_tx_clk_divider_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_8_LC_20_10_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_8_LC_20_10_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_8_LC_20_10_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_8_LC_20_10_7  (
            .in0(N__13143),
            .in1(N__13158),
            .in2(N__13128),
            .in3(N__12492),
            .lcout(\DUT.uart_inst0.un1_tx_clk_divider_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNI9B9Q2_1_LC_20_11_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNI9B9Q2_1_LC_20_11_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNI9B9Q2_1_LC_20_11_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \DUT.uart_inst0.tx_state_RNI9B9Q2_1_LC_20_11_4  (
            .in0(_gnd_net_),
            .in1(N__12282),
            .in2(_gnd_net_),
            .in3(N__12196),
            .lcout(\DUT.uart_inst0.N_147 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_21_9_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_21_9_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_21_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_21_9_0  (
            .in0(_gnd_net_),
            .in1(N__12849),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_21_9_0_),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_1_LC_21_9_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_1_LC_21_9_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_1_LC_21_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_1_LC_21_9_1  (
            .in0(_gnd_net_),
            .in1(N__12613),
            .in2(N__13042),
            .in3(N__12601),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_1 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_0 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_1 ),
            .clk(N__12825),
            .ce(),
            .sr(N__12637));
    defparam \DUT.uart_inst0.tx_clk_divider_2_LC_21_9_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_2_LC_21_9_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_2_LC_21_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_2_LC_21_9_2  (
            .in0(_gnd_net_),
            .in1(N__13008),
            .in2(N__12598),
            .in3(N__12583),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_2 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_1 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_2 ),
            .clk(N__12825),
            .ce(),
            .sr(N__12637));
    defparam \DUT.uart_inst0.tx_clk_divider_3_LC_21_9_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_3_LC_21_9_3 .SEQ_MODE=4'b1001;
    defparam \DUT.uart_inst0.tx_clk_divider_3_LC_21_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_3_LC_21_9_3  (
            .in0(_gnd_net_),
            .in1(N__12579),
            .in2(N__13043),
            .in3(N__12565),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_3 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_2 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_3 ),
            .clk(N__12825),
            .ce(),
            .sr(N__12637));
    defparam \DUT.uart_inst0.tx_clk_divider_4_LC_21_9_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_4_LC_21_9_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_4_LC_21_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_4_LC_21_9_4  (
            .in0(_gnd_net_),
            .in1(N__13012),
            .in2(N__12562),
            .in3(N__12547),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_4 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_3 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_4 ),
            .clk(N__12825),
            .ce(),
            .sr(N__12637));
    defparam \DUT.uart_inst0.tx_clk_divider_5_LC_21_9_5 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_5_LC_21_9_5 .SEQ_MODE=4'b1001;
    defparam \DUT.uart_inst0.tx_clk_divider_5_LC_21_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_5_LC_21_9_5  (
            .in0(_gnd_net_),
            .in1(N__12544),
            .in2(N__13044),
            .in3(N__12532),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_5 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_4 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_5 ),
            .clk(N__12825),
            .ce(),
            .sr(N__12637));
    defparam \DUT.uart_inst0.tx_clk_divider_6_LC_21_9_6 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_6_LC_21_9_6 .SEQ_MODE=4'b1001;
    defparam \DUT.uart_inst0.tx_clk_divider_6_LC_21_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_6_LC_21_9_6  (
            .in0(_gnd_net_),
            .in1(N__13016),
            .in2(N__12529),
            .in3(N__12514),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_6 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_5 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_6 ),
            .clk(N__12825),
            .ce(),
            .sr(N__12637));
    defparam \DUT.uart_inst0.tx_clk_divider_7_LC_21_9_7 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_7_LC_21_9_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_7_LC_21_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_7_LC_21_9_7  (
            .in0(_gnd_net_),
            .in1(N__12510),
            .in2(N__13045),
            .in3(N__12496),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_7 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_6 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_7 ),
            .clk(N__12825),
            .ce(),
            .sr(N__12637));
    defparam \DUT.uart_inst0.tx_clk_divider_8_LC_21_10_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_8_LC_21_10_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_8_LC_21_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_8_LC_21_10_0  (
            .in0(_gnd_net_),
            .in1(N__12493),
            .in2(N__13004),
            .in3(N__12481),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_8 ),
            .ltout(),
            .carryin(bfn_21_10_0_),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_8 ),
            .clk(N__12821),
            .ce(),
            .sr(N__12636));
    defparam \DUT.uart_inst0.tx_clk_divider_9_LC_21_10_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_9_LC_21_10_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_9_LC_21_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_9_LC_21_10_1  (
            .in0(_gnd_net_),
            .in1(N__12972),
            .in2(N__13162),
            .in3(N__13147),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_9 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_8 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_9 ),
            .clk(N__12821),
            .ce(),
            .sr(N__12636));
    defparam \DUT.uart_inst0.tx_clk_divider_10_LC_21_10_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_10_LC_21_10_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_10_LC_21_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_10_LC_21_10_2  (
            .in0(_gnd_net_),
            .in1(N__13144),
            .in2(N__13002),
            .in3(N__13132),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_10 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_9 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_10 ),
            .clk(N__12821),
            .ce(),
            .sr(N__12636));
    defparam \DUT.uart_inst0.tx_clk_divider_11_LC_21_10_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_11_LC_21_10_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_11_LC_21_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_11_LC_21_10_3  (
            .in0(_gnd_net_),
            .in1(N__12965),
            .in2(N__13129),
            .in3(N__13111),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_11 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_10 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_11 ),
            .clk(N__12821),
            .ce(),
            .sr(N__12636));
    defparam \DUT.uart_inst0.tx_clk_divider_12_LC_21_10_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_12_LC_21_10_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_12_LC_21_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_12_LC_21_10_4  (
            .in0(_gnd_net_),
            .in1(N__13108),
            .in2(N__13003),
            .in3(N__13096),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_12 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_11 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_12 ),
            .clk(N__12821),
            .ce(),
            .sr(N__12636));
    defparam \DUT.uart_inst0.tx_clk_divider_13_LC_21_10_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_13_LC_21_10_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_13_LC_21_10_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_13_LC_21_10_5  (
            .in0(_gnd_net_),
            .in1(N__13090),
            .in2(_gnd_net_),
            .in3(N__13093),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12821),
            .ce(),
            .sr(N__12636));
    defparam \DUT.uart_inst0.tx_clk_divider_0_LC_21_10_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_0_LC_21_10_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_0_LC_21_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_0_LC_21_10_7  (
            .in0(_gnd_net_),
            .in1(N__12961),
            .in2(_gnd_net_),
            .in3(N__12850),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12821),
            .ce(),
            .sr(N__12636));
endmodule // top
