// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Mar 28 2020 19:39:19

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    ioFifoData,
    P1A9,
    P1A1,
    P1A8,
    oRx_n,
    P1A7,
    P1A3,
    iTxE_n,
    iRxF_n,
    iClk,
    P1A2,
    BTN_N,
    BTN1,
    oTx_n);

    output [7:0] ioFifoData;
    output P1A9;
    input P1A1;
    output P1A8;
    output oRx_n;
    output P1A7;
    output P1A3;
    input iTxE_n;
    input iRxF_n;
    input iClk;
    output P1A2;
    input BTN_N;
    input BTN1;
    output oTx_n;

    wire N__13213;
    wire N__13199;
    wire N__13198;
    wire N__13197;
    wire N__13190;
    wire N__13189;
    wire N__13188;
    wire N__13181;
    wire N__13180;
    wire N__13179;
    wire N__13172;
    wire N__13171;
    wire N__13170;
    wire N__13163;
    wire N__13162;
    wire N__13161;
    wire N__13154;
    wire N__13153;
    wire N__13152;
    wire N__13145;
    wire N__13144;
    wire N__13143;
    wire N__13136;
    wire N__13135;
    wire N__13134;
    wire N__13127;
    wire N__13126;
    wire N__13125;
    wire N__13118;
    wire N__13117;
    wire N__13116;
    wire N__13109;
    wire N__13108;
    wire N__13107;
    wire N__13100;
    wire N__13099;
    wire N__13098;
    wire N__13091;
    wire N__13090;
    wire N__13089;
    wire N__13082;
    wire N__13081;
    wire N__13080;
    wire N__13073;
    wire N__13072;
    wire N__13071;
    wire N__13064;
    wire N__13063;
    wire N__13062;
    wire N__13055;
    wire N__13054;
    wire N__13053;
    wire N__13046;
    wire N__13045;
    wire N__13044;
    wire N__13037;
    wire N__13036;
    wire N__13035;
    wire N__13018;
    wire N__13015;
    wire N__13012;
    wire N__13009;
    wire N__13008;
    wire N__13005;
    wire N__13002;
    wire N__13001;
    wire N__13000;
    wire N__12999;
    wire N__12998;
    wire N__12997;
    wire N__12996;
    wire N__12995;
    wire N__12994;
    wire N__12993;
    wire N__12992;
    wire N__12991;
    wire N__12990;
    wire N__12989;
    wire N__12988;
    wire N__12987;
    wire N__12986;
    wire N__12985;
    wire N__12984;
    wire N__12983;
    wire N__12982;
    wire N__12981;
    wire N__12980;
    wire N__12979;
    wire N__12978;
    wire N__12977;
    wire N__12972;
    wire N__12967;
    wire N__12960;
    wire N__12957;
    wire N__12954;
    wire N__12951;
    wire N__12948;
    wire N__12947;
    wire N__12944;
    wire N__12941;
    wire N__12938;
    wire N__12935;
    wire N__12932;
    wire N__12929;
    wire N__12926;
    wire N__12923;
    wire N__12920;
    wire N__12917;
    wire N__12914;
    wire N__12911;
    wire N__12908;
    wire N__12905;
    wire N__12902;
    wire N__12899;
    wire N__12898;
    wire N__12897;
    wire N__12896;
    wire N__12895;
    wire N__12894;
    wire N__12893;
    wire N__12892;
    wire N__12889;
    wire N__12884;
    wire N__12879;
    wire N__12868;
    wire N__12859;
    wire N__12850;
    wire N__12847;
    wire N__12842;
    wire N__12835;
    wire N__12832;
    wire N__12829;
    wire N__12826;
    wire N__12823;
    wire N__12820;
    wire N__12817;
    wire N__12814;
    wire N__12811;
    wire N__12808;
    wire N__12799;
    wire N__12792;
    wire N__12785;
    wire N__12776;
    wire N__12763;
    wire N__12762;
    wire N__12759;
    wire N__12756;
    wire N__12751;
    wire N__12748;
    wire N__12745;
    wire N__12744;
    wire N__12741;
    wire N__12738;
    wire N__12735;
    wire N__12730;
    wire N__12729;
    wire N__12726;
    wire N__12723;
    wire N__12720;
    wire N__12717;
    wire N__12716;
    wire N__12711;
    wire N__12708;
    wire N__12703;
    wire N__12700;
    wire N__12697;
    wire N__12694;
    wire N__12693;
    wire N__12690;
    wire N__12687;
    wire N__12682;
    wire N__12679;
    wire N__12676;
    wire N__12675;
    wire N__12674;
    wire N__12673;
    wire N__12672;
    wire N__12671;
    wire N__12670;
    wire N__12667;
    wire N__12666;
    wire N__12663;
    wire N__12662;
    wire N__12659;
    wire N__12656;
    wire N__12655;
    wire N__12654;
    wire N__12653;
    wire N__12650;
    wire N__12647;
    wire N__12646;
    wire N__12645;
    wire N__12642;
    wire N__12639;
    wire N__12636;
    wire N__12631;
    wire N__12628;
    wire N__12625;
    wire N__12620;
    wire N__12619;
    wire N__12618;
    wire N__12617;
    wire N__12616;
    wire N__12615;
    wire N__12614;
    wire N__12611;
    wire N__12608;
    wire N__12601;
    wire N__12592;
    wire N__12591;
    wire N__12584;
    wire N__12577;
    wire N__12570;
    wire N__12567;
    wire N__12560;
    wire N__12557;
    wire N__12554;
    wire N__12541;
    wire N__12540;
    wire N__12539;
    wire N__12536;
    wire N__12535;
    wire N__12534;
    wire N__12531;
    wire N__12530;
    wire N__12529;
    wire N__12528;
    wire N__12521;
    wire N__12518;
    wire N__12513;
    wire N__12508;
    wire N__12505;
    wire N__12502;
    wire N__12499;
    wire N__12496;
    wire N__12495;
    wire N__12494;
    wire N__12493;
    wire N__12492;
    wire N__12491;
    wire N__12490;
    wire N__12489;
    wire N__12488;
    wire N__12487;
    wire N__12486;
    wire N__12485;
    wire N__12484;
    wire N__12451;
    wire N__12448;
    wire N__12445;
    wire N__12444;
    wire N__12443;
    wire N__12442;
    wire N__12439;
    wire N__12436;
    wire N__12435;
    wire N__12432;
    wire N__12429;
    wire N__12426;
    wire N__12423;
    wire N__12420;
    wire N__12417;
    wire N__12406;
    wire N__12405;
    wire N__12404;
    wire N__12401;
    wire N__12400;
    wire N__12397;
    wire N__12396;
    wire N__12393;
    wire N__12390;
    wire N__12389;
    wire N__12388;
    wire N__12387;
    wire N__12384;
    wire N__12379;
    wire N__12376;
    wire N__12373;
    wire N__12370;
    wire N__12365;
    wire N__12352;
    wire N__12349;
    wire N__12346;
    wire N__12343;
    wire N__12340;
    wire N__12339;
    wire N__12338;
    wire N__12337;
    wire N__12334;
    wire N__12329;
    wire N__12328;
    wire N__12325;
    wire N__12324;
    wire N__12323;
    wire N__12322;
    wire N__12321;
    wire N__12320;
    wire N__12319;
    wire N__12318;
    wire N__12317;
    wire N__12312;
    wire N__12307;
    wire N__12304;
    wire N__12299;
    wire N__12296;
    wire N__12289;
    wire N__12286;
    wire N__12283;
    wire N__12278;
    wire N__12275;
    wire N__12270;
    wire N__12267;
    wire N__12266;
    wire N__12265;
    wire N__12262;
    wire N__12259;
    wire N__12256;
    wire N__12251;
    wire N__12246;
    wire N__12235;
    wire N__12234;
    wire N__12233;
    wire N__12230;
    wire N__12225;
    wire N__12224;
    wire N__12223;
    wire N__12218;
    wire N__12217;
    wire N__12216;
    wire N__12213;
    wire N__12210;
    wire N__12207;
    wire N__12204;
    wire N__12201;
    wire N__12190;
    wire N__12187;
    wire N__12184;
    wire N__12181;
    wire N__12178;
    wire N__12175;
    wire N__12172;
    wire N__12169;
    wire N__12166;
    wire N__12165;
    wire N__12164;
    wire N__12161;
    wire N__12158;
    wire N__12155;
    wire N__12152;
    wire N__12147;
    wire N__12142;
    wire N__12139;
    wire N__12138;
    wire N__12137;
    wire N__12136;
    wire N__12135;
    wire N__12134;
    wire N__12133;
    wire N__12132;
    wire N__12131;
    wire N__12130;
    wire N__12129;
    wire N__12128;
    wire N__12127;
    wire N__12126;
    wire N__12125;
    wire N__12124;
    wire N__12123;
    wire N__12122;
    wire N__12121;
    wire N__12120;
    wire N__12119;
    wire N__12118;
    wire N__12117;
    wire N__12116;
    wire N__12115;
    wire N__12114;
    wire N__12113;
    wire N__12112;
    wire N__12111;
    wire N__12110;
    wire N__12109;
    wire N__12108;
    wire N__12107;
    wire N__12106;
    wire N__12105;
    wire N__12104;
    wire N__12103;
    wire N__12102;
    wire N__12101;
    wire N__12100;
    wire N__12099;
    wire N__12098;
    wire N__12097;
    wire N__12096;
    wire N__12095;
    wire N__12094;
    wire N__12093;
    wire N__12092;
    wire N__12091;
    wire N__12090;
    wire N__12089;
    wire N__12088;
    wire N__12087;
    wire N__12086;
    wire N__12085;
    wire N__12084;
    wire N__12083;
    wire N__12082;
    wire N__12081;
    wire N__12080;
    wire N__12079;
    wire N__12078;
    wire N__12077;
    wire N__12076;
    wire N__12075;
    wire N__11944;
    wire N__11941;
    wire N__11940;
    wire N__11939;
    wire N__11938;
    wire N__11937;
    wire N__11936;
    wire N__11935;
    wire N__11932;
    wire N__11931;
    wire N__11930;
    wire N__11929;
    wire N__11926;
    wire N__11925;
    wire N__11924;
    wire N__11923;
    wire N__11922;
    wire N__11921;
    wire N__11920;
    wire N__11919;
    wire N__11918;
    wire N__11915;
    wire N__11908;
    wire N__11905;
    wire N__11898;
    wire N__11893;
    wire N__11890;
    wire N__11887;
    wire N__11884;
    wire N__11881;
    wire N__11878;
    wire N__11875;
    wire N__11872;
    wire N__11869;
    wire N__11868;
    wire N__11867;
    wire N__11866;
    wire N__11863;
    wire N__11862;
    wire N__11859;
    wire N__11856;
    wire N__11853;
    wire N__11850;
    wire N__11849;
    wire N__11848;
    wire N__11847;
    wire N__11846;
    wire N__11845;
    wire N__11844;
    wire N__11843;
    wire N__11840;
    wire N__11837;
    wire N__11836;
    wire N__11833;
    wire N__11832;
    wire N__11829;
    wire N__11826;
    wire N__11823;
    wire N__11820;
    wire N__11817;
    wire N__11764;
    wire N__11761;
    wire N__11758;
    wire N__11757;
    wire N__11754;
    wire N__11751;
    wire N__11748;
    wire N__11743;
    wire N__11740;
    wire N__11739;
    wire N__11736;
    wire N__11733;
    wire N__11728;
    wire N__11725;
    wire N__11724;
    wire N__11721;
    wire N__11718;
    wire N__11713;
    wire N__11710;
    wire N__11709;
    wire N__11706;
    wire N__11703;
    wire N__11698;
    wire N__11695;
    wire N__11694;
    wire N__11691;
    wire N__11688;
    wire N__11683;
    wire N__11680;
    wire N__11679;
    wire N__11676;
    wire N__11673;
    wire N__11668;
    wire N__11665;
    wire N__11664;
    wire N__11661;
    wire N__11658;
    wire N__11653;
    wire N__11650;
    wire N__11649;
    wire N__11646;
    wire N__11643;
    wire N__11640;
    wire N__11635;
    wire N__11632;
    wire N__11629;
    wire N__11626;
    wire N__11623;
    wire N__11622;
    wire N__11621;
    wire N__11620;
    wire N__11619;
    wire N__11618;
    wire N__11617;
    wire N__11614;
    wire N__11611;
    wire N__11610;
    wire N__11609;
    wire N__11608;
    wire N__11603;
    wire N__11602;
    wire N__11599;
    wire N__11596;
    wire N__11593;
    wire N__11590;
    wire N__11587;
    wire N__11586;
    wire N__11579;
    wire N__11576;
    wire N__11573;
    wire N__11566;
    wire N__11561;
    wire N__11558;
    wire N__11553;
    wire N__11542;
    wire N__11539;
    wire N__11536;
    wire N__11535;
    wire N__11532;
    wire N__11531;
    wire N__11528;
    wire N__11527;
    wire N__11526;
    wire N__11525;
    wire N__11524;
    wire N__11521;
    wire N__11520;
    wire N__11517;
    wire N__11512;
    wire N__11507;
    wire N__11506;
    wire N__11503;
    wire N__11502;
    wire N__11501;
    wire N__11498;
    wire N__11495;
    wire N__11494;
    wire N__11489;
    wire N__11486;
    wire N__11483;
    wire N__11478;
    wire N__11475;
    wire N__11472;
    wire N__11469;
    wire N__11466;
    wire N__11463;
    wire N__11460;
    wire N__11457;
    wire N__11454;
    wire N__11451;
    wire N__11448;
    wire N__11445;
    wire N__11442;
    wire N__11435;
    wire N__11430;
    wire N__11427;
    wire N__11424;
    wire N__11417;
    wire N__11412;
    wire N__11409;
    wire N__11404;
    wire N__11401;
    wire N__11400;
    wire N__11399;
    wire N__11398;
    wire N__11397;
    wire N__11396;
    wire N__11395;
    wire N__11394;
    wire N__11393;
    wire N__11392;
    wire N__11389;
    wire N__11388;
    wire N__11383;
    wire N__11380;
    wire N__11377;
    wire N__11376;
    wire N__11375;
    wire N__11372;
    wire N__11363;
    wire N__11360;
    wire N__11357;
    wire N__11352;
    wire N__11349;
    wire N__11344;
    wire N__11329;
    wire N__11328;
    wire N__11323;
    wire N__11322;
    wire N__11319;
    wire N__11316;
    wire N__11311;
    wire N__11308;
    wire N__11307;
    wire N__11304;
    wire N__11301;
    wire N__11296;
    wire N__11293;
    wire N__11292;
    wire N__11289;
    wire N__11286;
    wire N__11281;
    wire N__11278;
    wire N__11277;
    wire N__11276;
    wire N__11273;
    wire N__11270;
    wire N__11267;
    wire N__11262;
    wire N__11257;
    wire N__11254;
    wire N__11253;
    wire N__11250;
    wire N__11247;
    wire N__11244;
    wire N__11239;
    wire N__11236;
    wire N__11235;
    wire N__11232;
    wire N__11229;
    wire N__11226;
    wire N__11221;
    wire N__11218;
    wire N__11217;
    wire N__11214;
    wire N__11211;
    wire N__11206;
    wire N__11203;
    wire N__11202;
    wire N__11201;
    wire N__11200;
    wire N__11197;
    wire N__11196;
    wire N__11195;
    wire N__11194;
    wire N__11191;
    wire N__11182;
    wire N__11181;
    wire N__11180;
    wire N__11179;
    wire N__11178;
    wire N__11177;
    wire N__11176;
    wire N__11175;
    wire N__11174;
    wire N__11169;
    wire N__11164;
    wire N__11163;
    wire N__11162;
    wire N__11161;
    wire N__11160;
    wire N__11157;
    wire N__11156;
    wire N__11153;
    wire N__11150;
    wire N__11147;
    wire N__11146;
    wire N__11145;
    wire N__11138;
    wire N__11135;
    wire N__11132;
    wire N__11129;
    wire N__11114;
    wire N__11105;
    wire N__11102;
    wire N__11097;
    wire N__11086;
    wire N__11083;
    wire N__11082;
    wire N__11079;
    wire N__11076;
    wire N__11073;
    wire N__11068;
    wire N__11065;
    wire N__11062;
    wire N__11061;
    wire N__11058;
    wire N__11055;
    wire N__11052;
    wire N__11049;
    wire N__11044;
    wire N__11043;
    wire N__11040;
    wire N__11037;
    wire N__11036;
    wire N__11035;
    wire N__11034;
    wire N__11031;
    wire N__11026;
    wire N__11021;
    wire N__11014;
    wire N__11013;
    wire N__11012;
    wire N__11011;
    wire N__11006;
    wire N__11005;
    wire N__11000;
    wire N__10997;
    wire N__10994;
    wire N__10991;
    wire N__10988;
    wire N__10981;
    wire N__10978;
    wire N__10975;
    wire N__10972;
    wire N__10969;
    wire N__10966;
    wire N__10965;
    wire N__10964;
    wire N__10963;
    wire N__10960;
    wire N__10953;
    wire N__10948;
    wire N__10945;
    wire N__10942;
    wire N__10939;
    wire N__10936;
    wire N__10933;
    wire N__10932;
    wire N__10931;
    wire N__10928;
    wire N__10923;
    wire N__10918;
    wire N__10915;
    wire N__10912;
    wire N__10909;
    wire N__10906;
    wire N__10905;
    wire N__10904;
    wire N__10901;
    wire N__10900;
    wire N__10899;
    wire N__10898;
    wire N__10897;
    wire N__10896;
    wire N__10893;
    wire N__10890;
    wire N__10883;
    wire N__10878;
    wire N__10875;
    wire N__10872;
    wire N__10871;
    wire N__10870;
    wire N__10869;
    wire N__10864;
    wire N__10859;
    wire N__10856;
    wire N__10849;
    wire N__10846;
    wire N__10843;
    wire N__10840;
    wire N__10831;
    wire N__10830;
    wire N__10827;
    wire N__10824;
    wire N__10821;
    wire N__10818;
    wire N__10815;
    wire N__10812;
    wire N__10809;
    wire N__10804;
    wire N__10801;
    wire N__10798;
    wire N__10797;
    wire N__10796;
    wire N__10793;
    wire N__10790;
    wire N__10787;
    wire N__10780;
    wire N__10777;
    wire N__10774;
    wire N__10771;
    wire N__10770;
    wire N__10769;
    wire N__10766;
    wire N__10761;
    wire N__10756;
    wire N__10753;
    wire N__10750;
    wire N__10747;
    wire N__10746;
    wire N__10745;
    wire N__10742;
    wire N__10737;
    wire N__10732;
    wire N__10729;
    wire N__10726;
    wire N__10723;
    wire N__10722;
    wire N__10721;
    wire N__10718;
    wire N__10715;
    wire N__10710;
    wire N__10705;
    wire N__10702;
    wire N__10699;
    wire N__10696;
    wire N__10695;
    wire N__10694;
    wire N__10691;
    wire N__10686;
    wire N__10681;
    wire N__10678;
    wire N__10675;
    wire N__10672;
    wire N__10669;
    wire N__10668;
    wire N__10667;
    wire N__10664;
    wire N__10661;
    wire N__10658;
    wire N__10651;
    wire N__10648;
    wire N__10645;
    wire N__10642;
    wire N__10641;
    wire N__10640;
    wire N__10637;
    wire N__10632;
    wire N__10627;
    wire N__10624;
    wire N__10621;
    wire N__10618;
    wire N__10615;
    wire N__10614;
    wire N__10613;
    wire N__10610;
    wire N__10607;
    wire N__10604;
    wire N__10597;
    wire N__10594;
    wire N__10591;
    wire N__10588;
    wire N__10587;
    wire N__10586;
    wire N__10583;
    wire N__10580;
    wire N__10577;
    wire N__10570;
    wire N__10567;
    wire N__10564;
    wire N__10561;
    wire N__10558;
    wire N__10557;
    wire N__10556;
    wire N__10553;
    wire N__10548;
    wire N__10543;
    wire N__10540;
    wire N__10537;
    wire N__10534;
    wire N__10531;
    wire N__10530;
    wire N__10527;
    wire N__10526;
    wire N__10523;
    wire N__10520;
    wire N__10517;
    wire N__10514;
    wire N__10511;
    wire N__10508;
    wire N__10501;
    wire N__10498;
    wire N__10495;
    wire N__10492;
    wire N__10489;
    wire N__10486;
    wire N__10485;
    wire N__10484;
    wire N__10481;
    wire N__10478;
    wire N__10475;
    wire N__10472;
    wire N__10469;
    wire N__10462;
    wire N__10459;
    wire N__10456;
    wire N__10453;
    wire N__10452;
    wire N__10451;
    wire N__10448;
    wire N__10445;
    wire N__10442;
    wire N__10435;
    wire N__10432;
    wire N__10429;
    wire N__10426;
    wire N__10425;
    wire N__10424;
    wire N__10421;
    wire N__10418;
    wire N__10415;
    wire N__10408;
    wire N__10405;
    wire N__10402;
    wire N__10399;
    wire N__10398;
    wire N__10397;
    wire N__10394;
    wire N__10391;
    wire N__10388;
    wire N__10381;
    wire N__10378;
    wire N__10375;
    wire N__10372;
    wire N__10371;
    wire N__10368;
    wire N__10367;
    wire N__10364;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10352;
    wire N__10345;
    wire N__10342;
    wire N__10339;
    wire N__10336;
    wire N__10333;
    wire N__10332;
    wire N__10331;
    wire N__10328;
    wire N__10327;
    wire N__10324;
    wire N__10321;
    wire N__10318;
    wire N__10315;
    wire N__10312;
    wire N__10309;
    wire N__10306;
    wire N__10297;
    wire N__10294;
    wire N__10291;
    wire N__10288;
    wire N__10285;
    wire N__10282;
    wire N__10279;
    wire N__10276;
    wire N__10275;
    wire N__10272;
    wire N__10269;
    wire N__10268;
    wire N__10267;
    wire N__10262;
    wire N__10259;
    wire N__10256;
    wire N__10249;
    wire N__10246;
    wire N__10243;
    wire N__10240;
    wire N__10237;
    wire N__10234;
    wire N__10233;
    wire N__10230;
    wire N__10229;
    wire N__10226;
    wire N__10223;
    wire N__10220;
    wire N__10217;
    wire N__10212;
    wire N__10211;
    wire N__10208;
    wire N__10205;
    wire N__10202;
    wire N__10195;
    wire N__10192;
    wire N__10189;
    wire N__10186;
    wire N__10183;
    wire N__10180;
    wire N__10177;
    wire N__10174;
    wire N__10171;
    wire N__10168;
    wire N__10167;
    wire N__10164;
    wire N__10161;
    wire N__10158;
    wire N__10153;
    wire N__10152;
    wire N__10151;
    wire N__10148;
    wire N__10145;
    wire N__10142;
    wire N__10139;
    wire N__10132;
    wire N__10129;
    wire N__10126;
    wire N__10123;
    wire N__10120;
    wire N__10117;
    wire N__10116;
    wire N__10113;
    wire N__10110;
    wire N__10107;
    wire N__10104;
    wire N__10101;
    wire N__10096;
    wire N__10093;
    wire N__10090;
    wire N__10089;
    wire N__10086;
    wire N__10083;
    wire N__10080;
    wire N__10075;
    wire N__10074;
    wire N__10071;
    wire N__10068;
    wire N__10065;
    wire N__10062;
    wire N__10057;
    wire N__10054;
    wire N__10053;
    wire N__10052;
    wire N__10049;
    wire N__10044;
    wire N__10043;
    wire N__10042;
    wire N__10041;
    wire N__10036;
    wire N__10031;
    wire N__10030;
    wire N__10027;
    wire N__10026;
    wire N__10023;
    wire N__10020;
    wire N__10017;
    wire N__10014;
    wire N__10011;
    wire N__10000;
    wire N__9997;
    wire N__9994;
    wire N__9993;
    wire N__9992;
    wire N__9991;
    wire N__9990;
    wire N__9989;
    wire N__9988;
    wire N__9987;
    wire N__9986;
    wire N__9985;
    wire N__9984;
    wire N__9983;
    wire N__9982;
    wire N__9979;
    wire N__9976;
    wire N__9969;
    wire N__9968;
    wire N__9967;
    wire N__9966;
    wire N__9965;
    wire N__9964;
    wire N__9961;
    wire N__9956;
    wire N__9953;
    wire N__9944;
    wire N__9937;
    wire N__9932;
    wire N__9925;
    wire N__9910;
    wire N__9907;
    wire N__9904;
    wire N__9903;
    wire N__9900;
    wire N__9897;
    wire N__9894;
    wire N__9889;
    wire N__9886;
    wire N__9885;
    wire N__9882;
    wire N__9879;
    wire N__9874;
    wire N__9871;
    wire N__9870;
    wire N__9867;
    wire N__9864;
    wire N__9861;
    wire N__9856;
    wire N__9855;
    wire N__9852;
    wire N__9851;
    wire N__9850;
    wire N__9849;
    wire N__9846;
    wire N__9843;
    wire N__9842;
    wire N__9839;
    wire N__9838;
    wire N__9837;
    wire N__9834;
    wire N__9833;
    wire N__9832;
    wire N__9831;
    wire N__9828;
    wire N__9825;
    wire N__9822;
    wire N__9819;
    wire N__9816;
    wire N__9813;
    wire N__9804;
    wire N__9801;
    wire N__9784;
    wire N__9781;
    wire N__9778;
    wire N__9775;
    wire N__9772;
    wire N__9771;
    wire N__9768;
    wire N__9767;
    wire N__9766;
    wire N__9765;
    wire N__9764;
    wire N__9763;
    wire N__9760;
    wire N__9759;
    wire N__9756;
    wire N__9755;
    wire N__9754;
    wire N__9753;
    wire N__9748;
    wire N__9745;
    wire N__9742;
    wire N__9741;
    wire N__9740;
    wire N__9737;
    wire N__9734;
    wire N__9731;
    wire N__9728;
    wire N__9725;
    wire N__9720;
    wire N__9717;
    wire N__9708;
    wire N__9691;
    wire N__9688;
    wire N__9685;
    wire N__9682;
    wire N__9679;
    wire N__9676;
    wire N__9675;
    wire N__9674;
    wire N__9673;
    wire N__9672;
    wire N__9671;
    wire N__9670;
    wire N__9667;
    wire N__9664;
    wire N__9661;
    wire N__9660;
    wire N__9659;
    wire N__9658;
    wire N__9657;
    wire N__9656;
    wire N__9653;
    wire N__9652;
    wire N__9651;
    wire N__9650;
    wire N__9649;
    wire N__9648;
    wire N__9647;
    wire N__9644;
    wire N__9643;
    wire N__9642;
    wire N__9639;
    wire N__9636;
    wire N__9631;
    wire N__9628;
    wire N__9621;
    wire N__9612;
    wire N__9599;
    wire N__9590;
    wire N__9577;
    wire N__9574;
    wire N__9571;
    wire N__9568;
    wire N__9565;
    wire N__9562;
    wire N__9559;
    wire N__9556;
    wire N__9553;
    wire N__9550;
    wire N__9547;
    wire N__9544;
    wire N__9541;
    wire N__9538;
    wire N__9535;
    wire N__9532;
    wire N__9529;
    wire N__9526;
    wire N__9523;
    wire N__9522;
    wire N__9521;
    wire N__9518;
    wire N__9517;
    wire N__9514;
    wire N__9513;
    wire N__9510;
    wire N__9509;
    wire N__9506;
    wire N__9505;
    wire N__9504;
    wire N__9503;
    wire N__9500;
    wire N__9497;
    wire N__9490;
    wire N__9487;
    wire N__9484;
    wire N__9481;
    wire N__9476;
    wire N__9463;
    wire N__9462;
    wire N__9461;
    wire N__9458;
    wire N__9457;
    wire N__9456;
    wire N__9453;
    wire N__9452;
    wire N__9451;
    wire N__9446;
    wire N__9443;
    wire N__9440;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9422;
    wire N__9409;
    wire N__9406;
    wire N__9405;
    wire N__9404;
    wire N__9403;
    wire N__9402;
    wire N__9401;
    wire N__9400;
    wire N__9399;
    wire N__9396;
    wire N__9387;
    wire N__9386;
    wire N__9385;
    wire N__9382;
    wire N__9379;
    wire N__9376;
    wire N__9373;
    wire N__9370;
    wire N__9365;
    wire N__9352;
    wire N__9349;
    wire N__9348;
    wire N__9347;
    wire N__9344;
    wire N__9343;
    wire N__9340;
    wire N__9339;
    wire N__9336;
    wire N__9335;
    wire N__9334;
    wire N__9333;
    wire N__9330;
    wire N__9327;
    wire N__9324;
    wire N__9321;
    wire N__9318;
    wire N__9311;
    wire N__9308;
    wire N__9295;
    wire N__9292;
    wire N__9291;
    wire N__9288;
    wire N__9285;
    wire N__9282;
    wire N__9277;
    wire N__9274;
    wire N__9271;
    wire N__9268;
    wire N__9265;
    wire N__9264;
    wire N__9261;
    wire N__9258;
    wire N__9253;
    wire N__9250;
    wire N__9249;
    wire N__9246;
    wire N__9243;
    wire N__9240;
    wire N__9235;
    wire N__9232;
    wire N__9229;
    wire N__9228;
    wire N__9225;
    wire N__9222;
    wire N__9217;
    wire N__9214;
    wire N__9211;
    wire N__9208;
    wire N__9207;
    wire N__9202;
    wire N__9199;
    wire N__9196;
    wire N__9193;
    wire N__9192;
    wire N__9189;
    wire N__9186;
    wire N__9181;
    wire N__9180;
    wire N__9177;
    wire N__9174;
    wire N__9169;
    wire N__9166;
    wire N__9165;
    wire N__9162;
    wire N__9161;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9145;
    wire N__9144;
    wire N__9143;
    wire N__9142;
    wire N__9137;
    wire N__9132;
    wire N__9131;
    wire N__9130;
    wire N__9129;
    wire N__9128;
    wire N__9127;
    wire N__9124;
    wire N__9121;
    wire N__9116;
    wire N__9111;
    wire N__9108;
    wire N__9097;
    wire N__9094;
    wire N__9093;
    wire N__9092;
    wire N__9087;
    wire N__9084;
    wire N__9081;
    wire N__9078;
    wire N__9075;
    wire N__9070;
    wire N__9069;
    wire N__9068;
    wire N__9063;
    wire N__9062;
    wire N__9059;
    wire N__9056;
    wire N__9053;
    wire N__9046;
    wire N__9045;
    wire N__9042;
    wire N__9039;
    wire N__9034;
    wire N__9031;
    wire N__9030;
    wire N__9027;
    wire N__9024;
    wire N__9019;
    wire N__9016;
    wire N__9013;
    wire N__9010;
    wire N__9007;
    wire N__9006;
    wire N__9003;
    wire N__9000;
    wire N__8997;
    wire N__8992;
    wire N__8991;
    wire N__8988;
    wire N__8985;
    wire N__8984;
    wire N__8983;
    wire N__8978;
    wire N__8975;
    wire N__8972;
    wire N__8967;
    wire N__8964;
    wire N__8961;
    wire N__8958;
    wire N__8955;
    wire N__8952;
    wire N__8947;
    wire N__8944;
    wire N__8941;
    wire N__8938;
    wire N__8937;
    wire N__8934;
    wire N__8933;
    wire N__8930;
    wire N__8929;
    wire N__8926;
    wire N__8923;
    wire N__8920;
    wire N__8917;
    wire N__8914;
    wire N__8911;
    wire N__8906;
    wire N__8903;
    wire N__8900;
    wire N__8897;
    wire N__8890;
    wire N__8887;
    wire N__8884;
    wire N__8881;
    wire N__8878;
    wire N__8877;
    wire N__8876;
    wire N__8873;
    wire N__8870;
    wire N__8867;
    wire N__8866;
    wire N__8863;
    wire N__8858;
    wire N__8855;
    wire N__8852;
    wire N__8847;
    wire N__8844;
    wire N__8841;
    wire N__8836;
    wire N__8833;
    wire N__8830;
    wire N__8827;
    wire N__8824;
    wire N__8821;
    wire N__8818;
    wire N__8815;
    wire N__8812;
    wire N__8809;
    wire N__8806;
    wire N__8803;
    wire N__8800;
    wire N__8797;
    wire N__8796;
    wire N__8793;
    wire N__8790;
    wire N__8787;
    wire N__8784;
    wire N__8779;
    wire N__8776;
    wire N__8773;
    wire N__8770;
    wire N__8767;
    wire N__8764;
    wire N__8761;
    wire N__8758;
    wire N__8755;
    wire N__8752;
    wire N__8749;
    wire N__8746;
    wire N__8743;
    wire N__8740;
    wire N__8739;
    wire N__8736;
    wire N__8733;
    wire N__8728;
    wire N__8725;
    wire N__8722;
    wire N__8719;
    wire N__8718;
    wire N__8715;
    wire N__8712;
    wire N__8707;
    wire N__8704;
    wire N__8701;
    wire N__8698;
    wire N__8695;
    wire N__8692;
    wire N__8689;
    wire N__8686;
    wire N__8683;
    wire N__8682;
    wire N__8681;
    wire N__8680;
    wire N__8677;
    wire N__8676;
    wire N__8675;
    wire N__8674;
    wire N__8673;
    wire N__8670;
    wire N__8667;
    wire N__8664;
    wire N__8661;
    wire N__8658;
    wire N__8651;
    wire N__8648;
    wire N__8643;
    wire N__8636;
    wire N__8629;
    wire N__8626;
    wire N__8623;
    wire N__8622;
    wire N__8621;
    wire N__8620;
    wire N__8617;
    wire N__8614;
    wire N__8609;
    wire N__8602;
    wire N__8599;
    wire N__8596;
    wire N__8593;
    wire N__8590;
    wire N__8587;
    wire N__8584;
    wire N__8581;
    wire N__8578;
    wire N__8577;
    wire N__8576;
    wire N__8575;
    wire N__8570;
    wire N__8565;
    wire N__8562;
    wire N__8559;
    wire N__8554;
    wire N__8551;
    wire N__8548;
    wire N__8545;
    wire N__8544;
    wire N__8541;
    wire N__8540;
    wire N__8537;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8521;
    wire N__8518;
    wire N__8515;
    wire N__8512;
    wire N__8509;
    wire N__8508;
    wire N__8505;
    wire N__8504;
    wire N__8501;
    wire N__8498;
    wire N__8495;
    wire N__8492;
    wire N__8485;
    wire N__8482;
    wire N__8479;
    wire N__8476;
    wire N__8475;
    wire N__8472;
    wire N__8469;
    wire N__8464;
    wire N__8463;
    wire N__8460;
    wire N__8459;
    wire N__8456;
    wire N__8451;
    wire N__8448;
    wire N__8443;
    wire N__8440;
    wire N__8437;
    wire N__8434;
    wire N__8431;
    wire N__8430;
    wire N__8427;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8419;
    wire N__8418;
    wire N__8417;
    wire N__8416;
    wire N__8415;
    wire N__8412;
    wire N__8409;
    wire N__8406;
    wire N__8401;
    wire N__8394;
    wire N__8383;
    wire N__8380;
    wire N__8377;
    wire N__8374;
    wire N__8371;
    wire N__8370;
    wire N__8369;
    wire N__8368;
    wire N__8367;
    wire N__8366;
    wire N__8363;
    wire N__8360;
    wire N__8359;
    wire N__8356;
    wire N__8355;
    wire N__8352;
    wire N__8349;
    wire N__8346;
    wire N__8343;
    wire N__8340;
    wire N__8337;
    wire N__8332;
    wire N__8327;
    wire N__8314;
    wire N__8313;
    wire N__8310;
    wire N__8307;
    wire N__8304;
    wire N__8301;
    wire N__8296;
    wire N__8293;
    wire N__8292;
    wire N__8291;
    wire N__8290;
    wire N__8289;
    wire N__8288;
    wire N__8285;
    wire N__8280;
    wire N__8275;
    wire N__8270;
    wire N__8263;
    wire N__8262;
    wire N__8261;
    wire N__8258;
    wire N__8255;
    wire N__8252;
    wire N__8249;
    wire N__8242;
    wire N__8241;
    wire N__8240;
    wire N__8239;
    wire N__8238;
    wire N__8233;
    wire N__8230;
    wire N__8229;
    wire N__8228;
    wire N__8225;
    wire N__8224;
    wire N__8223;
    wire N__8220;
    wire N__8217;
    wire N__8214;
    wire N__8211;
    wire N__8206;
    wire N__8203;
    wire N__8200;
    wire N__8197;
    wire N__8184;
    wire N__8183;
    wire N__8180;
    wire N__8177;
    wire N__8174;
    wire N__8167;
    wire N__8164;
    wire N__8161;
    wire N__8158;
    wire N__8157;
    wire N__8156;
    wire N__8155;
    wire N__8154;
    wire N__8153;
    wire N__8152;
    wire N__8151;
    wire N__8150;
    wire N__8147;
    wire N__8142;
    wire N__8139;
    wire N__8132;
    wire N__8127;
    wire N__8116;
    wire N__8113;
    wire N__8110;
    wire N__8107;
    wire N__8104;
    wire N__8103;
    wire N__8100;
    wire N__8097;
    wire N__8092;
    wire N__8089;
    wire N__8086;
    wire N__8083;
    wire N__8080;
    wire N__8079;
    wire N__8074;
    wire N__8071;
    wire N__8068;
    wire N__8065;
    wire N__8062;
    wire N__8059;
    wire N__8056;
    wire N__8053;
    wire N__8050;
    wire N__8047;
    wire N__8044;
    wire N__8041;
    wire N__8040;
    wire N__8039;
    wire N__8038;
    wire N__8031;
    wire N__8028;
    wire N__8023;
    wire N__8020;
    wire N__8017;
    wire N__8014;
    wire N__8013;
    wire N__8012;
    wire N__8011;
    wire N__8010;
    wire N__8009;
    wire N__8008;
    wire N__8007;
    wire N__8004;
    wire N__8001;
    wire N__7998;
    wire N__7993;
    wire N__7986;
    wire N__7975;
    wire N__7972;
    wire N__7969;
    wire N__7966;
    wire N__7965;
    wire N__7962;
    wire N__7959;
    wire N__7954;
    wire N__7951;
    wire N__7948;
    wire N__7945;
    wire N__7944;
    wire N__7941;
    wire N__7938;
    wire N__7937;
    wire N__7936;
    wire N__7933;
    wire N__7930;
    wire N__7927;
    wire N__7924;
    wire N__7915;
    wire N__7912;
    wire N__7909;
    wire N__7906;
    wire N__7903;
    wire N__7900;
    wire N__7897;
    wire N__7896;
    wire N__7893;
    wire N__7890;
    wire N__7885;
    wire N__7882;
    wire N__7879;
    wire N__7876;
    wire N__7873;
    wire N__7870;
    wire N__7869;
    wire N__7868;
    wire N__7865;
    wire N__7860;
    wire N__7855;
    wire N__7852;
    wire N__7849;
    wire N__7848;
    wire N__7847;
    wire N__7844;
    wire N__7839;
    wire N__7834;
    wire N__7833;
    wire N__7832;
    wire N__7829;
    wire N__7824;
    wire N__7819;
    wire N__7816;
    wire N__7813;
    wire N__7812;
    wire N__7811;
    wire N__7810;
    wire N__7807;
    wire N__7800;
    wire N__7795;
    wire N__7792;
    wire N__7789;
    wire N__7786;
    wire N__7783;
    wire N__7780;
    wire N__7777;
    wire N__7774;
    wire N__7771;
    wire N__7768;
    wire N__7767;
    wire N__7766;
    wire N__7763;
    wire N__7760;
    wire N__7757;
    wire N__7756;
    wire N__7751;
    wire N__7748;
    wire N__7745;
    wire N__7742;
    wire N__7737;
    wire N__7734;
    wire N__7731;
    wire N__7726;
    wire N__7723;
    wire N__7720;
    wire N__7717;
    wire N__7716;
    wire N__7715;
    wire N__7712;
    wire N__7709;
    wire N__7706;
    wire N__7705;
    wire N__7702;
    wire N__7697;
    wire N__7694;
    wire N__7691;
    wire N__7686;
    wire N__7683;
    wire N__7680;
    wire N__7675;
    wire N__7672;
    wire N__7669;
    wire N__7666;
    wire N__7663;
    wire N__7662;
    wire N__7661;
    wire N__7660;
    wire N__7657;
    wire N__7654;
    wire N__7651;
    wire N__7648;
    wire N__7639;
    wire N__7636;
    wire N__7633;
    wire N__7630;
    wire N__7627;
    wire N__7624;
    wire N__7621;
    wire N__7620;
    wire N__7619;
    wire N__7616;
    wire N__7613;
    wire N__7612;
    wire N__7611;
    wire N__7610;
    wire N__7609;
    wire N__7608;
    wire N__7605;
    wire N__7602;
    wire N__7599;
    wire N__7596;
    wire N__7591;
    wire N__7588;
    wire N__7585;
    wire N__7582;
    wire N__7575;
    wire N__7574;
    wire N__7569;
    wire N__7564;
    wire N__7561;
    wire N__7558;
    wire N__7549;
    wire N__7548;
    wire N__7547;
    wire N__7546;
    wire N__7545;
    wire N__7542;
    wire N__7541;
    wire N__7538;
    wire N__7535;
    wire N__7532;
    wire N__7529;
    wire N__7528;
    wire N__7525;
    wire N__7522;
    wire N__7519;
    wire N__7514;
    wire N__7511;
    wire N__7508;
    wire N__7505;
    wire N__7504;
    wire N__7503;
    wire N__7502;
    wire N__7497;
    wire N__7488;
    wire N__7481;
    wire N__7474;
    wire N__7473;
    wire N__7472;
    wire N__7471;
    wire N__7470;
    wire N__7467;
    wire N__7464;
    wire N__7457;
    wire N__7450;
    wire N__7447;
    wire N__7444;
    wire N__7441;
    wire N__7438;
    wire N__7435;
    wire N__7432;
    wire N__7429;
    wire N__7426;
    wire N__7423;
    wire N__7420;
    wire N__7417;
    wire N__7414;
    wire N__7411;
    wire N__7408;
    wire N__7405;
    wire N__7402;
    wire N__7399;
    wire N__7396;
    wire N__7393;
    wire N__7392;
    wire N__7391;
    wire N__7390;
    wire N__7387;
    wire N__7386;
    wire N__7385;
    wire N__7384;
    wire N__7383;
    wire N__7382;
    wire N__7381;
    wire N__7380;
    wire N__7377;
    wire N__7374;
    wire N__7367;
    wire N__7362;
    wire N__7353;
    wire N__7342;
    wire N__7339;
    wire N__7336;
    wire N__7333;
    wire N__7330;
    wire N__7327;
    wire N__7324;
    wire N__7321;
    wire N__7318;
    wire N__7315;
    wire N__7312;
    wire N__7311;
    wire N__7308;
    wire N__7305;
    wire N__7302;
    wire N__7297;
    wire N__7294;
    wire N__7293;
    wire N__7292;
    wire N__7291;
    wire N__7290;
    wire N__7281;
    wire N__7278;
    wire N__7273;
    wire N__7270;
    wire N__7267;
    wire N__7264;
    wire N__7263;
    wire N__7258;
    wire N__7255;
    wire N__7252;
    wire N__7249;
    wire N__7246;
    wire N__7243;
    wire N__7240;
    wire N__7237;
    wire N__7234;
    wire N__7233;
    wire N__7230;
    wire N__7227;
    wire N__7224;
    wire N__7221;
    wire N__7216;
    wire N__7213;
    wire N__7210;
    wire N__7207;
    wire N__7206;
    wire N__7203;
    wire N__7200;
    wire N__7195;
    wire N__7194;
    wire N__7193;
    wire N__7190;
    wire N__7187;
    wire N__7184;
    wire N__7177;
    wire N__7176;
    wire N__7173;
    wire N__7170;
    wire N__7169;
    wire N__7166;
    wire N__7161;
    wire N__7156;
    wire N__7153;
    wire N__7152;
    wire N__7149;
    wire N__7146;
    wire N__7143;
    wire N__7138;
    wire N__7137;
    wire N__7136;
    wire N__7135;
    wire N__7132;
    wire N__7127;
    wire N__7124;
    wire N__7119;
    wire N__7114;
    wire N__7111;
    wire N__7108;
    wire N__7105;
    wire N__7102;
    wire N__7101;
    wire N__7100;
    wire N__7097;
    wire N__7094;
    wire N__7093;
    wire N__7092;
    wire N__7091;
    wire N__7088;
    wire N__7085;
    wire N__7082;
    wire N__7079;
    wire N__7074;
    wire N__7063;
    wire N__7060;
    wire N__7057;
    wire N__7054;
    wire N__7051;
    wire N__7048;
    wire N__7045;
    wire N__7042;
    wire N__7039;
    wire N__7036;
    wire N__7033;
    wire N__7032;
    wire N__7031;
    wire N__7028;
    wire N__7025;
    wire N__7024;
    wire N__7021;
    wire N__7016;
    wire N__7013;
    wire N__7006;
    wire N__7003;
    wire N__7002;
    wire N__7001;
    wire N__6998;
    wire N__6995;
    wire N__6994;
    wire N__6993;
    wire N__6990;
    wire N__6985;
    wire N__6982;
    wire N__6979;
    wire N__6970;
    wire N__6967;
    wire N__6966;
    wire N__6965;
    wire N__6962;
    wire N__6959;
    wire N__6956;
    wire N__6955;
    wire N__6954;
    wire N__6951;
    wire N__6946;
    wire N__6943;
    wire N__6940;
    wire N__6931;
    wire N__6930;
    wire N__6927;
    wire N__6924;
    wire N__6923;
    wire N__6920;
    wire N__6917;
    wire N__6914;
    wire N__6913;
    wire N__6912;
    wire N__6909;
    wire N__6904;
    wire N__6901;
    wire N__6898;
    wire N__6889;
    wire N__6888;
    wire N__6885;
    wire N__6882;
    wire N__6881;
    wire N__6878;
    wire N__6875;
    wire N__6872;
    wire N__6871;
    wire N__6870;
    wire N__6863;
    wire N__6860;
    wire N__6857;
    wire N__6850;
    wire N__6849;
    wire N__6846;
    wire N__6843;
    wire N__6842;
    wire N__6839;
    wire N__6836;
    wire N__6833;
    wire N__6832;
    wire N__6831;
    wire N__6824;
    wire N__6821;
    wire N__6818;
    wire N__6811;
    wire N__6810;
    wire N__6807;
    wire N__6804;
    wire N__6803;
    wire N__6800;
    wire N__6797;
    wire N__6794;
    wire N__6793;
    wire N__6792;
    wire N__6785;
    wire N__6782;
    wire N__6779;
    wire N__6772;
    wire N__6769;
    wire N__6768;
    wire N__6765;
    wire N__6764;
    wire N__6761;
    wire N__6760;
    wire N__6759;
    wire N__6756;
    wire N__6753;
    wire N__6750;
    wire N__6747;
    wire N__6744;
    wire N__6733;
    wire N__6730;
    wire N__6729;
    wire N__6726;
    wire N__6725;
    wire N__6722;
    wire N__6721;
    wire N__6720;
    wire N__6715;
    wire N__6708;
    wire N__6703;
    wire N__6700;
    wire N__6697;
    wire N__6694;
    wire N__6693;
    wire N__6692;
    wire N__6691;
    wire N__6684;
    wire N__6681;
    wire N__6676;
    wire N__6675;
    wire N__6674;
    wire N__6667;
    wire N__6664;
    wire N__6661;
    wire N__6658;
    wire N__6655;
    wire N__6652;
    wire N__6649;
    wire N__6646;
    wire N__6643;
    wire N__6640;
    wire N__6637;
    wire N__6634;
    wire N__6631;
    wire N__6628;
    wire N__6625;
    wire N__6622;
    wire N__6619;
    wire N__6616;
    wire N__6613;
    wire N__6610;
    wire N__6607;
    wire N__6604;
    wire N__6601;
    wire N__6598;
    wire N__6595;
    wire N__6592;
    wire N__6589;
    wire N__6586;
    wire N__6583;
    wire N__6580;
    wire N__6579;
    wire N__6576;
    wire N__6573;
    wire N__6568;
    wire N__6565;
    wire N__6564;
    wire N__6559;
    wire N__6556;
    wire N__6553;
    wire N__6552;
    wire N__6551;
    wire N__6550;
    wire N__6549;
    wire N__6542;
    wire N__6539;
    wire N__6536;
    wire N__6529;
    wire N__6526;
    wire N__6523;
    wire N__6520;
    wire N__6517;
    wire N__6516;
    wire N__6515;
    wire N__6512;
    wire N__6509;
    wire N__6506;
    wire N__6499;
    wire N__6498;
    wire N__6497;
    wire N__6496;
    wire N__6493;
    wire N__6484;
    wire N__6481;
    wire N__6480;
    wire N__6479;
    wire N__6474;
    wire N__6471;
    wire N__6466;
    wire N__6463;
    wire N__6460;
    wire N__6457;
    wire N__6454;
    wire N__6451;
    wire N__6448;
    wire N__6445;
    wire N__6442;
    wire N__6439;
    wire N__6436;
    wire N__6433;
    wire N__6430;
    wire N__6427;
    wire N__6424;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire N__6414;
    wire N__6413;
    wire N__6412;
    wire N__6411;
    wire N__6410;
    wire N__6409;
    wire N__6408;
    wire N__6407;
    wire N__6404;
    wire N__6401;
    wire N__6400;
    wire N__6393;
    wire N__6392;
    wire N__6389;
    wire N__6386;
    wire N__6381;
    wire N__6378;
    wire N__6375;
    wire N__6372;
    wire N__6369;
    wire N__6366;
    wire N__6349;
    wire N__6346;
    wire N__6343;
    wire N__6340;
    wire N__6337;
    wire N__6334;
    wire N__6331;
    wire N__6328;
    wire N__6325;
    wire N__6322;
    wire N__6319;
    wire N__6316;
    wire N__6313;
    wire N__6310;
    wire N__6307;
    wire N__6304;
    wire N__6303;
    wire N__6300;
    wire N__6297;
    wire N__6292;
    wire N__6291;
    wire N__6288;
    wire N__6285;
    wire N__6280;
    wire N__6277;
    wire N__6274;
    wire N__6271;
    wire N__6268;
    wire N__6265;
    wire N__6262;
    wire N__6259;
    wire N__6256;
    wire N__6253;
    wire N__6250;
    wire N__6247;
    wire N__6244;
    wire N__6241;
    wire N__6238;
    wire N__6235;
    wire N__6232;
    wire N__6229;
    wire N__6226;
    wire N__6223;
    wire N__6220;
    wire N__6217;
    wire N__6214;
    wire N__6211;
    wire N__6208;
    wire N__6205;
    wire N__6204;
    wire N__6201;
    wire N__6198;
    wire N__6193;
    wire N__6192;
    wire N__6189;
    wire N__6186;
    wire N__6181;
    wire N__6178;
    wire N__6175;
    wire N__6172;
    wire N__6169;
    wire N__6166;
    wire N__6165;
    wire N__6162;
    wire N__6159;
    wire N__6154;
    wire N__6153;
    wire N__6150;
    wire N__6147;
    wire N__6146;
    wire N__6145;
    wire N__6144;
    wire N__6139;
    wire N__6132;
    wire N__6127;
    wire N__6124;
    wire N__6121;
    wire N__6118;
    wire N__6115;
    wire N__6114;
    wire N__6111;
    wire N__6108;
    wire N__6105;
    wire N__6102;
    wire N__6097;
    wire N__6094;
    wire N__6093;
    wire N__6088;
    wire N__6085;
    wire N__6084;
    wire N__6079;
    wire N__6076;
    wire N__6073;
    wire N__6070;
    wire N__6067;
    wire N__6066;
    wire N__6063;
    wire N__6062;
    wire N__6059;
    wire N__6058;
    wire N__6055;
    wire N__6050;
    wire N__6047;
    wire N__6040;
    wire N__6037;
    wire N__6036;
    wire N__6033;
    wire N__6030;
    wire N__6025;
    wire N__6024;
    wire N__6021;
    wire N__6018;
    wire N__6013;
    wire N__6012;
    wire N__6011;
    wire N__6010;
    wire N__6009;
    wire N__6008;
    wire N__6007;
    wire N__6004;
    wire N__6003;
    wire N__6002;
    wire N__6001;
    wire N__6000;
    wire N__5999;
    wire N__5998;
    wire N__5997;
    wire N__5996;
    wire N__5995;
    wire N__5994;
    wire N__5993;
    wire N__5976;
    wire N__5975;
    wire N__5974;
    wire N__5971;
    wire N__5968;
    wire N__5951;
    wire N__5948;
    wire N__5941;
    wire N__5938;
    wire N__5929;
    wire N__5926;
    wire N__5923;
    wire N__5920;
    wire N__5919;
    wire N__5918;
    wire N__5911;
    wire N__5908;
    wire N__5905;
    wire N__5904;
    wire N__5903;
    wire N__5902;
    wire N__5901;
    wire N__5900;
    wire N__5899;
    wire N__5898;
    wire N__5889;
    wire N__5888;
    wire N__5887;
    wire N__5886;
    wire N__5885;
    wire N__5884;
    wire N__5875;
    wire N__5872;
    wire N__5863;
    wire N__5860;
    wire N__5851;
    wire N__5848;
    wire N__5847;
    wire N__5844;
    wire N__5841;
    wire N__5836;
    wire N__5833;
    wire N__5832;
    wire N__5831;
    wire N__5828;
    wire N__5825;
    wire N__5824;
    wire N__5823;
    wire N__5820;
    wire N__5817;
    wire N__5814;
    wire N__5809;
    wire N__5800;
    wire N__5797;
    wire N__5794;
    wire N__5793;
    wire N__5790;
    wire N__5787;
    wire N__5782;
    wire N__5781;
    wire N__5778;
    wire N__5775;
    wire N__5770;
    wire N__5767;
    wire N__5764;
    wire N__5761;
    wire N__5758;
    wire N__5755;
    wire N__5752;
    wire N__5749;
    wire N__5746;
    wire N__5743;
    wire N__5740;
    wire N__5737;
    wire N__5734;
    wire N__5731;
    wire N__5728;
    wire N__5725;
    wire N__5722;
    wire N__5719;
    wire N__5716;
    wire N__5713;
    wire N__5710;
    wire N__5707;
    wire N__5706;
    wire N__5703;
    wire N__5700;
    wire N__5697;
    wire N__5694;
    wire N__5689;
    wire N__5688;
    wire N__5685;
    wire N__5682;
    wire N__5677;
    wire N__5674;
    wire N__5671;
    wire N__5670;
    wire N__5667;
    wire N__5664;
    wire N__5663;
    wire N__5660;
    wire N__5657;
    wire N__5654;
    wire N__5651;
    wire N__5650;
    wire N__5647;
    wire N__5642;
    wire N__5639;
    wire N__5632;
    wire N__5629;
    wire N__5626;
    wire N__5623;
    wire N__5620;
    wire N__5617;
    wire N__5614;
    wire N__5611;
    wire N__5608;
    wire N__5605;
    wire N__5602;
    wire N__5599;
    wire N__5596;
    wire N__5593;
    wire N__5590;
    wire N__5587;
    wire N__5584;
    wire N__5581;
    wire N__5578;
    wire N__5575;
    wire N__5572;
    wire N__5569;
    wire N__5566;
    wire N__5563;
    wire N__5560;
    wire N__5557;
    wire N__5556;
    wire N__5555;
    wire N__5552;
    wire N__5549;
    wire N__5548;
    wire N__5547;
    wire N__5546;
    wire N__5545;
    wire N__5542;
    wire N__5537;
    wire N__5528;
    wire N__5521;
    wire N__5520;
    wire N__5519;
    wire N__5518;
    wire N__5515;
    wire N__5514;
    wire N__5511;
    wire N__5508;
    wire N__5501;
    wire N__5494;
    wire N__5491;
    wire N__5490;
    wire N__5485;
    wire N__5482;
    wire N__5481;
    wire N__5476;
    wire N__5473;
    wire N__5472;
    wire N__5471;
    wire N__5470;
    wire N__5465;
    wire N__5460;
    wire N__5455;
    wire N__5454;
    wire N__5453;
    wire N__5452;
    wire N__5451;
    wire N__5450;
    wire N__5447;
    wire N__5440;
    wire N__5433;
    wire N__5428;
    wire N__5425;
    wire N__5424;
    wire N__5423;
    wire N__5422;
    wire N__5419;
    wire N__5418;
    wire N__5411;
    wire N__5406;
    wire N__5401;
    wire N__5398;
    wire N__5395;
    wire N__5392;
    wire N__5389;
    wire N__5386;
    wire N__5383;
    wire N__5380;
    wire N__5377;
    wire N__5374;
    wire N__5371;
    wire N__5368;
    wire N__5365;
    wire N__5362;
    wire N__5359;
    wire N__5356;
    wire N__5353;
    wire N__5350;
    wire N__5347;
    wire N__5344;
    wire N__5341;
    wire N__5338;
    wire N__5335;
    wire N__5332;
    wire N__5329;
    wire N__5326;
    wire N__5323;
    wire N__5320;
    wire N__5317;
    wire N__5314;
    wire N__5311;
    wire N__5308;
    wire N__5305;
    wire N__5302;
    wire N__5299;
    wire N__5296;
    wire N__5293;
    wire N__5290;
    wire N__5287;
    wire N__5284;
    wire N__5281;
    wire N__5278;
    wire N__5275;
    wire N__5272;
    wire N__5269;
    wire N__5266;
    wire N__5263;
    wire N__5260;
    wire N__5257;
    wire N__5254;
    wire N__5251;
    wire N__5250;
    wire N__5247;
    wire N__5244;
    wire N__5243;
    wire N__5242;
    wire N__5239;
    wire N__5236;
    wire N__5233;
    wire N__5230;
    wire N__5229;
    wire N__5220;
    wire N__5217;
    wire N__5216;
    wire N__5215;
    wire N__5214;
    wire N__5209;
    wire N__5206;
    wire N__5203;
    wire N__5200;
    wire N__5197;
    wire N__5194;
    wire N__5189;
    wire N__5184;
    wire N__5181;
    wire N__5178;
    wire N__5175;
    wire N__5172;
    wire N__5169;
    wire N__5166;
    wire N__5161;
    wire N__5158;
    wire N__5155;
    wire N__5152;
    wire N__5149;
    wire N__5146;
    wire N__5143;
    wire N__5140;
    wire N__5137;
    wire N__5134;
    wire N__5131;
    wire N__5128;
    wire N__5125;
    wire N__5122;
    wire N__5119;
    wire N__5116;
    wire N__5113;
    wire N__5110;
    wire N__5107;
    wire N__5104;
    wire N__5101;
    wire N__5098;
    wire N__5095;
    wire N__5092;
    wire N__5089;
    wire N__5086;
    wire N__5083;
    wire N__5080;
    wire N__5077;
    wire N__5074;
    wire N__5071;
    wire N__5068;
    wire N__5065;
    wire N__5062;
    wire N__5059;
    wire N__5056;
    wire N__5053;
    wire N__5050;
    wire N__5047;
    wire N__5044;
    wire N__5041;
    wire N__5038;
    wire N__5035;
    wire N__5032;
    wire N__5029;
    wire N__5026;
    wire N__5023;
    wire N__5020;
    wire N__5017;
    wire wRamRdData_6;
    wire wRamRdData_2;
    wire wRamRdData_3;
    wire wRamRdData_5;
    wire BTN_N_c;
    wire wRamRdData_7;
    wire wRamRdData_0;
    wire VCCG0;
    wire wRamRdData_4;
    wire wRamRdData_1;
    wire GNDG0;
    wire \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO ;
    wire \DUT.fifo_rx_inst.N_86_cascade_ ;
    wire \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1 ;
    wire \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1_cascade_ ;
    wire oTx_n_c_i;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_4 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_4 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_5 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_5 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_5 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_6 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_6 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_6 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_4 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_3 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_3 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_3 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_awe2 ;
    wire \DUT.fifo_rx_inst.rFifoData_awe2_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoDataro_3 ;
    wire \DUT.fifo_rx_inst.rFifoDataro_2 ;
    wire \DUT.fifo_rx_inst.N_42 ;
    wire \DUT.fifo_rx_inst.rWritePtrZ0Z_0 ;
    wire \DUT.fifo_rx_inst.N_42_cascade_ ;
    wire \DUT.fifo_rx_inst.rWritePtrZ0Z_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_awe1_cascade_ ;
    wire \DUT.fifo_tx_inst.un1_i11_i ;
    wire \DUT.fifo_tx_inst.un1_i11_i_cascade_ ;
    wire wRxBufferEmpty_i_0_cascade_;
    wire \DUT.fifo_rx_inst.un1_rFifoCount16_0_i_0 ;
    wire bfn_13_18_0_;
    wire \DUT.fifo_rx_inst.rFifoCount_RNIK3G92Z0Z_1 ;
    wire \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0 ;
    wire \DUT.fifo_rx_inst.un1_rFifoCount_1_axb_2 ;
    wire \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1 ;
    wire \DUT.fifo_rx_inst.rFifoCountZ0Z_2 ;
    wire \DUT.fifo_rx_inst.rFifoCountZ0Z_1 ;
    wire \DUT.fifo_tx_inst.N_35_cascade_ ;
    wire G_143_cascade_;
    wire \fifo_inst.ftdi_input_inst.SUMZ0Z_2_cascade_ ;
    wire \DUT.fifo_rx_inst.N_86 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_7 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_7 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_2 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_2 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_2 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1_cascade_ ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_7 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram0_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram3_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram2_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ;
    wire wRxBufferEmpty_i_0_0;
    wire \DUT.fifo_rx_inst.rFifoDataro_1 ;
    wire \DUT.fifo_rx_inst.rTxByte_42_0 ;
    wire \DUT.fifo_rx_inst.rTxByte_42_1_cascade_ ;
    wire wRxBufferEmpty_i_0;
    wire rFifoDatarff_0_RNIHJV05;
    wire \DUT.fifo_rx_inst.rReadPtrZ0Z_1 ;
    wire \DUT.fifo_rx_inst.rReadPtr_RNI4NC92Z0Z_0 ;
    wire \DUT.fifo_rx_inst.N_73 ;
    wire \DUT.fifo_rx_inst.rReadPtr_RNI4NC92Z0Z_0_cascade_ ;
    wire \DUT.fifo_rx_inst.rReadPtrZ0Z_0 ;
    wire \DUT.uart_inst0.recv_state_srsts_1_0_6_cascade_ ;
    wire \DUT.fifo_rx_inst.un1_rFifoCount16_0_0 ;
    wire \DUT.fifo_rx_inst.rFifoCountZ0Z_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_awe0 ;
    wire \DUT.fifo_rx_inst.rFifoDataro_0 ;
    wire oTx_n_c;
    wire P1A2_c;
    wire \DUT.fifo_tx_inst.rFifoCountZ0Z_0 ;
    wire \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0 ;
    wire bfn_14_19_0_;
    wire \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0 ;
    wire \DUT.fifo_tx_inst.N_35 ;
    wire \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1 ;
    wire \DUT.fifo_tx_inst.rFifoDataro_3 ;
    wire \DUT.fifo_tx_inst.rFifoDataro_2 ;
    wire \DUT.fifo_tx_inst.rFifoDataro_1 ;
    wire \DUT.fifo_tx_inst.rFifoDataro_0 ;
    wire \DUT.fifo_tx_inst.rFifoDataror_1_0_cascade_ ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ;
    wire \DUT.fifo_tx_inst.un1_i11_2_i_cascade_ ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_3 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_3 ;
    wire \DUT.fifo_tx_inst.CO0 ;
    wire \DUT.fifo_tx_inst.CO0_cascade_ ;
    wire \DUT.fifo_tx_inst.un1_i11_2_i ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_5 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_5 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_5 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_7 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_7 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_ ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_7 ;
    wire \DUT.fifo_tx_inst.N_33 ;
    wire \DUT.fifo_tx_inst.N_41 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_4 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_4 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_ ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_2 ;
    wire \DUT.rFifoDatarx_2_cascade_ ;
    wire \DUT.fifo_tx_inst.N_40 ;
    wire G_145_cascade_;
    wire G_145;
    wire G_142_cascade_;
    wire G_144;
    wire \fifo_inst.ftdi_input_inst.SUMZ0Z_3 ;
    wire G_147;
    wire G_142;
    wire G_141;
    wire G_141_cascade_;
    wire G_140;
    wire fifo_inst_ftdi_input_inst_oTxFull_0;
    wire G_140_cascade_;
    wire G_143;
    wire G_146;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_0 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_1 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_2 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_3 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_4 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_5 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_6 ;
    wire \DUT.fifo_rx_inst.rFifoData_ram1_7 ;
    wire \DUT.fifo_rx_inst.rFifoData_awe1 ;
    wire \DUT.wRxByte_0 ;
    wire \DUT.wRxByte_1 ;
    wire \DUT.wRxByte_2 ;
    wire \DUT.wRxByte_3 ;
    wire \DUT.wRxByte_4 ;
    wire \DUT.wRxByte_5 ;
    wire \DUT.wRxByte_6 ;
    wire \DUT.wRxByte_7 ;
    wire \DUT.uart_inst0.rx_bits_remaining_2_sqmuxa ;
    wire \DUT.uart_inst0.rx_countdown_3_2_cascade_ ;
    wire \DUT.wRcvd ;
    wire \DUT.uart_inst0.rx_countdown_8_i_o2_2_1_2_cascade_ ;
    wire \DUT.uart_inst0.rx_countdown_8_i_o2_2_2_cascade_ ;
    wire \DUT.uart_inst0.recv_state_RNO_0Z0Z_1_cascade_ ;
    wire \DUT.uart_inst0.un1_m2_e_0_cascade_ ;
    wire \DUT.uart_inst0.N_69 ;
    wire \DUT.uart_inst0.recv_state_RNITN8GJZ0Z_2_cascade_ ;
    wire \DUT.uart_inst0.recv_state_RNITN8GJZ0Z_2 ;
    wire \DUT.uart_inst0.rx_bits_remainingZ0Z_2 ;
    wire \DUT.uart_inst0.rx_bits_remainingZ0Z_1 ;
    wire \DUT.uart_inst0.rx_bits_remainingZ0Z_3 ;
    wire \DUT.uart_inst0.rx_bits_remainingZ0Z_0 ;
    wire \DUT.uart_inst0.N_98_4_cascade_ ;
    wire \DUT.uart_inst0.rx_m2_e_0 ;
    wire \DUT.uart_inst0.r_N_5_mux_cascade_ ;
    wire \DUT.uart_inst0.recv_stateZ0Z_2 ;
    wire \DUT.uart_inst0.N_98_4 ;
    wire \DUT.uart_inst0.r_N_3_mux_cascade_ ;
    wire \DUT.uart_inst0.recv_N_5_mux ;
    wire \DUT.uart_inst0.g3_cascade_ ;
    wire \DUT.uart_inst0.g3_1 ;
    wire \DUT.uart_inst0.tx_countdown_0_c3 ;
    wire \DUT.uart_inst0.un1_m7_3 ;
    wire \DUT.uart_inst0.un1_tx_state_0_a4_1_cascade_ ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_s1_sn_0_cascade_ ;
    wire \DUT.uart_inst0.tx_countdown_7_1_0_3 ;
    wire \DUT.uart_inst0.tx_countdown_RNO_0Z0Z_1_cascade_ ;
    wire \DUT.uart_inst0.g0_i_o4_0_4_cascade_ ;
    wire \DUT.fifo_tx_inst.rWritePtrZ0Z_1 ;
    wire \DUT.fifo_tx_inst.rWritePtrZ0Z_0 ;
    wire \DUT.fifo_tx_inst.rFifoCountZ0Z_2 ;
    wire \DUT.rFifoDatarxZ0Z_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_4 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4 ;
    wire \DUT.rFifoDatarx_4_cascade_ ;
    wire \DUT.uart_inst0.tx_data_RNO_0Z0Z_4 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram1_6 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram0_6 ;
    wire \DUT.fifo_tx_inst.rReadPtrZ0Z_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_ ;
    wire \DUT.uart_inst0.tx_data_RNO_0Z0Z_2 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_0 ;
    wire rTxByteZ0Z_2;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_2 ;
    wire rTxByteZ0Z_4;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_4 ;
    wire rTxByteZ0Z_5;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_5 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_6 ;
    wire rTxByteZ0Z_7;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_7 ;
    wire \DUT.fifo_tx_inst.rFifoData_awe3 ;
    wire \DUT.rFifoDatarx_7 ;
    wire G_152_cascade_;
    wire G_151;
    wire G_150;
    wire \fifo_inst.ftdi_input_inst.un1_rWrStateZ0Z_1 ;
    wire G_149;
    wire \fifo_inst.ftdi_input_inst.un2_oPacketAvail_iZ0 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_10_cascade_ ;
    wire \DUT.uart_inst0.rx_clk_divider_RNIKU472Z0Z_10 ;
    wire \DUT.uart_inst0.recv_state_RNO_0Z0Z_0 ;
    wire \DUT.uart_inst0.recv_state_RNO_1Z0Z_0_cascade_ ;
    wire \DUT.uart_inst0.recv_stateZ0Z_0 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_10 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_0_cascade_ ;
    wire \DUT.uart_inst0.rx_countdown_3_2 ;
    wire \DUT.uart_inst0.rx_countdown_8_i_o2_1_2_cascade_ ;
    wire \DUT.uart_inst0.recv_state_RNO_0Z0Z_4_cascade_ ;
    wire \DUT.uart_inst0.recv_stateZ0Z_4 ;
    wire \DUT.uart_inst0.recv_stateZ0Z_5 ;
    wire \DUT.uart_inst0.recv_stateZ0Z_3 ;
    wire P1A1_c;
    wire \DUT.uart_inst0.recv_stateZ0Z_1 ;
    wire \DUT.uart_inst0.recv_state_srsts_1_5 ;
    wire bfn_16_16_0_;
    wire \DUT.uart_inst0.rx_countdown_3_s1_1 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_0_s1 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_1_s1_THRU_CO ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_1_s1 ;
    wire \DUT.uart_inst0.rx_countdown_3_s1_3 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_2_s1 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_3_s1 ;
    wire \DUT.uart_inst0.rx_countdown_3_cry_4_s1 ;
    wire \DUT.uart_inst0.N_105 ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_1 ;
    wire \DUT.uart_inst0.N_102 ;
    wire \DUT.uart_inst0.rx_countdownZ1Z_3 ;
    wire \DUT.uart_inst0.rx_countdown_8_i_o2_1_1_2 ;
    wire \DUT.uart_inst0.rx_countdown_3_s1_4 ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_4 ;
    wire \DUT.uart_inst0.rx_countdown_RNO_0Z0Z_2 ;
    wire \DUT.uart_inst0.rx_countdown_8_i_o2_1_2 ;
    wire \DUT.uart_inst0.rx_countdown_RNO_1Z0Z_2 ;
    wire \DUT.uart_inst0.rx_countdown_8_i_o2_2_2 ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_2 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_6_cascade_ ;
    wire \DUT.uart_inst0.un1_tx_bits_remaining_axbxc2_N_4L5_1_1 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_0_cascade_ ;
    wire \DUT.uart_inst0.un1_tx_bits_remaining_axbxc2_N_4L5_1 ;
    wire rRxReadZ0;
    wire \DUT.fifo_tx_inst.rFifoCountZ0Z_1 ;
    wire \DUT.fifo_tx_inst.rFifoCount_RNIBPFMZ0Z_1 ;
    wire \DUT.uart_inst0.g0_0_0_a3_3_cascade_ ;
    wire \DUT.uart_inst0.g0_0_0_a3_5_cascade_ ;
    wire \DUT.uart_inst0.N_159_0_0 ;
    wire \DUT.N_37 ;
    wire \DUT.uart_inst0.tx_countdown_0_1_5_cascade_ ;
    wire \DUT.uart_inst0.g0_i_o4_0_5 ;
    wire \DUT.uart_inst0.N_14_cascade_ ;
    wire P1A7_c;
    wire \DUT.uart_inst0.N_6 ;
    wire \DUT.uart_inst0.un1_tx_bits_remaining_axbxc2_N_4L5_1_0 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_1 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_2 ;
    wire \DUT.rFifoDatarx_1_cascade_ ;
    wire \DUT.uart_inst0.tx_data_RNO_0Z0Z_1_cascade_ ;
    wire \DUT.uart_inst0.tx_dataZ0Z_1 ;
    wire \DUT.uart_inst0.tx_data_RNO_0Z0Z_0 ;
    wire \DUT.rFifoDatarx_5 ;
    wire \DUT.uart_inst0.tx_data_RNO_0Z0Z_5_cascade_ ;
    wire \DUT.uart_inst0.tx_dataZ0Z_5 ;
    wire rTxByteZ0Z_1;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_1 ;
    wire rTxByteZ0Z_0;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_0 ;
    wire rTxByteZ0Z_6;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_6 ;
    wire \DUT.uart_inst0.tx_data_8_321_a2_0 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_11 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_12 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_9_cascade_ ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_a_13 ;
    wire \DUT.uart_inst0.rx_countdown_3_s1_5 ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_5 ;
    wire \DUT.uart_inst0.un2_rx_clk_divider_0 ;
    wire \DUT.uart_inst0.N_70 ;
    wire \DUT.uart_inst0.rx_countdownZ0Z_3 ;
    wire G_148;
    wire \fifo_inst.ftdi_output_inst.N_95_cascade_ ;
    wire \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_3 ;
    wire \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2 ;
    wire \fifo_inst.ftdi_output_inst.N_95 ;
    wire \fifo_inst.ftdi_output_inst.m14_1_cascade_ ;
    wire \fifo_inst.ftdi_output_inst.N_86_0 ;
    wire \DUT.uart_inst0.tx_bits_remaining_RNO_1Z0Z_2 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_9 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_8 ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_7 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_3 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_5 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_2 ;
    wire \DUT.uart_inst0.tx_data_i_m_4_0_cascade_ ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_4 ;
    wire \DUT.uart_inst0.tx_countdown_0_c4_i ;
    wire \DUT.uart_inst0.tx_state_ns_0_o3_1_0_1 ;
    wire \DUT.rFifoDatarx_6 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_7 ;
    wire \DUT.uart_inst0.tx_data_RNO_0Z0Z_6_cascade_ ;
    wire \DUT.uart_inst0.tx_dataZ0Z_6 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_4 ;
    wire \DUT.rFifoDataror_0 ;
    wire \DUT.uart_inst0.tx_data_RNO_0Z0Z_3_cascade_ ;
    wire \DUT.uart_inst0.N_152_0 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_3 ;
    wire \DUT.uart_inst0.N_159 ;
    wire \DUT.uart_inst0.tx_dataZ0Z_0 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_1 ;
    wire \DUT.uart_inst0.g0_i_a4_0_4 ;
    wire \DUT.uart_inst0.tx_countdownZ0Z_0 ;
    wire \DUT.uart_inst0.g0_i_a4_0_5_cascade_ ;
    wire \DUT.uart_inst0.N_15 ;
    wire \DUT.uart_inst0.N_7 ;
    wire \DUT.fifo_tx_inst.rReadPtrZ0Z_1 ;
    wire \DUT.fifo_tx_inst.rFifoData_ram3_3 ;
    wire \DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3 ;
    wire \DUT.rFifoDatarx_3 ;
    wire \DUT.uart_inst0.tx_bits_remainingZ0Z_3 ;
    wire \DUT.uart_inst0.tx_state_ns_i_i_a2_0_0_0_cascade_ ;
    wire \DUT.uart_inst0.g0_i_a4_1_0 ;
    wire \DUT.uart_inst0.d_N_5_mux ;
    wire rTxByteZ0Z_3;
    wire \DUT.fifo_tx_inst.rFifoData_ram2_3 ;
    wire \DUT.fifo_tx_inst.N_39 ;
    wire \fifo_inst.ftdi_output_inst.rTxE_nZ0Z_1 ;
    wire iTxE_n_c;
    wire \fifo_inst.ftdi_output_inst.rTxE_nZ0Z_0 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_1 ;
    wire bfn_18_13_0_;
    wire \DUT.uart_inst0.rx_clk_dividerZ1Z_1 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_0 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_2 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_1 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_3 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_2_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_2 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_4 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_3 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_5 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_4_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_4 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_6 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_5_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_5 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_7 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_6 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_7 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_8 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO ;
    wire bfn_18_14_0_;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_9 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_8 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_10 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_9 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_11 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_10 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_12 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_11 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_13 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_12 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_14 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_13 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_15 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_14 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_15 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_16 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO ;
    wire bfn_18_15_0_;
    wire \DUT.uart_inst0.N_72 ;
    wire \DUT.uart_inst0.rx_clk_divider_1_cry_16 ;
    wire \DUT.uart_inst0.rx_clk_dividerZ0Z_17 ;
    wire \fifo_inst.wRamRdAddr_2 ;
    wire \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4 ;
    wire \fifo_inst.ftdi_output_inst.rWrDelayZ0 ;
    wire \fifo_inst.ftdi_output_inst.N_3_0 ;
    wire \fifo_inst.wRamRdAddr_0 ;
    wire \fifo_inst.ftdi_output_inst.N_3_0_cascade_ ;
    wire \fifo_inst.wRamRdAddr_1 ;
    wire \DUT.uart_inst0.tx_state_ns_i_i_a2_0_0_0 ;
    wire \DUT.uart_inst0.tx_state_0_sqmuxa_i_0 ;
    wire wPllLocked_iso_i;
    wire \DUT.uart_inst0.N_345_0_0 ;
    wire \DUT.uart_inst0.tx_bits_remaining_0_sqmuxa ;
    wire \DUT.rTransmitZ0 ;
    wire \DUT.uart_inst0.tx_clk_divider_0_sqmuxa ;
    wire wPllLocked;
    wire \DUT.uart_inst0.tx_clk_divider_0_sqmuxa_cascade_ ;
    wire \DUT.uart_inst0.un1_tx_clk_divider_0 ;
    wire \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0 ;
    wire \fifo_inst.ftdi_output_inst.rRxF_nZ0Z_1 ;
    wire \fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_0 ;
    wire bfn_18_19_0_;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_1 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_0 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_2 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_1 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_3 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_2 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_4 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_3 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_5 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_4 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_6 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_5 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_7 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_6 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_7 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_8 ;
    wire bfn_18_20_0_;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_9 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_8 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_10 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_9 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_11 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_10 ;
    wire CONSTANT_ONE_NET;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_12 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_11 ;
    wire \DUT.uart_inst0.tx_clk_divider_cry_12 ;
    wire \DUT.uart_inst0.tx_clk_dividerZ0Z_13 ;
    wire \DUT.uart_inst0.tx_clk_divider_1_sqmuxa_1_i ;
    wire \DUT.uart_inst0.tx_state_ns_i_i_0_0 ;
    wire \DUT.uart_inst0.N_345_0 ;
    wire \DUT.uart_inst0.tx_state_ns_i_i_a2_0_1_0 ;
    wire \DUT.tx_state_0 ;
    wire wPllLocked_iso_i_g;
    wire \DUT.uart_inst0.tx_bits_remainingZ0Z_2 ;
    wire \DUT.uart_inst0.tx_bits_remainingZ0Z_0 ;
    wire \DUT.uart_inst0.tx_bits_remaining_RNO_0Z0Z_3 ;
    wire \DUT.tx_state_1 ;
    wire \DUT.uart_inst0.tx_bits_remainingZ0Z_1 ;
    wire \DUT.uart_inst0.tx_bits_remaining_RNO_0Z0Z_2 ;
    wire iRxF_n_c;
    wire \fifo_inst.ftdi_output_inst.rRxF_nZ0Z_0 ;
    wire clk_48mhz;
    wire wPllLocked_g;
    wire _gnd_net_;

    defparam \fifo_inst.ftdi_input_inst.ram512x8_inst_physical .WRITE_MODE=1;
    defparam \fifo_inst.ftdi_input_inst.ram512x8_inst_physical .READ_MODE=1;
    SB_RAM40_4K \fifo_inst.ftdi_input_inst.ram512x8_inst_physical  (
            .RDATA({dangling_wire_0,wRamRdData_7,dangling_wire_1,wRamRdData_6,dangling_wire_2,wRamRdData_5,dangling_wire_3,wRamRdData_4,dangling_wire_4,wRamRdData_3,dangling_wire_5,wRamRdData_2,dangling_wire_6,wRamRdData_1,dangling_wire_7,wRamRdData_0}),
            .RADDR({dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,N__11068,N__10945,N__10975}),
            .WADDR({dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,N__7876,N__7855,N__7819}),
            .MASK({dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39}),
            .WDATA({dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55}),
            .RCLKE(),
            .RCLK(GNDG0),
            .RE(N__13008),
            .WCLKE(),
            .WCLK(N__12139),
            .WE(N__6523));
    defparam \top_pll_inst.top_pll_inst_pll .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \top_pll_inst.top_pll_inst_pll .TEST_MODE=1'b0;
    defparam \top_pll_inst.top_pll_inst_pll .SHIFTREG_DIV_MODE=2'b00;
    defparam \top_pll_inst.top_pll_inst_pll .PLLOUT_SELECT="GENCLK";
    defparam \top_pll_inst.top_pll_inst_pll .FILTER_RANGE=3'b001;
    defparam \top_pll_inst.top_pll_inst_pll .FEEDBACK_PATH="SIMPLE";
    defparam \top_pll_inst.top_pll_inst_pll .FDA_RELATIVE=4'b0000;
    defparam \top_pll_inst.top_pll_inst_pll .FDA_FEEDBACK=4'b0000;
    defparam \top_pll_inst.top_pll_inst_pll .ENABLE_ICEGATE=1'b0;
    defparam \top_pll_inst.top_pll_inst_pll .DIVR=4'b0000;
    defparam \top_pll_inst.top_pll_inst_pll .DIVQ=3'b100;
    defparam \top_pll_inst.top_pll_inst_pll .DIVF=7'b0111111;
    defparam \top_pll_inst.top_pll_inst_pll .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    PLL40 \top_pll_inst.top_pll_inst_pll  (
            .PLLOUTGLOBAL(clk_48mhz),
            .SDI(GNDG0),
            .BYPASS(GNDG0),
            .RESETB(N__5137),
            .PLLOUTCORE(),
            .LOCK(\PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO ),
            .SDO(),
            .SCLK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .EXTFEEDBACK(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLIN(N__13213));
    IO_PAD \top_pll_inst.top_pll_inst_iopad  (
            .OE(VCCG0),
            .DIN(),
            .DOUT(N__13213),
            .PACKAGEPIN(iClk));
    IO_PAD P1A8_obuft_iopad (
            .OE(N__13199),
            .DIN(N__13198),
            .DOUT(N__13197),
            .PACKAGEPIN(P1A8));
    defparam P1A8_obuft_preio.NEG_TRIGGER=1'b0;
    defparam P1A8_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO P1A8_obuft_preio (
            .PADOEN(N__13199),
            .PADOUT(N__13198),
            .PADIN(N__13197),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_1_iopad (
            .OE(N__13190),
            .DIN(N__13189),
            .DOUT(N__13188),
            .PACKAGEPIN(ioFifoData[1]));
    defparam ioFifoData_obuft_1_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_1_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_1_preio (
            .PADOEN(N__13190),
            .PADOUT(N__13189),
            .PADIN(N__13188),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5229),
            .DIN0(),
            .DOUT0(N__5161),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A9_obuft_iopad (
            .OE(N__13181),
            .DIN(N__13180),
            .DOUT(N__13179),
            .PACKAGEPIN(P1A9));
    defparam P1A9_obuft_preio.NEG_TRIGGER=1'b0;
    defparam P1A9_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO P1A9_obuft_preio (
            .PADOEN(N__13181),
            .PADOUT(N__13180),
            .PADIN(N__13179),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_4_iopad (
            .OE(N__13172),
            .DIN(N__13171),
            .DOUT(N__13170),
            .PACKAGEPIN(ioFifoData[4]));
    defparam ioFifoData_obuft_4_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_4_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_4_preio (
            .PADOEN(N__13172),
            .PADOUT(N__13171),
            .PADIN(N__13170),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5243),
            .DIN0(),
            .DOUT0(N__5086),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_0_iopad (
            .OE(N__13163),
            .DIN(N__13162),
            .DOUT(N__13161),
            .PACKAGEPIN(ioFifoData[0]));
    defparam ioFifoData_obuft_0_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_0_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_0_preio (
            .PADOEN(N__13163),
            .PADOUT(N__13162),
            .PADIN(N__13161),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5216),
            .DIN0(),
            .DOUT0(N__5107),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD oRx_n_obuf_iopad (
            .OE(N__13154),
            .DIN(N__13153),
            .DOUT(N__13152),
            .PACKAGEPIN(oRx_n));
    defparam oRx_n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam oRx_n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO oRx_n_obuf_preio (
            .PADOEN(N__13154),
            .PADOUT(N__13153),
            .PADIN(N__13152),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__13018),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A2_obuf_iopad (
            .OE(N__13145),
            .DIN(N__13144),
            .DOUT(N__13143),
            .PACKAGEPIN(P1A2));
    defparam P1A2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO P1A2_obuf_preio (
            .PADOEN(N__13145),
            .PADOUT(N__13144),
            .PADIN(N__13143),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6181),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_7_iopad (
            .OE(N__13136),
            .DIN(N__13135),
            .DOUT(N__13134),
            .PACKAGEPIN(ioFifoData[7]));
    defparam ioFifoData_obuft_7_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_7_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_7_preio (
            .PADOEN(N__13136),
            .PADOUT(N__13135),
            .PADIN(N__13134),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5215),
            .DIN0(),
            .DOUT0(N__5122),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD iRxF_n_ibuf_iopad (
            .OE(N__13127),
            .DIN(N__13126),
            .DOUT(N__13125),
            .PACKAGEPIN(iRxF_n));
    defparam iRxF_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam iRxF_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO iRxF_n_ibuf_preio (
            .PADOEN(N__13127),
            .PADOUT(N__13126),
            .PADIN(N__13125),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(iRxF_n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A3_obuf_iopad (
            .OE(N__13118),
            .DIN(N__13117),
            .DOUT(N__13116),
            .PACKAGEPIN(P1A3));
    defparam P1A3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO P1A3_obuf_preio (
            .PADOEN(N__13118),
            .PADOUT(N__13117),
            .PADIN(N__13116),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A7_obuf_iopad (
            .OE(N__13109),
            .DIN(N__13108),
            .DOUT(N__13107),
            .PACKAGEPIN(P1A7));
    defparam P1A7_obuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A7_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO P1A7_obuf_preio (
            .PADOEN(N__13109),
            .PADOUT(N__13108),
            .PADIN(N__13107),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8809),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BTN_N_ibuf_iopad (
            .OE(N__13100),
            .DIN(N__13099),
            .DOUT(N__13098),
            .PACKAGEPIN(BTN_N));
    defparam BTN_N_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam BTN_N_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO BTN_N_ibuf_preio (
            .PADOEN(N__13100),
            .PADOUT(N__13099),
            .PADIN(N__13098),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(BTN_N_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_3_iopad (
            .OE(N__13091),
            .DIN(N__13090),
            .DOUT(N__13089),
            .PACKAGEPIN(ioFifoData[3]));
    defparam ioFifoData_obuft_3_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_3_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_3_preio (
            .PADOEN(N__13091),
            .PADOUT(N__13090),
            .PADIN(N__13089),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5250),
            .DIN0(),
            .DOUT0(N__5044),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_6_iopad (
            .OE(N__13082),
            .DIN(N__13081),
            .DOUT(N__13080),
            .PACKAGEPIN(ioFifoData[6]));
    defparam ioFifoData_obuft_6_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_6_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_6_preio (
            .PADOEN(N__13082),
            .PADOUT(N__13081),
            .PADIN(N__13080),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5214),
            .DIN0(),
            .DOUT0(N__5074),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_5_iopad (
            .OE(N__13073),
            .DIN(N__13072),
            .DOUT(N__13071),
            .PACKAGEPIN(ioFifoData[5]));
    defparam ioFifoData_obuft_5_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_5_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_5_preio (
            .PADOEN(N__13073),
            .PADOUT(N__13072),
            .PADIN(N__13071),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5242),
            .DIN0(),
            .DOUT0(N__5026),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD oTx_n_obuf_iopad (
            .OE(N__13064),
            .DIN(N__13063),
            .DOUT(N__13062),
            .PACKAGEPIN(oTx_n));
    defparam oTx_n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam oTx_n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO oTx_n_obuf_preio (
            .PADOEN(N__13064),
            .PADOUT(N__13063),
            .PADIN(N__13062),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6214),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD iTxE_n_ibuf_iopad (
            .OE(N__13055),
            .DIN(N__13054),
            .DOUT(N__13053),
            .PACKAGEPIN(iTxE_n));
    defparam iTxE_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam iTxE_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO iTxE_n_ibuf_preio (
            .PADOEN(N__13055),
            .PADOUT(N__13054),
            .PADIN(N__13053),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(iTxE_n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_obuft_2_iopad (
            .OE(N__13046),
            .DIN(N__13045),
            .DOUT(N__13044),
            .PACKAGEPIN(ioFifoData[2]));
    defparam ioFifoData_obuft_2_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_obuft_2_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_obuft_2_preio (
            .PADOEN(N__13046),
            .PADOUT(N__13045),
            .PADIN(N__13044),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__5251),
            .DIN0(),
            .DOUT0(N__5062),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A1_ibuf_iopad (
            .OE(N__13037),
            .DIN(N__13036),
            .DOUT(N__13035),
            .PACKAGEPIN(P1A1));
    defparam P1A1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO P1A1_ibuf_preio (
            .PADOEN(N__13037),
            .PADOUT(N__13036),
            .PADIN(N__13035),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(P1A1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IoInMux I__3084 (
            .O(N__13018),
            .I(N__13015));
    LocalMux I__3083 (
            .O(N__13015),
            .I(N__13012));
    IoSpan4Mux I__3082 (
            .O(N__13012),
            .I(N__13009));
    Span4Mux_s3_v I__3081 (
            .O(N__13009),
            .I(N__13005));
    SRMux I__3080 (
            .O(N__13008),
            .I(N__13002));
    Span4Mux_v I__3079 (
            .O(N__13005),
            .I(N__12972));
    LocalMux I__3078 (
            .O(N__13002),
            .I(N__12972));
    InMux I__3077 (
            .O(N__13001),
            .I(N__12967));
    InMux I__3076 (
            .O(N__13000),
            .I(N__12967));
    InMux I__3075 (
            .O(N__12999),
            .I(N__12960));
    InMux I__3074 (
            .O(N__12998),
            .I(N__12960));
    InMux I__3073 (
            .O(N__12997),
            .I(N__12960));
    CascadeMux I__3072 (
            .O(N__12996),
            .I(N__12957));
    CascadeMux I__3071 (
            .O(N__12995),
            .I(N__12954));
    CascadeMux I__3070 (
            .O(N__12994),
            .I(N__12951));
    CascadeMux I__3069 (
            .O(N__12993),
            .I(N__12948));
    CascadeMux I__3068 (
            .O(N__12992),
            .I(N__12944));
    CascadeMux I__3067 (
            .O(N__12991),
            .I(N__12941));
    CascadeMux I__3066 (
            .O(N__12990),
            .I(N__12938));
    CascadeMux I__3065 (
            .O(N__12989),
            .I(N__12935));
    CascadeMux I__3064 (
            .O(N__12988),
            .I(N__12932));
    CascadeMux I__3063 (
            .O(N__12987),
            .I(N__12929));
    CascadeMux I__3062 (
            .O(N__12986),
            .I(N__12926));
    CascadeMux I__3061 (
            .O(N__12985),
            .I(N__12923));
    CascadeMux I__3060 (
            .O(N__12984),
            .I(N__12920));
    CascadeMux I__3059 (
            .O(N__12983),
            .I(N__12917));
    CascadeMux I__3058 (
            .O(N__12982),
            .I(N__12914));
    CascadeMux I__3057 (
            .O(N__12981),
            .I(N__12911));
    CascadeMux I__3056 (
            .O(N__12980),
            .I(N__12908));
    CascadeMux I__3055 (
            .O(N__12979),
            .I(N__12905));
    CascadeMux I__3054 (
            .O(N__12978),
            .I(N__12902));
    CascadeMux I__3053 (
            .O(N__12977),
            .I(N__12899));
    Span4Mux_v I__3052 (
            .O(N__12972),
            .I(N__12889));
    LocalMux I__3051 (
            .O(N__12967),
            .I(N__12884));
    LocalMux I__3050 (
            .O(N__12960),
            .I(N__12884));
    InMux I__3049 (
            .O(N__12957),
            .I(N__12879));
    InMux I__3048 (
            .O(N__12954),
            .I(N__12879));
    InMux I__3047 (
            .O(N__12951),
            .I(N__12868));
    InMux I__3046 (
            .O(N__12948),
            .I(N__12868));
    InMux I__3045 (
            .O(N__12947),
            .I(N__12868));
    InMux I__3044 (
            .O(N__12944),
            .I(N__12868));
    InMux I__3043 (
            .O(N__12941),
            .I(N__12868));
    InMux I__3042 (
            .O(N__12938),
            .I(N__12859));
    InMux I__3041 (
            .O(N__12935),
            .I(N__12859));
    InMux I__3040 (
            .O(N__12932),
            .I(N__12859));
    InMux I__3039 (
            .O(N__12929),
            .I(N__12859));
    InMux I__3038 (
            .O(N__12926),
            .I(N__12850));
    InMux I__3037 (
            .O(N__12923),
            .I(N__12850));
    InMux I__3036 (
            .O(N__12920),
            .I(N__12850));
    InMux I__3035 (
            .O(N__12917),
            .I(N__12850));
    InMux I__3034 (
            .O(N__12914),
            .I(N__12847));
    InMux I__3033 (
            .O(N__12911),
            .I(N__12842));
    InMux I__3032 (
            .O(N__12908),
            .I(N__12842));
    InMux I__3031 (
            .O(N__12905),
            .I(N__12835));
    InMux I__3030 (
            .O(N__12902),
            .I(N__12835));
    InMux I__3029 (
            .O(N__12899),
            .I(N__12835));
    CascadeMux I__3028 (
            .O(N__12898),
            .I(N__12832));
    CascadeMux I__3027 (
            .O(N__12897),
            .I(N__12829));
    CascadeMux I__3026 (
            .O(N__12896),
            .I(N__12826));
    CascadeMux I__3025 (
            .O(N__12895),
            .I(N__12823));
    CascadeMux I__3024 (
            .O(N__12894),
            .I(N__12820));
    CascadeMux I__3023 (
            .O(N__12893),
            .I(N__12817));
    CascadeMux I__3022 (
            .O(N__12892),
            .I(N__12814));
    Span4Mux_v I__3021 (
            .O(N__12889),
            .I(N__12811));
    Span4Mux_v I__3020 (
            .O(N__12884),
            .I(N__12808));
    LocalMux I__3019 (
            .O(N__12879),
            .I(N__12799));
    LocalMux I__3018 (
            .O(N__12868),
            .I(N__12799));
    LocalMux I__3017 (
            .O(N__12859),
            .I(N__12799));
    LocalMux I__3016 (
            .O(N__12850),
            .I(N__12799));
    LocalMux I__3015 (
            .O(N__12847),
            .I(N__12792));
    LocalMux I__3014 (
            .O(N__12842),
            .I(N__12792));
    LocalMux I__3013 (
            .O(N__12835),
            .I(N__12792));
    InMux I__3012 (
            .O(N__12832),
            .I(N__12785));
    InMux I__3011 (
            .O(N__12829),
            .I(N__12785));
    InMux I__3010 (
            .O(N__12826),
            .I(N__12785));
    InMux I__3009 (
            .O(N__12823),
            .I(N__12776));
    InMux I__3008 (
            .O(N__12820),
            .I(N__12776));
    InMux I__3007 (
            .O(N__12817),
            .I(N__12776));
    InMux I__3006 (
            .O(N__12814),
            .I(N__12776));
    Odrv4 I__3005 (
            .O(N__12811),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3004 (
            .O(N__12808),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__3003 (
            .O(N__12799),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__3002 (
            .O(N__12792),
            .I(CONSTANT_ONE_NET));
    LocalMux I__3001 (
            .O(N__12785),
            .I(CONSTANT_ONE_NET));
    LocalMux I__3000 (
            .O(N__12776),
            .I(CONSTANT_ONE_NET));
    InMux I__2999 (
            .O(N__12763),
            .I(N__12759));
    InMux I__2998 (
            .O(N__12762),
            .I(N__12756));
    LocalMux I__2997 (
            .O(N__12759),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_12 ));
    LocalMux I__2996 (
            .O(N__12756),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_12 ));
    InMux I__2995 (
            .O(N__12751),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_11 ));
    InMux I__2994 (
            .O(N__12748),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_12 ));
    CascadeMux I__2993 (
            .O(N__12745),
            .I(N__12741));
    InMux I__2992 (
            .O(N__12744),
            .I(N__12738));
    InMux I__2991 (
            .O(N__12741),
            .I(N__12735));
    LocalMux I__2990 (
            .O(N__12738),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_13 ));
    LocalMux I__2989 (
            .O(N__12735),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_13 ));
    SRMux I__2988 (
            .O(N__12730),
            .I(N__12726));
    SRMux I__2987 (
            .O(N__12729),
            .I(N__12723));
    LocalMux I__2986 (
            .O(N__12726),
            .I(N__12720));
    LocalMux I__2985 (
            .O(N__12723),
            .I(N__12717));
    Span4Mux_h I__2984 (
            .O(N__12720),
            .I(N__12711));
    Span4Mux_h I__2983 (
            .O(N__12717),
            .I(N__12711));
    SRMux I__2982 (
            .O(N__12716),
            .I(N__12708));
    Odrv4 I__2981 (
            .O(N__12711),
            .I(\DUT.uart_inst0.tx_clk_divider_1_sqmuxa_1_i ));
    LocalMux I__2980 (
            .O(N__12708),
            .I(\DUT.uart_inst0.tx_clk_divider_1_sqmuxa_1_i ));
    InMux I__2979 (
            .O(N__12703),
            .I(N__12700));
    LocalMux I__2978 (
            .O(N__12700),
            .I(\DUT.uart_inst0.tx_state_ns_i_i_0_0 ));
    InMux I__2977 (
            .O(N__12697),
            .I(N__12694));
    LocalMux I__2976 (
            .O(N__12694),
            .I(N__12690));
    InMux I__2975 (
            .O(N__12693),
            .I(N__12687));
    Odrv4 I__2974 (
            .O(N__12690),
            .I(\DUT.uart_inst0.N_345_0 ));
    LocalMux I__2973 (
            .O(N__12687),
            .I(\DUT.uart_inst0.N_345_0 ));
    InMux I__2972 (
            .O(N__12682),
            .I(N__12679));
    LocalMux I__2971 (
            .O(N__12679),
            .I(\DUT.uart_inst0.tx_state_ns_i_i_a2_0_1_0 ));
    CascadeMux I__2970 (
            .O(N__12676),
            .I(N__12667));
    CascadeMux I__2969 (
            .O(N__12675),
            .I(N__12663));
    InMux I__2968 (
            .O(N__12674),
            .I(N__12659));
    CascadeMux I__2967 (
            .O(N__12673),
            .I(N__12656));
    InMux I__2966 (
            .O(N__12672),
            .I(N__12650));
    CascadeMux I__2965 (
            .O(N__12671),
            .I(N__12647));
    InMux I__2964 (
            .O(N__12670),
            .I(N__12642));
    InMux I__2963 (
            .O(N__12667),
            .I(N__12639));
    InMux I__2962 (
            .O(N__12666),
            .I(N__12636));
    InMux I__2961 (
            .O(N__12663),
            .I(N__12631));
    InMux I__2960 (
            .O(N__12662),
            .I(N__12631));
    LocalMux I__2959 (
            .O(N__12659),
            .I(N__12628));
    InMux I__2958 (
            .O(N__12656),
            .I(N__12625));
    InMux I__2957 (
            .O(N__12655),
            .I(N__12620));
    InMux I__2956 (
            .O(N__12654),
            .I(N__12620));
    InMux I__2955 (
            .O(N__12653),
            .I(N__12611));
    LocalMux I__2954 (
            .O(N__12650),
            .I(N__12608));
    InMux I__2953 (
            .O(N__12647),
            .I(N__12601));
    InMux I__2952 (
            .O(N__12646),
            .I(N__12601));
    InMux I__2951 (
            .O(N__12645),
            .I(N__12601));
    LocalMux I__2950 (
            .O(N__12642),
            .I(N__12592));
    LocalMux I__2949 (
            .O(N__12639),
            .I(N__12592));
    LocalMux I__2948 (
            .O(N__12636),
            .I(N__12592));
    LocalMux I__2947 (
            .O(N__12631),
            .I(N__12592));
    Span4Mux_v I__2946 (
            .O(N__12628),
            .I(N__12584));
    LocalMux I__2945 (
            .O(N__12625),
            .I(N__12584));
    LocalMux I__2944 (
            .O(N__12620),
            .I(N__12584));
    InMux I__2943 (
            .O(N__12619),
            .I(N__12577));
    InMux I__2942 (
            .O(N__12618),
            .I(N__12577));
    InMux I__2941 (
            .O(N__12617),
            .I(N__12577));
    InMux I__2940 (
            .O(N__12616),
            .I(N__12570));
    InMux I__2939 (
            .O(N__12615),
            .I(N__12570));
    InMux I__2938 (
            .O(N__12614),
            .I(N__12570));
    LocalMux I__2937 (
            .O(N__12611),
            .I(N__12567));
    Span4Mux_v I__2936 (
            .O(N__12608),
            .I(N__12560));
    LocalMux I__2935 (
            .O(N__12601),
            .I(N__12560));
    Span4Mux_v I__2934 (
            .O(N__12592),
            .I(N__12560));
    InMux I__2933 (
            .O(N__12591),
            .I(N__12557));
    Span4Mux_h I__2932 (
            .O(N__12584),
            .I(N__12554));
    LocalMux I__2931 (
            .O(N__12577),
            .I(\DUT.tx_state_0 ));
    LocalMux I__2930 (
            .O(N__12570),
            .I(\DUT.tx_state_0 ));
    Odrv4 I__2929 (
            .O(N__12567),
            .I(\DUT.tx_state_0 ));
    Odrv4 I__2928 (
            .O(N__12560),
            .I(\DUT.tx_state_0 ));
    LocalMux I__2927 (
            .O(N__12557),
            .I(\DUT.tx_state_0 ));
    Odrv4 I__2926 (
            .O(N__12554),
            .I(\DUT.tx_state_0 ));
    CascadeMux I__2925 (
            .O(N__12541),
            .I(N__12536));
    CascadeMux I__2924 (
            .O(N__12540),
            .I(N__12531));
    InMux I__2923 (
            .O(N__12539),
            .I(N__12521));
    InMux I__2922 (
            .O(N__12536),
            .I(N__12521));
    InMux I__2921 (
            .O(N__12535),
            .I(N__12521));
    InMux I__2920 (
            .O(N__12534),
            .I(N__12518));
    InMux I__2919 (
            .O(N__12531),
            .I(N__12513));
    InMux I__2918 (
            .O(N__12530),
            .I(N__12513));
    InMux I__2917 (
            .O(N__12529),
            .I(N__12508));
    InMux I__2916 (
            .O(N__12528),
            .I(N__12508));
    LocalMux I__2915 (
            .O(N__12521),
            .I(N__12505));
    LocalMux I__2914 (
            .O(N__12518),
            .I(N__12502));
    LocalMux I__2913 (
            .O(N__12513),
            .I(N__12499));
    LocalMux I__2912 (
            .O(N__12508),
            .I(N__12496));
    Glb2LocalMux I__2911 (
            .O(N__12505),
            .I(N__12451));
    Glb2LocalMux I__2910 (
            .O(N__12502),
            .I(N__12451));
    Glb2LocalMux I__2909 (
            .O(N__12499),
            .I(N__12451));
    Glb2LocalMux I__2908 (
            .O(N__12496),
            .I(N__12451));
    SRMux I__2907 (
            .O(N__12495),
            .I(N__12451));
    SRMux I__2906 (
            .O(N__12494),
            .I(N__12451));
    SRMux I__2905 (
            .O(N__12493),
            .I(N__12451));
    SRMux I__2904 (
            .O(N__12492),
            .I(N__12451));
    SRMux I__2903 (
            .O(N__12491),
            .I(N__12451));
    SRMux I__2902 (
            .O(N__12490),
            .I(N__12451));
    SRMux I__2901 (
            .O(N__12489),
            .I(N__12451));
    SRMux I__2900 (
            .O(N__12488),
            .I(N__12451));
    SRMux I__2899 (
            .O(N__12487),
            .I(N__12451));
    SRMux I__2898 (
            .O(N__12486),
            .I(N__12451));
    SRMux I__2897 (
            .O(N__12485),
            .I(N__12451));
    SRMux I__2896 (
            .O(N__12484),
            .I(N__12451));
    GlobalMux I__2895 (
            .O(N__12451),
            .I(N__12448));
    gio2CtrlBuf I__2894 (
            .O(N__12448),
            .I(wPllLocked_iso_i_g));
    InMux I__2893 (
            .O(N__12445),
            .I(N__12439));
    InMux I__2892 (
            .O(N__12444),
            .I(N__12436));
    InMux I__2891 (
            .O(N__12443),
            .I(N__12432));
    InMux I__2890 (
            .O(N__12442),
            .I(N__12429));
    LocalMux I__2889 (
            .O(N__12439),
            .I(N__12426));
    LocalMux I__2888 (
            .O(N__12436),
            .I(N__12423));
    InMux I__2887 (
            .O(N__12435),
            .I(N__12420));
    LocalMux I__2886 (
            .O(N__12432),
            .I(N__12417));
    LocalMux I__2885 (
            .O(N__12429),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_2 ));
    Odrv4 I__2884 (
            .O(N__12426),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_2 ));
    Odrv4 I__2883 (
            .O(N__12423),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_2 ));
    LocalMux I__2882 (
            .O(N__12420),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_2 ));
    Odrv4 I__2881 (
            .O(N__12417),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_2 ));
    InMux I__2880 (
            .O(N__12406),
            .I(N__12401));
    CascadeMux I__2879 (
            .O(N__12405),
            .I(N__12397));
    InMux I__2878 (
            .O(N__12404),
            .I(N__12393));
    LocalMux I__2877 (
            .O(N__12401),
            .I(N__12390));
    InMux I__2876 (
            .O(N__12400),
            .I(N__12384));
    InMux I__2875 (
            .O(N__12397),
            .I(N__12379));
    InMux I__2874 (
            .O(N__12396),
            .I(N__12379));
    LocalMux I__2873 (
            .O(N__12393),
            .I(N__12376));
    Span4Mux_v I__2872 (
            .O(N__12390),
            .I(N__12373));
    InMux I__2871 (
            .O(N__12389),
            .I(N__12370));
    InMux I__2870 (
            .O(N__12388),
            .I(N__12365));
    InMux I__2869 (
            .O(N__12387),
            .I(N__12365));
    LocalMux I__2868 (
            .O(N__12384),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_0 ));
    LocalMux I__2867 (
            .O(N__12379),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_0 ));
    Odrv12 I__2866 (
            .O(N__12376),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_0 ));
    Odrv4 I__2865 (
            .O(N__12373),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_0 ));
    LocalMux I__2864 (
            .O(N__12370),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_0 ));
    LocalMux I__2863 (
            .O(N__12365),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_0 ));
    CascadeMux I__2862 (
            .O(N__12352),
            .I(N__12349));
    InMux I__2861 (
            .O(N__12349),
            .I(N__12346));
    LocalMux I__2860 (
            .O(N__12346),
            .I(N__12343));
    Odrv4 I__2859 (
            .O(N__12343),
            .I(\DUT.uart_inst0.tx_bits_remaining_RNO_0Z0Z_3 ));
    InMux I__2858 (
            .O(N__12340),
            .I(N__12334));
    InMux I__2857 (
            .O(N__12339),
            .I(N__12329));
    InMux I__2856 (
            .O(N__12338),
            .I(N__12329));
    CascadeMux I__2855 (
            .O(N__12337),
            .I(N__12325));
    LocalMux I__2854 (
            .O(N__12334),
            .I(N__12312));
    LocalMux I__2853 (
            .O(N__12329),
            .I(N__12312));
    InMux I__2852 (
            .O(N__12328),
            .I(N__12307));
    InMux I__2851 (
            .O(N__12325),
            .I(N__12307));
    InMux I__2850 (
            .O(N__12324),
            .I(N__12304));
    InMux I__2849 (
            .O(N__12323),
            .I(N__12299));
    InMux I__2848 (
            .O(N__12322),
            .I(N__12299));
    InMux I__2847 (
            .O(N__12321),
            .I(N__12296));
    InMux I__2846 (
            .O(N__12320),
            .I(N__12289));
    InMux I__2845 (
            .O(N__12319),
            .I(N__12289));
    InMux I__2844 (
            .O(N__12318),
            .I(N__12289));
    InMux I__2843 (
            .O(N__12317),
            .I(N__12286));
    Span4Mux_v I__2842 (
            .O(N__12312),
            .I(N__12283));
    LocalMux I__2841 (
            .O(N__12307),
            .I(N__12278));
    LocalMux I__2840 (
            .O(N__12304),
            .I(N__12278));
    LocalMux I__2839 (
            .O(N__12299),
            .I(N__12275));
    LocalMux I__2838 (
            .O(N__12296),
            .I(N__12270));
    LocalMux I__2837 (
            .O(N__12289),
            .I(N__12270));
    LocalMux I__2836 (
            .O(N__12286),
            .I(N__12267));
    Span4Mux_h I__2835 (
            .O(N__12283),
            .I(N__12262));
    Span4Mux_v I__2834 (
            .O(N__12278),
            .I(N__12259));
    Span4Mux_h I__2833 (
            .O(N__12275),
            .I(N__12256));
    Span4Mux_v I__2832 (
            .O(N__12270),
            .I(N__12251));
    Span4Mux_h I__2831 (
            .O(N__12267),
            .I(N__12251));
    InMux I__2830 (
            .O(N__12266),
            .I(N__12246));
    InMux I__2829 (
            .O(N__12265),
            .I(N__12246));
    Odrv4 I__2828 (
            .O(N__12262),
            .I(\DUT.tx_state_1 ));
    Odrv4 I__2827 (
            .O(N__12259),
            .I(\DUT.tx_state_1 ));
    Odrv4 I__2826 (
            .O(N__12256),
            .I(\DUT.tx_state_1 ));
    Odrv4 I__2825 (
            .O(N__12251),
            .I(\DUT.tx_state_1 ));
    LocalMux I__2824 (
            .O(N__12246),
            .I(\DUT.tx_state_1 ));
    InMux I__2823 (
            .O(N__12235),
            .I(N__12230));
    InMux I__2822 (
            .O(N__12234),
            .I(N__12225));
    InMux I__2821 (
            .O(N__12233),
            .I(N__12225));
    LocalMux I__2820 (
            .O(N__12230),
            .I(N__12218));
    LocalMux I__2819 (
            .O(N__12225),
            .I(N__12218));
    InMux I__2818 (
            .O(N__12224),
            .I(N__12213));
    InMux I__2817 (
            .O(N__12223),
            .I(N__12210));
    Span4Mux_v I__2816 (
            .O(N__12218),
            .I(N__12207));
    InMux I__2815 (
            .O(N__12217),
            .I(N__12204));
    InMux I__2814 (
            .O(N__12216),
            .I(N__12201));
    LocalMux I__2813 (
            .O(N__12213),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_1 ));
    LocalMux I__2812 (
            .O(N__12210),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_1 ));
    Odrv4 I__2811 (
            .O(N__12207),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_1 ));
    LocalMux I__2810 (
            .O(N__12204),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_1 ));
    LocalMux I__2809 (
            .O(N__12201),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_1 ));
    CascadeMux I__2808 (
            .O(N__12190),
            .I(N__12187));
    InMux I__2807 (
            .O(N__12187),
            .I(N__12184));
    LocalMux I__2806 (
            .O(N__12184),
            .I(N__12181));
    Span4Mux_h I__2805 (
            .O(N__12181),
            .I(N__12178));
    Odrv4 I__2804 (
            .O(N__12178),
            .I(\DUT.uart_inst0.tx_bits_remaining_RNO_0Z0Z_2 ));
    InMux I__2803 (
            .O(N__12175),
            .I(N__12172));
    LocalMux I__2802 (
            .O(N__12172),
            .I(N__12169));
    Odrv12 I__2801 (
            .O(N__12169),
            .I(iRxF_n_c));
    CascadeMux I__2800 (
            .O(N__12166),
            .I(N__12161));
    InMux I__2799 (
            .O(N__12165),
            .I(N__12158));
    InMux I__2798 (
            .O(N__12164),
            .I(N__12155));
    InMux I__2797 (
            .O(N__12161),
            .I(N__12152));
    LocalMux I__2796 (
            .O(N__12158),
            .I(N__12147));
    LocalMux I__2795 (
            .O(N__12155),
            .I(N__12147));
    LocalMux I__2794 (
            .O(N__12152),
            .I(N__12142));
    Sp12to4 I__2793 (
            .O(N__12147),
            .I(N__12142));
    Odrv12 I__2792 (
            .O(N__12142),
            .I(\fifo_inst.ftdi_output_inst.rRxF_nZ0Z_0 ));
    ClkMux I__2791 (
            .O(N__12139),
            .I(N__11944));
    ClkMux I__2790 (
            .O(N__12138),
            .I(N__11944));
    ClkMux I__2789 (
            .O(N__12137),
            .I(N__11944));
    ClkMux I__2788 (
            .O(N__12136),
            .I(N__11944));
    ClkMux I__2787 (
            .O(N__12135),
            .I(N__11944));
    ClkMux I__2786 (
            .O(N__12134),
            .I(N__11944));
    ClkMux I__2785 (
            .O(N__12133),
            .I(N__11944));
    ClkMux I__2784 (
            .O(N__12132),
            .I(N__11944));
    ClkMux I__2783 (
            .O(N__12131),
            .I(N__11944));
    ClkMux I__2782 (
            .O(N__12130),
            .I(N__11944));
    ClkMux I__2781 (
            .O(N__12129),
            .I(N__11944));
    ClkMux I__2780 (
            .O(N__12128),
            .I(N__11944));
    ClkMux I__2779 (
            .O(N__12127),
            .I(N__11944));
    ClkMux I__2778 (
            .O(N__12126),
            .I(N__11944));
    ClkMux I__2777 (
            .O(N__12125),
            .I(N__11944));
    ClkMux I__2776 (
            .O(N__12124),
            .I(N__11944));
    ClkMux I__2775 (
            .O(N__12123),
            .I(N__11944));
    ClkMux I__2774 (
            .O(N__12122),
            .I(N__11944));
    ClkMux I__2773 (
            .O(N__12121),
            .I(N__11944));
    ClkMux I__2772 (
            .O(N__12120),
            .I(N__11944));
    ClkMux I__2771 (
            .O(N__12119),
            .I(N__11944));
    ClkMux I__2770 (
            .O(N__12118),
            .I(N__11944));
    ClkMux I__2769 (
            .O(N__12117),
            .I(N__11944));
    ClkMux I__2768 (
            .O(N__12116),
            .I(N__11944));
    ClkMux I__2767 (
            .O(N__12115),
            .I(N__11944));
    ClkMux I__2766 (
            .O(N__12114),
            .I(N__11944));
    ClkMux I__2765 (
            .O(N__12113),
            .I(N__11944));
    ClkMux I__2764 (
            .O(N__12112),
            .I(N__11944));
    ClkMux I__2763 (
            .O(N__12111),
            .I(N__11944));
    ClkMux I__2762 (
            .O(N__12110),
            .I(N__11944));
    ClkMux I__2761 (
            .O(N__12109),
            .I(N__11944));
    ClkMux I__2760 (
            .O(N__12108),
            .I(N__11944));
    ClkMux I__2759 (
            .O(N__12107),
            .I(N__11944));
    ClkMux I__2758 (
            .O(N__12106),
            .I(N__11944));
    ClkMux I__2757 (
            .O(N__12105),
            .I(N__11944));
    ClkMux I__2756 (
            .O(N__12104),
            .I(N__11944));
    ClkMux I__2755 (
            .O(N__12103),
            .I(N__11944));
    ClkMux I__2754 (
            .O(N__12102),
            .I(N__11944));
    ClkMux I__2753 (
            .O(N__12101),
            .I(N__11944));
    ClkMux I__2752 (
            .O(N__12100),
            .I(N__11944));
    ClkMux I__2751 (
            .O(N__12099),
            .I(N__11944));
    ClkMux I__2750 (
            .O(N__12098),
            .I(N__11944));
    ClkMux I__2749 (
            .O(N__12097),
            .I(N__11944));
    ClkMux I__2748 (
            .O(N__12096),
            .I(N__11944));
    ClkMux I__2747 (
            .O(N__12095),
            .I(N__11944));
    ClkMux I__2746 (
            .O(N__12094),
            .I(N__11944));
    ClkMux I__2745 (
            .O(N__12093),
            .I(N__11944));
    ClkMux I__2744 (
            .O(N__12092),
            .I(N__11944));
    ClkMux I__2743 (
            .O(N__12091),
            .I(N__11944));
    ClkMux I__2742 (
            .O(N__12090),
            .I(N__11944));
    ClkMux I__2741 (
            .O(N__12089),
            .I(N__11944));
    ClkMux I__2740 (
            .O(N__12088),
            .I(N__11944));
    ClkMux I__2739 (
            .O(N__12087),
            .I(N__11944));
    ClkMux I__2738 (
            .O(N__12086),
            .I(N__11944));
    ClkMux I__2737 (
            .O(N__12085),
            .I(N__11944));
    ClkMux I__2736 (
            .O(N__12084),
            .I(N__11944));
    ClkMux I__2735 (
            .O(N__12083),
            .I(N__11944));
    ClkMux I__2734 (
            .O(N__12082),
            .I(N__11944));
    ClkMux I__2733 (
            .O(N__12081),
            .I(N__11944));
    ClkMux I__2732 (
            .O(N__12080),
            .I(N__11944));
    ClkMux I__2731 (
            .O(N__12079),
            .I(N__11944));
    ClkMux I__2730 (
            .O(N__12078),
            .I(N__11944));
    ClkMux I__2729 (
            .O(N__12077),
            .I(N__11944));
    ClkMux I__2728 (
            .O(N__12076),
            .I(N__11944));
    ClkMux I__2727 (
            .O(N__12075),
            .I(N__11944));
    GlobalMux I__2726 (
            .O(N__11944),
            .I(clk_48mhz));
    CascadeMux I__2725 (
            .O(N__11941),
            .I(N__11932));
    CascadeMux I__2724 (
            .O(N__11940),
            .I(N__11926));
    InMux I__2723 (
            .O(N__11939),
            .I(N__11915));
    InMux I__2722 (
            .O(N__11938),
            .I(N__11908));
    InMux I__2721 (
            .O(N__11937),
            .I(N__11908));
    InMux I__2720 (
            .O(N__11936),
            .I(N__11908));
    InMux I__2719 (
            .O(N__11935),
            .I(N__11905));
    InMux I__2718 (
            .O(N__11932),
            .I(N__11898));
    InMux I__2717 (
            .O(N__11931),
            .I(N__11898));
    InMux I__2716 (
            .O(N__11930),
            .I(N__11898));
    InMux I__2715 (
            .O(N__11929),
            .I(N__11893));
    InMux I__2714 (
            .O(N__11926),
            .I(N__11893));
    InMux I__2713 (
            .O(N__11925),
            .I(N__11890));
    InMux I__2712 (
            .O(N__11924),
            .I(N__11887));
    InMux I__2711 (
            .O(N__11923),
            .I(N__11884));
    InMux I__2710 (
            .O(N__11922),
            .I(N__11881));
    InMux I__2709 (
            .O(N__11921),
            .I(N__11878));
    InMux I__2708 (
            .O(N__11920),
            .I(N__11875));
    InMux I__2707 (
            .O(N__11919),
            .I(N__11872));
    InMux I__2706 (
            .O(N__11918),
            .I(N__11869));
    LocalMux I__2705 (
            .O(N__11915),
            .I(N__11863));
    LocalMux I__2704 (
            .O(N__11908),
            .I(N__11859));
    LocalMux I__2703 (
            .O(N__11905),
            .I(N__11856));
    LocalMux I__2702 (
            .O(N__11898),
            .I(N__11853));
    LocalMux I__2701 (
            .O(N__11893),
            .I(N__11850));
    LocalMux I__2700 (
            .O(N__11890),
            .I(N__11840));
    LocalMux I__2699 (
            .O(N__11887),
            .I(N__11837));
    LocalMux I__2698 (
            .O(N__11884),
            .I(N__11833));
    LocalMux I__2697 (
            .O(N__11881),
            .I(N__11829));
    LocalMux I__2696 (
            .O(N__11878),
            .I(N__11826));
    LocalMux I__2695 (
            .O(N__11875),
            .I(N__11823));
    LocalMux I__2694 (
            .O(N__11872),
            .I(N__11820));
    LocalMux I__2693 (
            .O(N__11869),
            .I(N__11817));
    CEMux I__2692 (
            .O(N__11868),
            .I(N__11764));
    CEMux I__2691 (
            .O(N__11867),
            .I(N__11764));
    CEMux I__2690 (
            .O(N__11866),
            .I(N__11764));
    Glb2LocalMux I__2689 (
            .O(N__11863),
            .I(N__11764));
    CEMux I__2688 (
            .O(N__11862),
            .I(N__11764));
    Glb2LocalMux I__2687 (
            .O(N__11859),
            .I(N__11764));
    Glb2LocalMux I__2686 (
            .O(N__11856),
            .I(N__11764));
    Glb2LocalMux I__2685 (
            .O(N__11853),
            .I(N__11764));
    Glb2LocalMux I__2684 (
            .O(N__11850),
            .I(N__11764));
    CEMux I__2683 (
            .O(N__11849),
            .I(N__11764));
    CEMux I__2682 (
            .O(N__11848),
            .I(N__11764));
    CEMux I__2681 (
            .O(N__11847),
            .I(N__11764));
    CEMux I__2680 (
            .O(N__11846),
            .I(N__11764));
    CEMux I__2679 (
            .O(N__11845),
            .I(N__11764));
    CEMux I__2678 (
            .O(N__11844),
            .I(N__11764));
    CEMux I__2677 (
            .O(N__11843),
            .I(N__11764));
    Glb2LocalMux I__2676 (
            .O(N__11840),
            .I(N__11764));
    Glb2LocalMux I__2675 (
            .O(N__11837),
            .I(N__11764));
    CEMux I__2674 (
            .O(N__11836),
            .I(N__11764));
    Glb2LocalMux I__2673 (
            .O(N__11833),
            .I(N__11764));
    CEMux I__2672 (
            .O(N__11832),
            .I(N__11764));
    Glb2LocalMux I__2671 (
            .O(N__11829),
            .I(N__11764));
    Glb2LocalMux I__2670 (
            .O(N__11826),
            .I(N__11764));
    Glb2LocalMux I__2669 (
            .O(N__11823),
            .I(N__11764));
    Glb2LocalMux I__2668 (
            .O(N__11820),
            .I(N__11764));
    Glb2LocalMux I__2667 (
            .O(N__11817),
            .I(N__11764));
    GlobalMux I__2666 (
            .O(N__11764),
            .I(N__11761));
    gio2CtrlBuf I__2665 (
            .O(N__11761),
            .I(wPllLocked_g));
    InMux I__2664 (
            .O(N__11758),
            .I(N__11754));
    InMux I__2663 (
            .O(N__11757),
            .I(N__11751));
    LocalMux I__2662 (
            .O(N__11754),
            .I(N__11748));
    LocalMux I__2661 (
            .O(N__11751),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_4 ));
    Odrv4 I__2660 (
            .O(N__11748),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_4 ));
    InMux I__2659 (
            .O(N__11743),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_3 ));
    InMux I__2658 (
            .O(N__11740),
            .I(N__11736));
    InMux I__2657 (
            .O(N__11739),
            .I(N__11733));
    LocalMux I__2656 (
            .O(N__11736),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_5 ));
    LocalMux I__2655 (
            .O(N__11733),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_5 ));
    InMux I__2654 (
            .O(N__11728),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_4 ));
    InMux I__2653 (
            .O(N__11725),
            .I(N__11721));
    InMux I__2652 (
            .O(N__11724),
            .I(N__11718));
    LocalMux I__2651 (
            .O(N__11721),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_6 ));
    LocalMux I__2650 (
            .O(N__11718),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_6 ));
    InMux I__2649 (
            .O(N__11713),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_5 ));
    InMux I__2648 (
            .O(N__11710),
            .I(N__11706));
    InMux I__2647 (
            .O(N__11709),
            .I(N__11703));
    LocalMux I__2646 (
            .O(N__11706),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_7 ));
    LocalMux I__2645 (
            .O(N__11703),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_7 ));
    InMux I__2644 (
            .O(N__11698),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_6 ));
    InMux I__2643 (
            .O(N__11695),
            .I(N__11691));
    InMux I__2642 (
            .O(N__11694),
            .I(N__11688));
    LocalMux I__2641 (
            .O(N__11691),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_8 ));
    LocalMux I__2640 (
            .O(N__11688),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_8 ));
    InMux I__2639 (
            .O(N__11683),
            .I(bfn_18_20_0_));
    InMux I__2638 (
            .O(N__11680),
            .I(N__11676));
    InMux I__2637 (
            .O(N__11679),
            .I(N__11673));
    LocalMux I__2636 (
            .O(N__11676),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_9 ));
    LocalMux I__2635 (
            .O(N__11673),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_9 ));
    InMux I__2634 (
            .O(N__11668),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_8 ));
    InMux I__2633 (
            .O(N__11665),
            .I(N__11661));
    InMux I__2632 (
            .O(N__11664),
            .I(N__11658));
    LocalMux I__2631 (
            .O(N__11661),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_10 ));
    LocalMux I__2630 (
            .O(N__11658),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_10 ));
    InMux I__2629 (
            .O(N__11653),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_9 ));
    CascadeMux I__2628 (
            .O(N__11650),
            .I(N__11646));
    InMux I__2627 (
            .O(N__11649),
            .I(N__11643));
    InMux I__2626 (
            .O(N__11646),
            .I(N__11640));
    LocalMux I__2625 (
            .O(N__11643),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_11 ));
    LocalMux I__2624 (
            .O(N__11640),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_11 ));
    InMux I__2623 (
            .O(N__11635),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_10 ));
    SRMux I__2622 (
            .O(N__11632),
            .I(N__11629));
    LocalMux I__2621 (
            .O(N__11629),
            .I(N__11626));
    Odrv12 I__2620 (
            .O(N__11626),
            .I(\DUT.uart_inst0.tx_bits_remaining_0_sqmuxa ));
    CascadeMux I__2619 (
            .O(N__11623),
            .I(N__11614));
    InMux I__2618 (
            .O(N__11622),
            .I(N__11611));
    InMux I__2617 (
            .O(N__11621),
            .I(N__11603));
    InMux I__2616 (
            .O(N__11620),
            .I(N__11603));
    InMux I__2615 (
            .O(N__11619),
            .I(N__11599));
    InMux I__2614 (
            .O(N__11618),
            .I(N__11596));
    InMux I__2613 (
            .O(N__11617),
            .I(N__11593));
    InMux I__2612 (
            .O(N__11614),
            .I(N__11590));
    LocalMux I__2611 (
            .O(N__11611),
            .I(N__11587));
    InMux I__2610 (
            .O(N__11610),
            .I(N__11579));
    InMux I__2609 (
            .O(N__11609),
            .I(N__11579));
    InMux I__2608 (
            .O(N__11608),
            .I(N__11579));
    LocalMux I__2607 (
            .O(N__11603),
            .I(N__11576));
    InMux I__2606 (
            .O(N__11602),
            .I(N__11573));
    LocalMux I__2605 (
            .O(N__11599),
            .I(N__11566));
    LocalMux I__2604 (
            .O(N__11596),
            .I(N__11566));
    LocalMux I__2603 (
            .O(N__11593),
            .I(N__11566));
    LocalMux I__2602 (
            .O(N__11590),
            .I(N__11561));
    Span4Mux_h I__2601 (
            .O(N__11587),
            .I(N__11561));
    InMux I__2600 (
            .O(N__11586),
            .I(N__11558));
    LocalMux I__2599 (
            .O(N__11579),
            .I(N__11553));
    Span4Mux_h I__2598 (
            .O(N__11576),
            .I(N__11553));
    LocalMux I__2597 (
            .O(N__11573),
            .I(\DUT.rTransmitZ0 ));
    Odrv12 I__2596 (
            .O(N__11566),
            .I(\DUT.rTransmitZ0 ));
    Odrv4 I__2595 (
            .O(N__11561),
            .I(\DUT.rTransmitZ0 ));
    LocalMux I__2594 (
            .O(N__11558),
            .I(\DUT.rTransmitZ0 ));
    Odrv4 I__2593 (
            .O(N__11553),
            .I(\DUT.rTransmitZ0 ));
    InMux I__2592 (
            .O(N__11542),
            .I(N__11539));
    LocalMux I__2591 (
            .O(N__11539),
            .I(\DUT.uart_inst0.tx_clk_divider_0_sqmuxa ));
    IoInMux I__2590 (
            .O(N__11536),
            .I(N__11532));
    CascadeMux I__2589 (
            .O(N__11535),
            .I(N__11528));
    LocalMux I__2588 (
            .O(N__11532),
            .I(N__11521));
    InMux I__2587 (
            .O(N__11531),
            .I(N__11517));
    InMux I__2586 (
            .O(N__11528),
            .I(N__11512));
    InMux I__2585 (
            .O(N__11527),
            .I(N__11512));
    InMux I__2584 (
            .O(N__11526),
            .I(N__11507));
    InMux I__2583 (
            .O(N__11525),
            .I(N__11507));
    CascadeMux I__2582 (
            .O(N__11524),
            .I(N__11503));
    Span4Mux_s1_v I__2581 (
            .O(N__11521),
            .I(N__11498));
    CascadeMux I__2580 (
            .O(N__11520),
            .I(N__11495));
    LocalMux I__2579 (
            .O(N__11517),
            .I(N__11489));
    LocalMux I__2578 (
            .O(N__11512),
            .I(N__11489));
    LocalMux I__2577 (
            .O(N__11507),
            .I(N__11486));
    InMux I__2576 (
            .O(N__11506),
            .I(N__11483));
    InMux I__2575 (
            .O(N__11503),
            .I(N__11478));
    InMux I__2574 (
            .O(N__11502),
            .I(N__11478));
    InMux I__2573 (
            .O(N__11501),
            .I(N__11475));
    Sp12to4 I__2572 (
            .O(N__11498),
            .I(N__11472));
    InMux I__2571 (
            .O(N__11495),
            .I(N__11469));
    InMux I__2570 (
            .O(N__11494),
            .I(N__11466));
    Span4Mux_v I__2569 (
            .O(N__11489),
            .I(N__11463));
    Span4Mux_v I__2568 (
            .O(N__11486),
            .I(N__11460));
    LocalMux I__2567 (
            .O(N__11483),
            .I(N__11457));
    LocalMux I__2566 (
            .O(N__11478),
            .I(N__11454));
    LocalMux I__2565 (
            .O(N__11475),
            .I(N__11451));
    Span12Mux_h I__2564 (
            .O(N__11472),
            .I(N__11448));
    LocalMux I__2563 (
            .O(N__11469),
            .I(N__11445));
    LocalMux I__2562 (
            .O(N__11466),
            .I(N__11442));
    Span4Mux_h I__2561 (
            .O(N__11463),
            .I(N__11435));
    Span4Mux_h I__2560 (
            .O(N__11460),
            .I(N__11435));
    Span4Mux_v I__2559 (
            .O(N__11457),
            .I(N__11435));
    Span4Mux_v I__2558 (
            .O(N__11454),
            .I(N__11430));
    Span4Mux_v I__2557 (
            .O(N__11451),
            .I(N__11430));
    Span12Mux_v I__2556 (
            .O(N__11448),
            .I(N__11427));
    Span12Mux_v I__2555 (
            .O(N__11445),
            .I(N__11424));
    Span12Mux_h I__2554 (
            .O(N__11442),
            .I(N__11417));
    Sp12to4 I__2553 (
            .O(N__11435),
            .I(N__11417));
    Sp12to4 I__2552 (
            .O(N__11430),
            .I(N__11417));
    Span12Mux_v I__2551 (
            .O(N__11427),
            .I(N__11412));
    Span12Mux_h I__2550 (
            .O(N__11424),
            .I(N__11412));
    Span12Mux_h I__2549 (
            .O(N__11417),
            .I(N__11409));
    Odrv12 I__2548 (
            .O(N__11412),
            .I(wPllLocked));
    Odrv12 I__2547 (
            .O(N__11409),
            .I(wPllLocked));
    CascadeMux I__2546 (
            .O(N__11404),
            .I(\DUT.uart_inst0.tx_clk_divider_0_sqmuxa_cascade_ ));
    InMux I__2545 (
            .O(N__11401),
            .I(N__11389));
    InMux I__2544 (
            .O(N__11400),
            .I(N__11383));
    InMux I__2543 (
            .O(N__11399),
            .I(N__11383));
    InMux I__2542 (
            .O(N__11398),
            .I(N__11380));
    InMux I__2541 (
            .O(N__11397),
            .I(N__11377));
    InMux I__2540 (
            .O(N__11396),
            .I(N__11372));
    InMux I__2539 (
            .O(N__11395),
            .I(N__11363));
    InMux I__2538 (
            .O(N__11394),
            .I(N__11363));
    InMux I__2537 (
            .O(N__11393),
            .I(N__11363));
    InMux I__2536 (
            .O(N__11392),
            .I(N__11363));
    LocalMux I__2535 (
            .O(N__11389),
            .I(N__11360));
    InMux I__2534 (
            .O(N__11388),
            .I(N__11357));
    LocalMux I__2533 (
            .O(N__11383),
            .I(N__11352));
    LocalMux I__2532 (
            .O(N__11380),
            .I(N__11352));
    LocalMux I__2531 (
            .O(N__11377),
            .I(N__11349));
    InMux I__2530 (
            .O(N__11376),
            .I(N__11344));
    InMux I__2529 (
            .O(N__11375),
            .I(N__11344));
    LocalMux I__2528 (
            .O(N__11372),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0 ));
    LocalMux I__2527 (
            .O(N__11363),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0 ));
    Odrv4 I__2526 (
            .O(N__11360),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0 ));
    LocalMux I__2525 (
            .O(N__11357),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0 ));
    Odrv4 I__2524 (
            .O(N__11352),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0 ));
    Odrv4 I__2523 (
            .O(N__11349),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0 ));
    LocalMux I__2522 (
            .O(N__11344),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0 ));
    InMux I__2521 (
            .O(N__11329),
            .I(N__11323));
    InMux I__2520 (
            .O(N__11328),
            .I(N__11323));
    LocalMux I__2519 (
            .O(N__11323),
            .I(N__11319));
    InMux I__2518 (
            .O(N__11322),
            .I(N__11316));
    Odrv4 I__2517 (
            .O(N__11319),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0 ));
    LocalMux I__2516 (
            .O(N__11316),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0 ));
    InMux I__2515 (
            .O(N__11311),
            .I(N__11308));
    LocalMux I__2514 (
            .O(N__11308),
            .I(N__11304));
    InMux I__2513 (
            .O(N__11307),
            .I(N__11301));
    Odrv4 I__2512 (
            .O(N__11304),
            .I(\fifo_inst.ftdi_output_inst.rRxF_nZ0Z_1 ));
    LocalMux I__2511 (
            .O(N__11301),
            .I(\fifo_inst.ftdi_output_inst.rRxF_nZ0Z_1 ));
    InMux I__2510 (
            .O(N__11296),
            .I(N__11293));
    LocalMux I__2509 (
            .O(N__11293),
            .I(N__11289));
    InMux I__2508 (
            .O(N__11292),
            .I(N__11286));
    Odrv12 I__2507 (
            .O(N__11289),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1 ));
    LocalMux I__2506 (
            .O(N__11286),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1 ));
    InMux I__2505 (
            .O(N__11281),
            .I(N__11278));
    LocalMux I__2504 (
            .O(N__11278),
            .I(N__11273));
    InMux I__2503 (
            .O(N__11277),
            .I(N__11270));
    InMux I__2502 (
            .O(N__11276),
            .I(N__11267));
    Span4Mux_h I__2501 (
            .O(N__11273),
            .I(N__11262));
    LocalMux I__2500 (
            .O(N__11270),
            .I(N__11262));
    LocalMux I__2499 (
            .O(N__11267),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_0 ));
    Odrv4 I__2498 (
            .O(N__11262),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_0 ));
    InMux I__2497 (
            .O(N__11257),
            .I(N__11254));
    LocalMux I__2496 (
            .O(N__11254),
            .I(N__11250));
    InMux I__2495 (
            .O(N__11253),
            .I(N__11247));
    Span4Mux_v I__2494 (
            .O(N__11250),
            .I(N__11244));
    LocalMux I__2493 (
            .O(N__11247),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_1 ));
    Odrv4 I__2492 (
            .O(N__11244),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_1 ));
    InMux I__2491 (
            .O(N__11239),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_0 ));
    CascadeMux I__2490 (
            .O(N__11236),
            .I(N__11232));
    InMux I__2489 (
            .O(N__11235),
            .I(N__11229));
    InMux I__2488 (
            .O(N__11232),
            .I(N__11226));
    LocalMux I__2487 (
            .O(N__11229),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_2 ));
    LocalMux I__2486 (
            .O(N__11226),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_2 ));
    InMux I__2485 (
            .O(N__11221),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_1 ));
    InMux I__2484 (
            .O(N__11218),
            .I(N__11214));
    InMux I__2483 (
            .O(N__11217),
            .I(N__11211));
    LocalMux I__2482 (
            .O(N__11214),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_3 ));
    LocalMux I__2481 (
            .O(N__11211),
            .I(\DUT.uart_inst0.tx_clk_dividerZ0Z_3 ));
    InMux I__2480 (
            .O(N__11206),
            .I(\DUT.uart_inst0.tx_clk_divider_cry_2 ));
    CascadeMux I__2479 (
            .O(N__11203),
            .I(N__11197));
    InMux I__2478 (
            .O(N__11202),
            .I(N__11191));
    InMux I__2477 (
            .O(N__11201),
            .I(N__11182));
    InMux I__2476 (
            .O(N__11200),
            .I(N__11182));
    InMux I__2475 (
            .O(N__11197),
            .I(N__11182));
    InMux I__2474 (
            .O(N__11196),
            .I(N__11182));
    InMux I__2473 (
            .O(N__11195),
            .I(N__11169));
    InMux I__2472 (
            .O(N__11194),
            .I(N__11169));
    LocalMux I__2471 (
            .O(N__11191),
            .I(N__11164));
    LocalMux I__2470 (
            .O(N__11182),
            .I(N__11164));
    CascadeMux I__2469 (
            .O(N__11181),
            .I(N__11157));
    CascadeMux I__2468 (
            .O(N__11180),
            .I(N__11153));
    CascadeMux I__2467 (
            .O(N__11179),
            .I(N__11150));
    CascadeMux I__2466 (
            .O(N__11178),
            .I(N__11147));
    InMux I__2465 (
            .O(N__11177),
            .I(N__11138));
    InMux I__2464 (
            .O(N__11176),
            .I(N__11138));
    InMux I__2463 (
            .O(N__11175),
            .I(N__11138));
    InMux I__2462 (
            .O(N__11174),
            .I(N__11135));
    LocalMux I__2461 (
            .O(N__11169),
            .I(N__11132));
    Span4Mux_h I__2460 (
            .O(N__11164),
            .I(N__11129));
    InMux I__2459 (
            .O(N__11163),
            .I(N__11114));
    InMux I__2458 (
            .O(N__11162),
            .I(N__11114));
    InMux I__2457 (
            .O(N__11161),
            .I(N__11114));
    InMux I__2456 (
            .O(N__11160),
            .I(N__11114));
    InMux I__2455 (
            .O(N__11157),
            .I(N__11114));
    InMux I__2454 (
            .O(N__11156),
            .I(N__11114));
    InMux I__2453 (
            .O(N__11153),
            .I(N__11114));
    InMux I__2452 (
            .O(N__11150),
            .I(N__11105));
    InMux I__2451 (
            .O(N__11147),
            .I(N__11105));
    InMux I__2450 (
            .O(N__11146),
            .I(N__11105));
    InMux I__2449 (
            .O(N__11145),
            .I(N__11105));
    LocalMux I__2448 (
            .O(N__11138),
            .I(N__11102));
    LocalMux I__2447 (
            .O(N__11135),
            .I(N__11097));
    Span4Mux_h I__2446 (
            .O(N__11132),
            .I(N__11097));
    Odrv4 I__2445 (
            .O(N__11129),
            .I(\DUT.uart_inst0.N_72 ));
    LocalMux I__2444 (
            .O(N__11114),
            .I(\DUT.uart_inst0.N_72 ));
    LocalMux I__2443 (
            .O(N__11105),
            .I(\DUT.uart_inst0.N_72 ));
    Odrv12 I__2442 (
            .O(N__11102),
            .I(\DUT.uart_inst0.N_72 ));
    Odrv4 I__2441 (
            .O(N__11097),
            .I(\DUT.uart_inst0.N_72 ));
    InMux I__2440 (
            .O(N__11086),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_16 ));
    CascadeMux I__2439 (
            .O(N__11083),
            .I(N__11079));
    InMux I__2438 (
            .O(N__11082),
            .I(N__11076));
    InMux I__2437 (
            .O(N__11079),
            .I(N__11073));
    LocalMux I__2436 (
            .O(N__11076),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_17 ));
    LocalMux I__2435 (
            .O(N__11073),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_17 ));
    CascadeMux I__2434 (
            .O(N__11068),
            .I(N__11065));
    InMux I__2433 (
            .O(N__11065),
            .I(N__11062));
    LocalMux I__2432 (
            .O(N__11062),
            .I(N__11058));
    CascadeMux I__2431 (
            .O(N__11061),
            .I(N__11055));
    Span4Mux_v I__2430 (
            .O(N__11058),
            .I(N__11052));
    InMux I__2429 (
            .O(N__11055),
            .I(N__11049));
    Odrv4 I__2428 (
            .O(N__11052),
            .I(\fifo_inst.wRamRdAddr_2 ));
    LocalMux I__2427 (
            .O(N__11049),
            .I(\fifo_inst.wRamRdAddr_2 ));
    InMux I__2426 (
            .O(N__11044),
            .I(N__11040));
    CascadeMux I__2425 (
            .O(N__11043),
            .I(N__11037));
    LocalMux I__2424 (
            .O(N__11040),
            .I(N__11031));
    InMux I__2423 (
            .O(N__11037),
            .I(N__11026));
    InMux I__2422 (
            .O(N__11036),
            .I(N__11026));
    InMux I__2421 (
            .O(N__11035),
            .I(N__11021));
    InMux I__2420 (
            .O(N__11034),
            .I(N__11021));
    Odrv4 I__2419 (
            .O(N__11031),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4 ));
    LocalMux I__2418 (
            .O(N__11026),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4 ));
    LocalMux I__2417 (
            .O(N__11021),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4 ));
    InMux I__2416 (
            .O(N__11014),
            .I(N__11006));
    InMux I__2415 (
            .O(N__11013),
            .I(N__11006));
    InMux I__2414 (
            .O(N__11012),
            .I(N__11000));
    InMux I__2413 (
            .O(N__11011),
            .I(N__11000));
    LocalMux I__2412 (
            .O(N__11006),
            .I(N__10997));
    InMux I__2411 (
            .O(N__11005),
            .I(N__10994));
    LocalMux I__2410 (
            .O(N__11000),
            .I(N__10991));
    Span4Mux_h I__2409 (
            .O(N__10997),
            .I(N__10988));
    LocalMux I__2408 (
            .O(N__10994),
            .I(\fifo_inst.ftdi_output_inst.rWrDelayZ0 ));
    Odrv4 I__2407 (
            .O(N__10991),
            .I(\fifo_inst.ftdi_output_inst.rWrDelayZ0 ));
    Odrv4 I__2406 (
            .O(N__10988),
            .I(\fifo_inst.ftdi_output_inst.rWrDelayZ0 ));
    InMux I__2405 (
            .O(N__10981),
            .I(N__10978));
    LocalMux I__2404 (
            .O(N__10978),
            .I(\fifo_inst.ftdi_output_inst.N_3_0 ));
    CascadeMux I__2403 (
            .O(N__10975),
            .I(N__10972));
    InMux I__2402 (
            .O(N__10972),
            .I(N__10969));
    LocalMux I__2401 (
            .O(N__10969),
            .I(N__10966));
    Span4Mux_v I__2400 (
            .O(N__10966),
            .I(N__10960));
    InMux I__2399 (
            .O(N__10965),
            .I(N__10953));
    InMux I__2398 (
            .O(N__10964),
            .I(N__10953));
    InMux I__2397 (
            .O(N__10963),
            .I(N__10953));
    Odrv4 I__2396 (
            .O(N__10960),
            .I(\fifo_inst.wRamRdAddr_0 ));
    LocalMux I__2395 (
            .O(N__10953),
            .I(\fifo_inst.wRamRdAddr_0 ));
    CascadeMux I__2394 (
            .O(N__10948),
            .I(\fifo_inst.ftdi_output_inst.N_3_0_cascade_ ));
    CascadeMux I__2393 (
            .O(N__10945),
            .I(N__10942));
    InMux I__2392 (
            .O(N__10942),
            .I(N__10939));
    LocalMux I__2391 (
            .O(N__10939),
            .I(N__10936));
    Span4Mux_v I__2390 (
            .O(N__10936),
            .I(N__10933));
    Span4Mux_v I__2389 (
            .O(N__10933),
            .I(N__10928));
    InMux I__2388 (
            .O(N__10932),
            .I(N__10923));
    InMux I__2387 (
            .O(N__10931),
            .I(N__10923));
    Odrv4 I__2386 (
            .O(N__10928),
            .I(\fifo_inst.wRamRdAddr_1 ));
    LocalMux I__2385 (
            .O(N__10923),
            .I(\fifo_inst.wRamRdAddr_1 ));
    InMux I__2384 (
            .O(N__10918),
            .I(N__10915));
    LocalMux I__2383 (
            .O(N__10915),
            .I(N__10912));
    Span4Mux_h I__2382 (
            .O(N__10912),
            .I(N__10909));
    Odrv4 I__2381 (
            .O(N__10909),
            .I(\DUT.uart_inst0.tx_state_ns_i_i_a2_0_0_0 ));
    CascadeMux I__2380 (
            .O(N__10906),
            .I(N__10901));
    InMux I__2379 (
            .O(N__10905),
            .I(N__10893));
    InMux I__2378 (
            .O(N__10904),
            .I(N__10890));
    InMux I__2377 (
            .O(N__10901),
            .I(N__10883));
    InMux I__2376 (
            .O(N__10900),
            .I(N__10883));
    InMux I__2375 (
            .O(N__10899),
            .I(N__10883));
    InMux I__2374 (
            .O(N__10898),
            .I(N__10878));
    InMux I__2373 (
            .O(N__10897),
            .I(N__10878));
    InMux I__2372 (
            .O(N__10896),
            .I(N__10875));
    LocalMux I__2371 (
            .O(N__10893),
            .I(N__10872));
    LocalMux I__2370 (
            .O(N__10890),
            .I(N__10864));
    LocalMux I__2369 (
            .O(N__10883),
            .I(N__10864));
    LocalMux I__2368 (
            .O(N__10878),
            .I(N__10859));
    LocalMux I__2367 (
            .O(N__10875),
            .I(N__10859));
    Span4Mux_h I__2366 (
            .O(N__10872),
            .I(N__10856));
    InMux I__2365 (
            .O(N__10871),
            .I(N__10849));
    InMux I__2364 (
            .O(N__10870),
            .I(N__10849));
    InMux I__2363 (
            .O(N__10869),
            .I(N__10849));
    Span4Mux_v I__2362 (
            .O(N__10864),
            .I(N__10846));
    Span4Mux_h I__2361 (
            .O(N__10859),
            .I(N__10843));
    Span4Mux_v I__2360 (
            .O(N__10856),
            .I(N__10840));
    LocalMux I__2359 (
            .O(N__10849),
            .I(\DUT.uart_inst0.tx_state_0_sqmuxa_i_0 ));
    Odrv4 I__2358 (
            .O(N__10846),
            .I(\DUT.uart_inst0.tx_state_0_sqmuxa_i_0 ));
    Odrv4 I__2357 (
            .O(N__10843),
            .I(\DUT.uart_inst0.tx_state_0_sqmuxa_i_0 ));
    Odrv4 I__2356 (
            .O(N__10840),
            .I(\DUT.uart_inst0.tx_state_0_sqmuxa_i_0 ));
    InMux I__2355 (
            .O(N__10831),
            .I(N__10827));
    IoInMux I__2354 (
            .O(N__10830),
            .I(N__10824));
    LocalMux I__2353 (
            .O(N__10827),
            .I(N__10821));
    LocalMux I__2352 (
            .O(N__10824),
            .I(N__10818));
    Span4Mux_v I__2351 (
            .O(N__10821),
            .I(N__10815));
    Span12Mux_s10_v I__2350 (
            .O(N__10818),
            .I(N__10812));
    Span4Mux_h I__2349 (
            .O(N__10815),
            .I(N__10809));
    Odrv12 I__2348 (
            .O(N__10812),
            .I(wPllLocked_iso_i));
    Odrv4 I__2347 (
            .O(N__10809),
            .I(wPllLocked_iso_i));
    CEMux I__2346 (
            .O(N__10804),
            .I(N__10801));
    LocalMux I__2345 (
            .O(N__10801),
            .I(\DUT.uart_inst0.N_345_0_0 ));
    InMux I__2344 (
            .O(N__10798),
            .I(N__10793));
    InMux I__2343 (
            .O(N__10797),
            .I(N__10790));
    InMux I__2342 (
            .O(N__10796),
            .I(N__10787));
    LocalMux I__2341 (
            .O(N__10793),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_9 ));
    LocalMux I__2340 (
            .O(N__10790),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_9 ));
    LocalMux I__2339 (
            .O(N__10787),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_9 ));
    InMux I__2338 (
            .O(N__10780),
            .I(N__10777));
    LocalMux I__2337 (
            .O(N__10777),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO ));
    InMux I__2336 (
            .O(N__10774),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_8 ));
    InMux I__2335 (
            .O(N__10771),
            .I(N__10766));
    InMux I__2334 (
            .O(N__10770),
            .I(N__10761));
    InMux I__2333 (
            .O(N__10769),
            .I(N__10761));
    LocalMux I__2332 (
            .O(N__10766),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_10 ));
    LocalMux I__2331 (
            .O(N__10761),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_10 ));
    InMux I__2330 (
            .O(N__10756),
            .I(N__10753));
    LocalMux I__2329 (
            .O(N__10753),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO ));
    InMux I__2328 (
            .O(N__10750),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_9 ));
    InMux I__2327 (
            .O(N__10747),
            .I(N__10742));
    InMux I__2326 (
            .O(N__10746),
            .I(N__10737));
    InMux I__2325 (
            .O(N__10745),
            .I(N__10737));
    LocalMux I__2324 (
            .O(N__10742),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_11 ));
    LocalMux I__2323 (
            .O(N__10737),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_11 ));
    InMux I__2322 (
            .O(N__10732),
            .I(N__10729));
    LocalMux I__2321 (
            .O(N__10729),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO ));
    InMux I__2320 (
            .O(N__10726),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_10 ));
    CascadeMux I__2319 (
            .O(N__10723),
            .I(N__10718));
    InMux I__2318 (
            .O(N__10722),
            .I(N__10715));
    InMux I__2317 (
            .O(N__10721),
            .I(N__10710));
    InMux I__2316 (
            .O(N__10718),
            .I(N__10710));
    LocalMux I__2315 (
            .O(N__10715),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_12 ));
    LocalMux I__2314 (
            .O(N__10710),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_12 ));
    InMux I__2313 (
            .O(N__10705),
            .I(N__10702));
    LocalMux I__2312 (
            .O(N__10702),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO ));
    InMux I__2311 (
            .O(N__10699),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_11 ));
    InMux I__2310 (
            .O(N__10696),
            .I(N__10691));
    InMux I__2309 (
            .O(N__10695),
            .I(N__10686));
    InMux I__2308 (
            .O(N__10694),
            .I(N__10686));
    LocalMux I__2307 (
            .O(N__10691),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_13 ));
    LocalMux I__2306 (
            .O(N__10686),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_13 ));
    CascadeMux I__2305 (
            .O(N__10681),
            .I(N__10678));
    InMux I__2304 (
            .O(N__10678),
            .I(N__10675));
    LocalMux I__2303 (
            .O(N__10675),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO ));
    InMux I__2302 (
            .O(N__10672),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_12 ));
    InMux I__2301 (
            .O(N__10669),
            .I(N__10664));
    InMux I__2300 (
            .O(N__10668),
            .I(N__10661));
    InMux I__2299 (
            .O(N__10667),
            .I(N__10658));
    LocalMux I__2298 (
            .O(N__10664),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_14 ));
    LocalMux I__2297 (
            .O(N__10661),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_14 ));
    LocalMux I__2296 (
            .O(N__10658),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_14 ));
    InMux I__2295 (
            .O(N__10651),
            .I(N__10648));
    LocalMux I__2294 (
            .O(N__10648),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO ));
    InMux I__2293 (
            .O(N__10645),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_13 ));
    InMux I__2292 (
            .O(N__10642),
            .I(N__10637));
    InMux I__2291 (
            .O(N__10641),
            .I(N__10632));
    InMux I__2290 (
            .O(N__10640),
            .I(N__10632));
    LocalMux I__2289 (
            .O(N__10637),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_15 ));
    LocalMux I__2288 (
            .O(N__10632),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_15 ));
    CascadeMux I__2287 (
            .O(N__10627),
            .I(N__10624));
    InMux I__2286 (
            .O(N__10624),
            .I(N__10621));
    LocalMux I__2285 (
            .O(N__10621),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO ));
    InMux I__2284 (
            .O(N__10618),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_14 ));
    InMux I__2283 (
            .O(N__10615),
            .I(N__10610));
    InMux I__2282 (
            .O(N__10614),
            .I(N__10607));
    InMux I__2281 (
            .O(N__10613),
            .I(N__10604));
    LocalMux I__2280 (
            .O(N__10610),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_16 ));
    LocalMux I__2279 (
            .O(N__10607),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_16 ));
    LocalMux I__2278 (
            .O(N__10604),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_16 ));
    InMux I__2277 (
            .O(N__10597),
            .I(N__10594));
    LocalMux I__2276 (
            .O(N__10594),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO ));
    InMux I__2275 (
            .O(N__10591),
            .I(bfn_18_15_0_));
    InMux I__2274 (
            .O(N__10588),
            .I(N__10583));
    InMux I__2273 (
            .O(N__10587),
            .I(N__10580));
    InMux I__2272 (
            .O(N__10586),
            .I(N__10577));
    LocalMux I__2271 (
            .O(N__10583),
            .I(\DUT.uart_inst0.rx_clk_dividerZ1Z_1 ));
    LocalMux I__2270 (
            .O(N__10580),
            .I(\DUT.uart_inst0.rx_clk_dividerZ1Z_1 ));
    LocalMux I__2269 (
            .O(N__10577),
            .I(\DUT.uart_inst0.rx_clk_dividerZ1Z_1 ));
    InMux I__2268 (
            .O(N__10570),
            .I(N__10567));
    LocalMux I__2267 (
            .O(N__10567),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO ));
    InMux I__2266 (
            .O(N__10564),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_0 ));
    InMux I__2265 (
            .O(N__10561),
            .I(N__10558));
    LocalMux I__2264 (
            .O(N__10558),
            .I(N__10553));
    InMux I__2263 (
            .O(N__10557),
            .I(N__10548));
    InMux I__2262 (
            .O(N__10556),
            .I(N__10548));
    Odrv4 I__2261 (
            .O(N__10553),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_2 ));
    LocalMux I__2260 (
            .O(N__10548),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_2 ));
    InMux I__2259 (
            .O(N__10543),
            .I(N__10540));
    LocalMux I__2258 (
            .O(N__10540),
            .I(N__10537));
    Odrv4 I__2257 (
            .O(N__10537),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO ));
    InMux I__2256 (
            .O(N__10534),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_1 ));
    InMux I__2255 (
            .O(N__10531),
            .I(N__10527));
    CascadeMux I__2254 (
            .O(N__10530),
            .I(N__10523));
    LocalMux I__2253 (
            .O(N__10527),
            .I(N__10520));
    InMux I__2252 (
            .O(N__10526),
            .I(N__10517));
    InMux I__2251 (
            .O(N__10523),
            .I(N__10514));
    Span4Mux_h I__2250 (
            .O(N__10520),
            .I(N__10511));
    LocalMux I__2249 (
            .O(N__10517),
            .I(N__10508));
    LocalMux I__2248 (
            .O(N__10514),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_3 ));
    Odrv4 I__2247 (
            .O(N__10511),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_3 ));
    Odrv4 I__2246 (
            .O(N__10508),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_3 ));
    InMux I__2245 (
            .O(N__10501),
            .I(N__10498));
    LocalMux I__2244 (
            .O(N__10498),
            .I(N__10495));
    Span4Mux_v I__2243 (
            .O(N__10495),
            .I(N__10492));
    Odrv4 I__2242 (
            .O(N__10492),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_2_THRU_CO ));
    InMux I__2241 (
            .O(N__10489),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_2 ));
    CascadeMux I__2240 (
            .O(N__10486),
            .I(N__10481));
    CascadeMux I__2239 (
            .O(N__10485),
            .I(N__10478));
    InMux I__2238 (
            .O(N__10484),
            .I(N__10475));
    InMux I__2237 (
            .O(N__10481),
            .I(N__10472));
    InMux I__2236 (
            .O(N__10478),
            .I(N__10469));
    LocalMux I__2235 (
            .O(N__10475),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_4 ));
    LocalMux I__2234 (
            .O(N__10472),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_4 ));
    LocalMux I__2233 (
            .O(N__10469),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_4 ));
    InMux I__2232 (
            .O(N__10462),
            .I(N__10459));
    LocalMux I__2231 (
            .O(N__10459),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO ));
    InMux I__2230 (
            .O(N__10456),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_3 ));
    InMux I__2229 (
            .O(N__10453),
            .I(N__10448));
    InMux I__2228 (
            .O(N__10452),
            .I(N__10445));
    InMux I__2227 (
            .O(N__10451),
            .I(N__10442));
    LocalMux I__2226 (
            .O(N__10448),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_5 ));
    LocalMux I__2225 (
            .O(N__10445),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_5 ));
    LocalMux I__2224 (
            .O(N__10442),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_5 ));
    InMux I__2223 (
            .O(N__10435),
            .I(N__10432));
    LocalMux I__2222 (
            .O(N__10432),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_4_THRU_CO ));
    InMux I__2221 (
            .O(N__10429),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_4 ));
    InMux I__2220 (
            .O(N__10426),
            .I(N__10421));
    InMux I__2219 (
            .O(N__10425),
            .I(N__10418));
    InMux I__2218 (
            .O(N__10424),
            .I(N__10415));
    LocalMux I__2217 (
            .O(N__10421),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_6 ));
    LocalMux I__2216 (
            .O(N__10418),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_6 ));
    LocalMux I__2215 (
            .O(N__10415),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_6 ));
    InMux I__2214 (
            .O(N__10408),
            .I(N__10405));
    LocalMux I__2213 (
            .O(N__10405),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_5_THRU_CO ));
    InMux I__2212 (
            .O(N__10402),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_5 ));
    InMux I__2211 (
            .O(N__10399),
            .I(N__10394));
    InMux I__2210 (
            .O(N__10398),
            .I(N__10391));
    InMux I__2209 (
            .O(N__10397),
            .I(N__10388));
    LocalMux I__2208 (
            .O(N__10394),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_7 ));
    LocalMux I__2207 (
            .O(N__10391),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_7 ));
    LocalMux I__2206 (
            .O(N__10388),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_7 ));
    InMux I__2205 (
            .O(N__10381),
            .I(N__10378));
    LocalMux I__2204 (
            .O(N__10378),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO ));
    InMux I__2203 (
            .O(N__10375),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_6 ));
    CascadeMux I__2202 (
            .O(N__10372),
            .I(N__10368));
    InMux I__2201 (
            .O(N__10371),
            .I(N__10364));
    InMux I__2200 (
            .O(N__10368),
            .I(N__10361));
    InMux I__2199 (
            .O(N__10367),
            .I(N__10358));
    LocalMux I__2198 (
            .O(N__10364),
            .I(N__10355));
    LocalMux I__2197 (
            .O(N__10361),
            .I(N__10352));
    LocalMux I__2196 (
            .O(N__10358),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_8 ));
    Odrv4 I__2195 (
            .O(N__10355),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_8 ));
    Odrv4 I__2194 (
            .O(N__10352),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_8 ));
    InMux I__2193 (
            .O(N__10345),
            .I(N__10342));
    LocalMux I__2192 (
            .O(N__10342),
            .I(N__10339));
    Odrv4 I__2191 (
            .O(N__10339),
            .I(\DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO ));
    InMux I__2190 (
            .O(N__10336),
            .I(bfn_18_14_0_));
    CascadeMux I__2189 (
            .O(N__10333),
            .I(N__10328));
    InMux I__2188 (
            .O(N__10332),
            .I(N__10324));
    CascadeMux I__2187 (
            .O(N__10331),
            .I(N__10321));
    InMux I__2186 (
            .O(N__10328),
            .I(N__10318));
    InMux I__2185 (
            .O(N__10327),
            .I(N__10315));
    LocalMux I__2184 (
            .O(N__10324),
            .I(N__10312));
    InMux I__2183 (
            .O(N__10321),
            .I(N__10309));
    LocalMux I__2182 (
            .O(N__10318),
            .I(N__10306));
    LocalMux I__2181 (
            .O(N__10315),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_3 ));
    Odrv4 I__2180 (
            .O(N__10312),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_3 ));
    LocalMux I__2179 (
            .O(N__10309),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_3 ));
    Odrv4 I__2178 (
            .O(N__10306),
            .I(\DUT.uart_inst0.tx_bits_remainingZ0Z_3 ));
    CascadeMux I__2177 (
            .O(N__10297),
            .I(\DUT.uart_inst0.tx_state_ns_i_i_a2_0_0_0_cascade_ ));
    InMux I__2176 (
            .O(N__10294),
            .I(N__10291));
    LocalMux I__2175 (
            .O(N__10291),
            .I(\DUT.uart_inst0.g0_i_a4_1_0 ));
    InMux I__2174 (
            .O(N__10288),
            .I(N__10285));
    LocalMux I__2173 (
            .O(N__10285),
            .I(N__10282));
    Span4Mux_h I__2172 (
            .O(N__10282),
            .I(N__10279));
    Odrv4 I__2171 (
            .O(N__10279),
            .I(\DUT.uart_inst0.d_N_5_mux ));
    InMux I__2170 (
            .O(N__10276),
            .I(N__10272));
    InMux I__2169 (
            .O(N__10275),
            .I(N__10269));
    LocalMux I__2168 (
            .O(N__10272),
            .I(N__10262));
    LocalMux I__2167 (
            .O(N__10269),
            .I(N__10262));
    InMux I__2166 (
            .O(N__10268),
            .I(N__10259));
    InMux I__2165 (
            .O(N__10267),
            .I(N__10256));
    Span12Mux_h I__2164 (
            .O(N__10262),
            .I(N__10249));
    LocalMux I__2163 (
            .O(N__10259),
            .I(N__10249));
    LocalMux I__2162 (
            .O(N__10256),
            .I(N__10249));
    Odrv12 I__2161 (
            .O(N__10249),
            .I(rTxByteZ0Z_3));
    InMux I__2160 (
            .O(N__10246),
            .I(N__10243));
    LocalMux I__2159 (
            .O(N__10243),
            .I(N__10240));
    Odrv4 I__2158 (
            .O(N__10240),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_3 ));
    CEMux I__2157 (
            .O(N__10237),
            .I(N__10234));
    LocalMux I__2156 (
            .O(N__10234),
            .I(N__10230));
    CEMux I__2155 (
            .O(N__10233),
            .I(N__10226));
    Span4Mux_v I__2154 (
            .O(N__10230),
            .I(N__10223));
    CEMux I__2153 (
            .O(N__10229),
            .I(N__10220));
    LocalMux I__2152 (
            .O(N__10226),
            .I(N__10217));
    Span4Mux_h I__2151 (
            .O(N__10223),
            .I(N__10212));
    LocalMux I__2150 (
            .O(N__10220),
            .I(N__10212));
    Span12Mux_h I__2149 (
            .O(N__10217),
            .I(N__10208));
    Span4Mux_v I__2148 (
            .O(N__10212),
            .I(N__10205));
    CEMux I__2147 (
            .O(N__10211),
            .I(N__10202));
    Odrv12 I__2146 (
            .O(N__10208),
            .I(\DUT.fifo_tx_inst.N_39 ));
    Odrv4 I__2145 (
            .O(N__10205),
            .I(\DUT.fifo_tx_inst.N_39 ));
    LocalMux I__2144 (
            .O(N__10202),
            .I(\DUT.fifo_tx_inst.N_39 ));
    InMux I__2143 (
            .O(N__10195),
            .I(N__10192));
    LocalMux I__2142 (
            .O(N__10192),
            .I(N__10189));
    Span4Mux_v I__2141 (
            .O(N__10189),
            .I(N__10186));
    Odrv4 I__2140 (
            .O(N__10186),
            .I(\fifo_inst.ftdi_output_inst.rTxE_nZ0Z_1 ));
    InMux I__2139 (
            .O(N__10183),
            .I(N__10180));
    LocalMux I__2138 (
            .O(N__10180),
            .I(N__10177));
    Span4Mux_v I__2137 (
            .O(N__10177),
            .I(N__10174));
    Odrv4 I__2136 (
            .O(N__10174),
            .I(iTxE_n_c));
    InMux I__2135 (
            .O(N__10171),
            .I(N__10168));
    LocalMux I__2134 (
            .O(N__10168),
            .I(N__10164));
    InMux I__2133 (
            .O(N__10167),
            .I(N__10161));
    Span4Mux_v I__2132 (
            .O(N__10164),
            .I(N__10158));
    LocalMux I__2131 (
            .O(N__10161),
            .I(\fifo_inst.ftdi_output_inst.rTxE_nZ0Z_0 ));
    Odrv4 I__2130 (
            .O(N__10158),
            .I(\fifo_inst.ftdi_output_inst.rTxE_nZ0Z_0 ));
    InMux I__2129 (
            .O(N__10153),
            .I(N__10148));
    InMux I__2128 (
            .O(N__10152),
            .I(N__10145));
    InMux I__2127 (
            .O(N__10151),
            .I(N__10142));
    LocalMux I__2126 (
            .O(N__10148),
            .I(N__10139));
    LocalMux I__2125 (
            .O(N__10145),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_1 ));
    LocalMux I__2124 (
            .O(N__10142),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_1 ));
    Odrv4 I__2123 (
            .O(N__10139),
            .I(\DUT.uart_inst0.rx_clk_dividerZ0Z_1 ));
    InMux I__2122 (
            .O(N__10132),
            .I(N__10129));
    LocalMux I__2121 (
            .O(N__10129),
            .I(N__10126));
    Span4Mux_h I__2120 (
            .O(N__10126),
            .I(N__10123));
    Odrv4 I__2119 (
            .O(N__10123),
            .I(\DUT.rFifoDatarx_6 ));
    CascadeMux I__2118 (
            .O(N__10120),
            .I(N__10117));
    InMux I__2117 (
            .O(N__10117),
            .I(N__10113));
    CascadeMux I__2116 (
            .O(N__10116),
            .I(N__10110));
    LocalMux I__2115 (
            .O(N__10113),
            .I(N__10107));
    InMux I__2114 (
            .O(N__10110),
            .I(N__10104));
    Span4Mux_h I__2113 (
            .O(N__10107),
            .I(N__10101));
    LocalMux I__2112 (
            .O(N__10104),
            .I(\DUT.uart_inst0.tx_dataZ0Z_7 ));
    Odrv4 I__2111 (
            .O(N__10101),
            .I(\DUT.uart_inst0.tx_dataZ0Z_7 ));
    CascadeMux I__2110 (
            .O(N__10096),
            .I(\DUT.uart_inst0.tx_data_RNO_0Z0Z_6_cascade_ ));
    InMux I__2109 (
            .O(N__10093),
            .I(N__10090));
    LocalMux I__2108 (
            .O(N__10090),
            .I(N__10086));
    InMux I__2107 (
            .O(N__10089),
            .I(N__10083));
    Span4Mux_h I__2106 (
            .O(N__10086),
            .I(N__10080));
    LocalMux I__2105 (
            .O(N__10083),
            .I(\DUT.uart_inst0.tx_dataZ0Z_6 ));
    Odrv4 I__2104 (
            .O(N__10080),
            .I(\DUT.uart_inst0.tx_dataZ0Z_6 ));
    CascadeMux I__2103 (
            .O(N__10075),
            .I(N__10071));
    CascadeMux I__2102 (
            .O(N__10074),
            .I(N__10068));
    InMux I__2101 (
            .O(N__10071),
            .I(N__10065));
    InMux I__2100 (
            .O(N__10068),
            .I(N__10062));
    LocalMux I__2099 (
            .O(N__10065),
            .I(N__10057));
    LocalMux I__2098 (
            .O(N__10062),
            .I(N__10057));
    Odrv4 I__2097 (
            .O(N__10057),
            .I(\DUT.uart_inst0.tx_dataZ0Z_4 ));
    InMux I__2096 (
            .O(N__10054),
            .I(N__10049));
    InMux I__2095 (
            .O(N__10053),
            .I(N__10044));
    InMux I__2094 (
            .O(N__10052),
            .I(N__10044));
    LocalMux I__2093 (
            .O(N__10049),
            .I(N__10036));
    LocalMux I__2092 (
            .O(N__10044),
            .I(N__10036));
    InMux I__2091 (
            .O(N__10043),
            .I(N__10031));
    InMux I__2090 (
            .O(N__10042),
            .I(N__10031));
    InMux I__2089 (
            .O(N__10041),
            .I(N__10027));
    Span4Mux_v I__2088 (
            .O(N__10036),
            .I(N__10023));
    LocalMux I__2087 (
            .O(N__10031),
            .I(N__10020));
    InMux I__2086 (
            .O(N__10030),
            .I(N__10017));
    LocalMux I__2085 (
            .O(N__10027),
            .I(N__10014));
    InMux I__2084 (
            .O(N__10026),
            .I(N__10011));
    Odrv4 I__2083 (
            .O(N__10023),
            .I(\DUT.rFifoDataror_0 ));
    Odrv4 I__2082 (
            .O(N__10020),
            .I(\DUT.rFifoDataror_0 ));
    LocalMux I__2081 (
            .O(N__10017),
            .I(\DUT.rFifoDataror_0 ));
    Odrv4 I__2080 (
            .O(N__10014),
            .I(\DUT.rFifoDataror_0 ));
    LocalMux I__2079 (
            .O(N__10011),
            .I(\DUT.rFifoDataror_0 ));
    CascadeMux I__2078 (
            .O(N__10000),
            .I(\DUT.uart_inst0.tx_data_RNO_0Z0Z_3_cascade_ ));
    CEMux I__2077 (
            .O(N__9997),
            .I(N__9994));
    LocalMux I__2076 (
            .O(N__9994),
            .I(N__9979));
    InMux I__2075 (
            .O(N__9993),
            .I(N__9976));
    InMux I__2074 (
            .O(N__9992),
            .I(N__9969));
    InMux I__2073 (
            .O(N__9991),
            .I(N__9969));
    InMux I__2072 (
            .O(N__9990),
            .I(N__9969));
    InMux I__2071 (
            .O(N__9989),
            .I(N__9961));
    InMux I__2070 (
            .O(N__9988),
            .I(N__9956));
    InMux I__2069 (
            .O(N__9987),
            .I(N__9956));
    InMux I__2068 (
            .O(N__9986),
            .I(N__9953));
    InMux I__2067 (
            .O(N__9985),
            .I(N__9944));
    InMux I__2066 (
            .O(N__9984),
            .I(N__9944));
    InMux I__2065 (
            .O(N__9983),
            .I(N__9944));
    InMux I__2064 (
            .O(N__9982),
            .I(N__9944));
    Span4Mux_v I__2063 (
            .O(N__9979),
            .I(N__9937));
    LocalMux I__2062 (
            .O(N__9976),
            .I(N__9937));
    LocalMux I__2061 (
            .O(N__9969),
            .I(N__9937));
    InMux I__2060 (
            .O(N__9968),
            .I(N__9932));
    InMux I__2059 (
            .O(N__9967),
            .I(N__9932));
    InMux I__2058 (
            .O(N__9966),
            .I(N__9925));
    InMux I__2057 (
            .O(N__9965),
            .I(N__9925));
    InMux I__2056 (
            .O(N__9964),
            .I(N__9925));
    LocalMux I__2055 (
            .O(N__9961),
            .I(\DUT.uart_inst0.N_152_0 ));
    LocalMux I__2054 (
            .O(N__9956),
            .I(\DUT.uart_inst0.N_152_0 ));
    LocalMux I__2053 (
            .O(N__9953),
            .I(\DUT.uart_inst0.N_152_0 ));
    LocalMux I__2052 (
            .O(N__9944),
            .I(\DUT.uart_inst0.N_152_0 ));
    Odrv4 I__2051 (
            .O(N__9937),
            .I(\DUT.uart_inst0.N_152_0 ));
    LocalMux I__2050 (
            .O(N__9932),
            .I(\DUT.uart_inst0.N_152_0 ));
    LocalMux I__2049 (
            .O(N__9925),
            .I(\DUT.uart_inst0.N_152_0 ));
    InMux I__2048 (
            .O(N__9910),
            .I(N__9907));
    LocalMux I__2047 (
            .O(N__9907),
            .I(N__9904));
    Span4Mux_v I__2046 (
            .O(N__9904),
            .I(N__9900));
    InMux I__2045 (
            .O(N__9903),
            .I(N__9897));
    Span4Mux_h I__2044 (
            .O(N__9900),
            .I(N__9894));
    LocalMux I__2043 (
            .O(N__9897),
            .I(\DUT.uart_inst0.tx_dataZ0Z_3 ));
    Odrv4 I__2042 (
            .O(N__9894),
            .I(\DUT.uart_inst0.tx_dataZ0Z_3 ));
    InMux I__2041 (
            .O(N__9889),
            .I(N__9886));
    LocalMux I__2040 (
            .O(N__9886),
            .I(N__9882));
    InMux I__2039 (
            .O(N__9885),
            .I(N__9879));
    Odrv4 I__2038 (
            .O(N__9882),
            .I(\DUT.uart_inst0.N_159 ));
    LocalMux I__2037 (
            .O(N__9879),
            .I(\DUT.uart_inst0.N_159 ));
    CascadeMux I__2036 (
            .O(N__9874),
            .I(N__9871));
    InMux I__2035 (
            .O(N__9871),
            .I(N__9867));
    InMux I__2034 (
            .O(N__9870),
            .I(N__9864));
    LocalMux I__2033 (
            .O(N__9867),
            .I(N__9861));
    LocalMux I__2032 (
            .O(N__9864),
            .I(\DUT.uart_inst0.tx_dataZ0Z_0 ));
    Odrv4 I__2031 (
            .O(N__9861),
            .I(\DUT.uart_inst0.tx_dataZ0Z_0 ));
    InMux I__2030 (
            .O(N__9856),
            .I(N__9852));
    InMux I__2029 (
            .O(N__9855),
            .I(N__9846));
    LocalMux I__2028 (
            .O(N__9852),
            .I(N__9843));
    InMux I__2027 (
            .O(N__9851),
            .I(N__9839));
    CascadeMux I__2026 (
            .O(N__9850),
            .I(N__9834));
    InMux I__2025 (
            .O(N__9849),
            .I(N__9828));
    LocalMux I__2024 (
            .O(N__9846),
            .I(N__9825));
    Span4Mux_h I__2023 (
            .O(N__9843),
            .I(N__9822));
    InMux I__2022 (
            .O(N__9842),
            .I(N__9819));
    LocalMux I__2021 (
            .O(N__9839),
            .I(N__9816));
    InMux I__2020 (
            .O(N__9838),
            .I(N__9813));
    InMux I__2019 (
            .O(N__9837),
            .I(N__9804));
    InMux I__2018 (
            .O(N__9834),
            .I(N__9804));
    InMux I__2017 (
            .O(N__9833),
            .I(N__9804));
    InMux I__2016 (
            .O(N__9832),
            .I(N__9804));
    InMux I__2015 (
            .O(N__9831),
            .I(N__9801));
    LocalMux I__2014 (
            .O(N__9828),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_1 ));
    Odrv4 I__2013 (
            .O(N__9825),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_1 ));
    Odrv4 I__2012 (
            .O(N__9822),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_1 ));
    LocalMux I__2011 (
            .O(N__9819),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_1 ));
    Odrv12 I__2010 (
            .O(N__9816),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_1 ));
    LocalMux I__2009 (
            .O(N__9813),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_1 ));
    LocalMux I__2008 (
            .O(N__9804),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_1 ));
    LocalMux I__2007 (
            .O(N__9801),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_1 ));
    InMux I__2006 (
            .O(N__9784),
            .I(N__9781));
    LocalMux I__2005 (
            .O(N__9781),
            .I(N__9778));
    Span4Mux_h I__2004 (
            .O(N__9778),
            .I(N__9775));
    Odrv4 I__2003 (
            .O(N__9775),
            .I(\DUT.uart_inst0.g0_i_a4_0_4 ));
    InMux I__2002 (
            .O(N__9772),
            .I(N__9768));
    InMux I__2001 (
            .O(N__9771),
            .I(N__9760));
    LocalMux I__2000 (
            .O(N__9768),
            .I(N__9756));
    InMux I__1999 (
            .O(N__9767),
            .I(N__9748));
    InMux I__1998 (
            .O(N__9766),
            .I(N__9748));
    CascadeMux I__1997 (
            .O(N__9765),
            .I(N__9745));
    CascadeMux I__1996 (
            .O(N__9764),
            .I(N__9742));
    InMux I__1995 (
            .O(N__9763),
            .I(N__9737));
    LocalMux I__1994 (
            .O(N__9760),
            .I(N__9734));
    InMux I__1993 (
            .O(N__9759),
            .I(N__9731));
    Span4Mux_v I__1992 (
            .O(N__9756),
            .I(N__9728));
    InMux I__1991 (
            .O(N__9755),
            .I(N__9725));
    InMux I__1990 (
            .O(N__9754),
            .I(N__9720));
    InMux I__1989 (
            .O(N__9753),
            .I(N__9720));
    LocalMux I__1988 (
            .O(N__9748),
            .I(N__9717));
    InMux I__1987 (
            .O(N__9745),
            .I(N__9708));
    InMux I__1986 (
            .O(N__9742),
            .I(N__9708));
    InMux I__1985 (
            .O(N__9741),
            .I(N__9708));
    InMux I__1984 (
            .O(N__9740),
            .I(N__9708));
    LocalMux I__1983 (
            .O(N__9737),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_0 ));
    Odrv4 I__1982 (
            .O(N__9734),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_0 ));
    LocalMux I__1981 (
            .O(N__9731),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_0 ));
    Odrv4 I__1980 (
            .O(N__9728),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_0 ));
    LocalMux I__1979 (
            .O(N__9725),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_0 ));
    LocalMux I__1978 (
            .O(N__9720),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_0 ));
    Odrv12 I__1977 (
            .O(N__9717),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_0 ));
    LocalMux I__1976 (
            .O(N__9708),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_0 ));
    CascadeMux I__1975 (
            .O(N__9691),
            .I(\DUT.uart_inst0.g0_i_a4_0_5_cascade_ ));
    InMux I__1974 (
            .O(N__9688),
            .I(N__9685));
    LocalMux I__1973 (
            .O(N__9685),
            .I(\DUT.uart_inst0.N_15 ));
    InMux I__1972 (
            .O(N__9682),
            .I(N__9679));
    LocalMux I__1971 (
            .O(N__9679),
            .I(\DUT.uart_inst0.N_7 ));
    InMux I__1970 (
            .O(N__9676),
            .I(N__9667));
    InMux I__1969 (
            .O(N__9675),
            .I(N__9664));
    CascadeMux I__1968 (
            .O(N__9674),
            .I(N__9661));
    CascadeMux I__1967 (
            .O(N__9673),
            .I(N__9653));
    CascadeMux I__1966 (
            .O(N__9672),
            .I(N__9644));
    CascadeMux I__1965 (
            .O(N__9671),
            .I(N__9639));
    CascadeMux I__1964 (
            .O(N__9670),
            .I(N__9636));
    LocalMux I__1963 (
            .O(N__9667),
            .I(N__9631));
    LocalMux I__1962 (
            .O(N__9664),
            .I(N__9631));
    InMux I__1961 (
            .O(N__9661),
            .I(N__9628));
    InMux I__1960 (
            .O(N__9660),
            .I(N__9621));
    InMux I__1959 (
            .O(N__9659),
            .I(N__9621));
    InMux I__1958 (
            .O(N__9658),
            .I(N__9621));
    InMux I__1957 (
            .O(N__9657),
            .I(N__9612));
    InMux I__1956 (
            .O(N__9656),
            .I(N__9612));
    InMux I__1955 (
            .O(N__9653),
            .I(N__9612));
    InMux I__1954 (
            .O(N__9652),
            .I(N__9612));
    InMux I__1953 (
            .O(N__9651),
            .I(N__9599));
    InMux I__1952 (
            .O(N__9650),
            .I(N__9599));
    InMux I__1951 (
            .O(N__9649),
            .I(N__9599));
    InMux I__1950 (
            .O(N__9648),
            .I(N__9599));
    InMux I__1949 (
            .O(N__9647),
            .I(N__9599));
    InMux I__1948 (
            .O(N__9644),
            .I(N__9599));
    InMux I__1947 (
            .O(N__9643),
            .I(N__9590));
    InMux I__1946 (
            .O(N__9642),
            .I(N__9590));
    InMux I__1945 (
            .O(N__9639),
            .I(N__9590));
    InMux I__1944 (
            .O(N__9636),
            .I(N__9590));
    Odrv4 I__1943 (
            .O(N__9631),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__1942 (
            .O(N__9628),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__1941 (
            .O(N__9621),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__1940 (
            .O(N__9612),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__1939 (
            .O(N__9599),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__1938 (
            .O(N__9590),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ));
    CascadeMux I__1937 (
            .O(N__9577),
            .I(N__9574));
    InMux I__1936 (
            .O(N__9574),
            .I(N__9571));
    LocalMux I__1935 (
            .O(N__9571),
            .I(N__9568));
    Span4Mux_h I__1934 (
            .O(N__9568),
            .I(N__9565));
    Odrv4 I__1933 (
            .O(N__9565),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_3 ));
    InMux I__1932 (
            .O(N__9562),
            .I(N__9559));
    LocalMux I__1931 (
            .O(N__9559),
            .I(N__9556));
    Odrv4 I__1930 (
            .O(N__9556),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3 ));
    InMux I__1929 (
            .O(N__9553),
            .I(N__9550));
    LocalMux I__1928 (
            .O(N__9550),
            .I(\DUT.rFifoDatarx_3 ));
    InMux I__1927 (
            .O(N__9547),
            .I(N__9544));
    LocalMux I__1926 (
            .O(N__9544),
            .I(\DUT.uart_inst0.tx_bits_remaining_RNO_1Z0Z_2 ));
    InMux I__1925 (
            .O(N__9541),
            .I(N__9538));
    LocalMux I__1924 (
            .O(N__9538),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_9 ));
    InMux I__1923 (
            .O(N__9535),
            .I(N__9532));
    LocalMux I__1922 (
            .O(N__9532),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_8 ));
    InMux I__1921 (
            .O(N__9529),
            .I(N__9526));
    LocalMux I__1920 (
            .O(N__9526),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_7 ));
    CascadeMux I__1919 (
            .O(N__9523),
            .I(N__9518));
    InMux I__1918 (
            .O(N__9522),
            .I(N__9514));
    CascadeMux I__1917 (
            .O(N__9521),
            .I(N__9510));
    InMux I__1916 (
            .O(N__9518),
            .I(N__9506));
    CascadeMux I__1915 (
            .O(N__9517),
            .I(N__9500));
    LocalMux I__1914 (
            .O(N__9514),
            .I(N__9497));
    InMux I__1913 (
            .O(N__9513),
            .I(N__9490));
    InMux I__1912 (
            .O(N__9510),
            .I(N__9490));
    InMux I__1911 (
            .O(N__9509),
            .I(N__9490));
    LocalMux I__1910 (
            .O(N__9506),
            .I(N__9487));
    InMux I__1909 (
            .O(N__9505),
            .I(N__9484));
    InMux I__1908 (
            .O(N__9504),
            .I(N__9481));
    InMux I__1907 (
            .O(N__9503),
            .I(N__9476));
    InMux I__1906 (
            .O(N__9500),
            .I(N__9476));
    Odrv4 I__1905 (
            .O(N__9497),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_3 ));
    LocalMux I__1904 (
            .O(N__9490),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_3 ));
    Odrv12 I__1903 (
            .O(N__9487),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_3 ));
    LocalMux I__1902 (
            .O(N__9484),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_3 ));
    LocalMux I__1901 (
            .O(N__9481),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_3 ));
    LocalMux I__1900 (
            .O(N__9476),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_3 ));
    CascadeMux I__1899 (
            .O(N__9463),
            .I(N__9458));
    CascadeMux I__1898 (
            .O(N__9462),
            .I(N__9453));
    InMux I__1897 (
            .O(N__9461),
            .I(N__9446));
    InMux I__1896 (
            .O(N__9458),
            .I(N__9446));
    CascadeMux I__1895 (
            .O(N__9457),
            .I(N__9443));
    CascadeMux I__1894 (
            .O(N__9456),
            .I(N__9440));
    InMux I__1893 (
            .O(N__9453),
            .I(N__9437));
    InMux I__1892 (
            .O(N__9452),
            .I(N__9434));
    InMux I__1891 (
            .O(N__9451),
            .I(N__9431));
    LocalMux I__1890 (
            .O(N__9446),
            .I(N__9428));
    InMux I__1889 (
            .O(N__9443),
            .I(N__9425));
    InMux I__1888 (
            .O(N__9440),
            .I(N__9422));
    LocalMux I__1887 (
            .O(N__9437),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_5 ));
    LocalMux I__1886 (
            .O(N__9434),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_5 ));
    LocalMux I__1885 (
            .O(N__9431),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_5 ));
    Odrv4 I__1884 (
            .O(N__9428),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_5 ));
    LocalMux I__1883 (
            .O(N__9425),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_5 ));
    LocalMux I__1882 (
            .O(N__9422),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_5 ));
    InMux I__1881 (
            .O(N__9409),
            .I(N__9406));
    LocalMux I__1880 (
            .O(N__9406),
            .I(N__9396));
    InMux I__1879 (
            .O(N__9405),
            .I(N__9387));
    InMux I__1878 (
            .O(N__9404),
            .I(N__9387));
    InMux I__1877 (
            .O(N__9403),
            .I(N__9387));
    InMux I__1876 (
            .O(N__9402),
            .I(N__9387));
    InMux I__1875 (
            .O(N__9401),
            .I(N__9382));
    InMux I__1874 (
            .O(N__9400),
            .I(N__9379));
    InMux I__1873 (
            .O(N__9399),
            .I(N__9376));
    Span4Mux_h I__1872 (
            .O(N__9396),
            .I(N__9373));
    LocalMux I__1871 (
            .O(N__9387),
            .I(N__9370));
    InMux I__1870 (
            .O(N__9386),
            .I(N__9365));
    InMux I__1869 (
            .O(N__9385),
            .I(N__9365));
    LocalMux I__1868 (
            .O(N__9382),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_2 ));
    LocalMux I__1867 (
            .O(N__9379),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_2 ));
    LocalMux I__1866 (
            .O(N__9376),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_2 ));
    Odrv4 I__1865 (
            .O(N__9373),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_2 ));
    Odrv4 I__1864 (
            .O(N__9370),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_2 ));
    LocalMux I__1863 (
            .O(N__9365),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_2 ));
    CascadeMux I__1862 (
            .O(N__9352),
            .I(\DUT.uart_inst0.tx_data_i_m_4_0_cascade_ ));
    InMux I__1861 (
            .O(N__9349),
            .I(N__9344));
    InMux I__1860 (
            .O(N__9348),
            .I(N__9340));
    InMux I__1859 (
            .O(N__9347),
            .I(N__9336));
    LocalMux I__1858 (
            .O(N__9344),
            .I(N__9330));
    InMux I__1857 (
            .O(N__9343),
            .I(N__9327));
    LocalMux I__1856 (
            .O(N__9340),
            .I(N__9324));
    InMux I__1855 (
            .O(N__9339),
            .I(N__9321));
    LocalMux I__1854 (
            .O(N__9336),
            .I(N__9318));
    InMux I__1853 (
            .O(N__9335),
            .I(N__9311));
    InMux I__1852 (
            .O(N__9334),
            .I(N__9311));
    InMux I__1851 (
            .O(N__9333),
            .I(N__9311));
    Span4Mux_h I__1850 (
            .O(N__9330),
            .I(N__9308));
    LocalMux I__1849 (
            .O(N__9327),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_4 ));
    Odrv4 I__1848 (
            .O(N__9324),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_4 ));
    LocalMux I__1847 (
            .O(N__9321),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_4 ));
    Odrv4 I__1846 (
            .O(N__9318),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_4 ));
    LocalMux I__1845 (
            .O(N__9311),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_4 ));
    Odrv4 I__1844 (
            .O(N__9308),
            .I(\DUT.uart_inst0.tx_countdownZ0Z_4 ));
    CascadeMux I__1843 (
            .O(N__9295),
            .I(N__9292));
    InMux I__1842 (
            .O(N__9292),
            .I(N__9288));
    InMux I__1841 (
            .O(N__9291),
            .I(N__9285));
    LocalMux I__1840 (
            .O(N__9288),
            .I(N__9282));
    LocalMux I__1839 (
            .O(N__9285),
            .I(\DUT.uart_inst0.tx_countdown_0_c4_i ));
    Odrv4 I__1838 (
            .O(N__9282),
            .I(\DUT.uart_inst0.tx_countdown_0_c4_i ));
    InMux I__1837 (
            .O(N__9277),
            .I(N__9274));
    LocalMux I__1836 (
            .O(N__9274),
            .I(\DUT.uart_inst0.tx_state_ns_0_o3_1_0_1 ));
    InMux I__1835 (
            .O(N__9271),
            .I(N__9268));
    LocalMux I__1834 (
            .O(N__9268),
            .I(N__9265));
    Span4Mux_v I__1833 (
            .O(N__9265),
            .I(N__9261));
    InMux I__1832 (
            .O(N__9264),
            .I(N__9258));
    Odrv4 I__1831 (
            .O(N__9261),
            .I(G_148));
    LocalMux I__1830 (
            .O(N__9258),
            .I(G_148));
    CascadeMux I__1829 (
            .O(N__9253),
            .I(\fifo_inst.ftdi_output_inst.N_95_cascade_ ));
    InMux I__1828 (
            .O(N__9250),
            .I(N__9246));
    InMux I__1827 (
            .O(N__9249),
            .I(N__9243));
    LocalMux I__1826 (
            .O(N__9246),
            .I(N__9240));
    LocalMux I__1825 (
            .O(N__9243),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_3 ));
    Odrv4 I__1824 (
            .O(N__9240),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_3 ));
    InMux I__1823 (
            .O(N__9235),
            .I(N__9232));
    LocalMux I__1822 (
            .O(N__9232),
            .I(N__9229));
    Span4Mux_h I__1821 (
            .O(N__9229),
            .I(N__9225));
    InMux I__1820 (
            .O(N__9228),
            .I(N__9222));
    Odrv4 I__1819 (
            .O(N__9225),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2 ));
    LocalMux I__1818 (
            .O(N__9222),
            .I(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2 ));
    InMux I__1817 (
            .O(N__9217),
            .I(N__9214));
    LocalMux I__1816 (
            .O(N__9214),
            .I(\fifo_inst.ftdi_output_inst.N_95 ));
    CascadeMux I__1815 (
            .O(N__9211),
            .I(\fifo_inst.ftdi_output_inst.m14_1_cascade_ ));
    InMux I__1814 (
            .O(N__9208),
            .I(N__9202));
    InMux I__1813 (
            .O(N__9207),
            .I(N__9202));
    LocalMux I__1812 (
            .O(N__9202),
            .I(\fifo_inst.ftdi_output_inst.N_86_0 ));
    CascadeMux I__1811 (
            .O(N__9199),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_9_cascade_ ));
    InMux I__1810 (
            .O(N__9196),
            .I(N__9193));
    LocalMux I__1809 (
            .O(N__9193),
            .I(N__9189));
    InMux I__1808 (
            .O(N__9192),
            .I(N__9186));
    Odrv4 I__1807 (
            .O(N__9189),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_13 ));
    LocalMux I__1806 (
            .O(N__9186),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_13 ));
    InMux I__1805 (
            .O(N__9181),
            .I(N__9177));
    InMux I__1804 (
            .O(N__9180),
            .I(N__9174));
    LocalMux I__1803 (
            .O(N__9177),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_5 ));
    LocalMux I__1802 (
            .O(N__9174),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_5 ));
    CascadeMux I__1801 (
            .O(N__9169),
            .I(N__9166));
    InMux I__1800 (
            .O(N__9166),
            .I(N__9162));
    InMux I__1799 (
            .O(N__9165),
            .I(N__9158));
    LocalMux I__1798 (
            .O(N__9162),
            .I(N__9155));
    InMux I__1797 (
            .O(N__9161),
            .I(N__9152));
    LocalMux I__1796 (
            .O(N__9158),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_5 ));
    Odrv4 I__1795 (
            .O(N__9155),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_5 ));
    LocalMux I__1794 (
            .O(N__9152),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_5 ));
    InMux I__1793 (
            .O(N__9145),
            .I(N__9137));
    InMux I__1792 (
            .O(N__9144),
            .I(N__9137));
    InMux I__1791 (
            .O(N__9143),
            .I(N__9132));
    InMux I__1790 (
            .O(N__9142),
            .I(N__9132));
    LocalMux I__1789 (
            .O(N__9137),
            .I(N__9124));
    LocalMux I__1788 (
            .O(N__9132),
            .I(N__9121));
    InMux I__1787 (
            .O(N__9131),
            .I(N__9116));
    InMux I__1786 (
            .O(N__9130),
            .I(N__9116));
    InMux I__1785 (
            .O(N__9129),
            .I(N__9111));
    InMux I__1784 (
            .O(N__9128),
            .I(N__9111));
    InMux I__1783 (
            .O(N__9127),
            .I(N__9108));
    Odrv4 I__1782 (
            .O(N__9124),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    Odrv4 I__1781 (
            .O(N__9121),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    LocalMux I__1780 (
            .O(N__9116),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    LocalMux I__1779 (
            .O(N__9111),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    LocalMux I__1778 (
            .O(N__9108),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0 ));
    CascadeMux I__1777 (
            .O(N__9097),
            .I(N__9094));
    InMux I__1776 (
            .O(N__9094),
            .I(N__9087));
    InMux I__1775 (
            .O(N__9093),
            .I(N__9087));
    InMux I__1774 (
            .O(N__9092),
            .I(N__9084));
    LocalMux I__1773 (
            .O(N__9087),
            .I(N__9081));
    LocalMux I__1772 (
            .O(N__9084),
            .I(N__9078));
    Span4Mux_h I__1771 (
            .O(N__9081),
            .I(N__9075));
    Odrv4 I__1770 (
            .O(N__9078),
            .I(\DUT.uart_inst0.N_70 ));
    Odrv4 I__1769 (
            .O(N__9075),
            .I(\DUT.uart_inst0.N_70 ));
    InMux I__1768 (
            .O(N__9070),
            .I(N__9063));
    InMux I__1767 (
            .O(N__9069),
            .I(N__9063));
    InMux I__1766 (
            .O(N__9068),
            .I(N__9059));
    LocalMux I__1765 (
            .O(N__9063),
            .I(N__9056));
    InMux I__1764 (
            .O(N__9062),
            .I(N__9053));
    LocalMux I__1763 (
            .O(N__9059),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    Odrv12 I__1762 (
            .O(N__9056),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    LocalMux I__1761 (
            .O(N__9053),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_3 ));
    InMux I__1760 (
            .O(N__9046),
            .I(N__9042));
    InMux I__1759 (
            .O(N__9045),
            .I(N__9039));
    LocalMux I__1758 (
            .O(N__9042),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_11 ));
    LocalMux I__1757 (
            .O(N__9039),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_11 ));
    CascadeMux I__1756 (
            .O(N__9034),
            .I(N__9031));
    InMux I__1755 (
            .O(N__9031),
            .I(N__9027));
    InMux I__1754 (
            .O(N__9030),
            .I(N__9024));
    LocalMux I__1753 (
            .O(N__9027),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_12 ));
    LocalMux I__1752 (
            .O(N__9024),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_12 ));
    InMux I__1751 (
            .O(N__9019),
            .I(N__9016));
    LocalMux I__1750 (
            .O(N__9016),
            .I(N__9013));
    Odrv4 I__1749 (
            .O(N__9013),
            .I(\DUT.rFifoDatarx_5 ));
    CascadeMux I__1748 (
            .O(N__9010),
            .I(\DUT.uart_inst0.tx_data_RNO_0Z0Z_5_cascade_ ));
    InMux I__1747 (
            .O(N__9007),
            .I(N__9003));
    InMux I__1746 (
            .O(N__9006),
            .I(N__9000));
    LocalMux I__1745 (
            .O(N__9003),
            .I(N__8997));
    LocalMux I__1744 (
            .O(N__9000),
            .I(\DUT.uart_inst0.tx_dataZ0Z_5 ));
    Odrv4 I__1743 (
            .O(N__8997),
            .I(\DUT.uart_inst0.tx_dataZ0Z_5 ));
    InMux I__1742 (
            .O(N__8992),
            .I(N__8988));
    InMux I__1741 (
            .O(N__8991),
            .I(N__8985));
    LocalMux I__1740 (
            .O(N__8988),
            .I(N__8978));
    LocalMux I__1739 (
            .O(N__8985),
            .I(N__8978));
    InMux I__1738 (
            .O(N__8984),
            .I(N__8975));
    InMux I__1737 (
            .O(N__8983),
            .I(N__8972));
    Span4Mux_h I__1736 (
            .O(N__8978),
            .I(N__8967));
    LocalMux I__1735 (
            .O(N__8975),
            .I(N__8967));
    LocalMux I__1734 (
            .O(N__8972),
            .I(N__8964));
    Span4Mux_v I__1733 (
            .O(N__8967),
            .I(N__8961));
    Span4Mux_h I__1732 (
            .O(N__8964),
            .I(N__8958));
    Span4Mux_v I__1731 (
            .O(N__8961),
            .I(N__8955));
    Span4Mux_v I__1730 (
            .O(N__8958),
            .I(N__8952));
    Odrv4 I__1729 (
            .O(N__8955),
            .I(rTxByteZ0Z_1));
    Odrv4 I__1728 (
            .O(N__8952),
            .I(rTxByteZ0Z_1));
    InMux I__1727 (
            .O(N__8947),
            .I(N__8944));
    LocalMux I__1726 (
            .O(N__8944),
            .I(N__8941));
    Odrv4 I__1725 (
            .O(N__8941),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_1 ));
    InMux I__1724 (
            .O(N__8938),
            .I(N__8934));
    InMux I__1723 (
            .O(N__8937),
            .I(N__8930));
    LocalMux I__1722 (
            .O(N__8934),
            .I(N__8926));
    InMux I__1721 (
            .O(N__8933),
            .I(N__8923));
    LocalMux I__1720 (
            .O(N__8930),
            .I(N__8920));
    InMux I__1719 (
            .O(N__8929),
            .I(N__8917));
    Span4Mux_v I__1718 (
            .O(N__8926),
            .I(N__8914));
    LocalMux I__1717 (
            .O(N__8923),
            .I(N__8911));
    Span4Mux_v I__1716 (
            .O(N__8920),
            .I(N__8906));
    LocalMux I__1715 (
            .O(N__8917),
            .I(N__8906));
    Span4Mux_v I__1714 (
            .O(N__8914),
            .I(N__8903));
    Span12Mux_v I__1713 (
            .O(N__8911),
            .I(N__8900));
    Span4Mux_v I__1712 (
            .O(N__8906),
            .I(N__8897));
    Odrv4 I__1711 (
            .O(N__8903),
            .I(rTxByteZ0Z_0));
    Odrv12 I__1710 (
            .O(N__8900),
            .I(rTxByteZ0Z_0));
    Odrv4 I__1709 (
            .O(N__8897),
            .I(rTxByteZ0Z_0));
    InMux I__1708 (
            .O(N__8890),
            .I(N__8887));
    LocalMux I__1707 (
            .O(N__8887),
            .I(N__8884));
    Span4Mux_v I__1706 (
            .O(N__8884),
            .I(N__8881));
    Odrv4 I__1705 (
            .O(N__8881),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_0 ));
    InMux I__1704 (
            .O(N__8878),
            .I(N__8873));
    InMux I__1703 (
            .O(N__8877),
            .I(N__8870));
    InMux I__1702 (
            .O(N__8876),
            .I(N__8867));
    LocalMux I__1701 (
            .O(N__8873),
            .I(N__8863));
    LocalMux I__1700 (
            .O(N__8870),
            .I(N__8858));
    LocalMux I__1699 (
            .O(N__8867),
            .I(N__8858));
    InMux I__1698 (
            .O(N__8866),
            .I(N__8855));
    Span4Mux_v I__1697 (
            .O(N__8863),
            .I(N__8852));
    Span4Mux_h I__1696 (
            .O(N__8858),
            .I(N__8847));
    LocalMux I__1695 (
            .O(N__8855),
            .I(N__8847));
    Span4Mux_v I__1694 (
            .O(N__8852),
            .I(N__8844));
    Span4Mux_v I__1693 (
            .O(N__8847),
            .I(N__8841));
    Odrv4 I__1692 (
            .O(N__8844),
            .I(rTxByteZ0Z_6));
    Odrv4 I__1691 (
            .O(N__8841),
            .I(rTxByteZ0Z_6));
    InMux I__1690 (
            .O(N__8836),
            .I(N__8833));
    LocalMux I__1689 (
            .O(N__8833),
            .I(N__8830));
    Odrv4 I__1688 (
            .O(N__8830),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_6 ));
    InMux I__1687 (
            .O(N__8827),
            .I(N__8824));
    LocalMux I__1686 (
            .O(N__8824),
            .I(\DUT.uart_inst0.tx_data_8_321_a2_0 ));
    CascadeMux I__1685 (
            .O(N__8821),
            .I(\DUT.uart_inst0.tx_countdown_0_1_5_cascade_ ));
    InMux I__1684 (
            .O(N__8818),
            .I(N__8815));
    LocalMux I__1683 (
            .O(N__8815),
            .I(\DUT.uart_inst0.g0_i_o4_0_5 ));
    CascadeMux I__1682 (
            .O(N__8812),
            .I(\DUT.uart_inst0.N_14_cascade_ ));
    IoInMux I__1681 (
            .O(N__8809),
            .I(N__8806));
    LocalMux I__1680 (
            .O(N__8806),
            .I(N__8803));
    Span4Mux_s1_v I__1679 (
            .O(N__8803),
            .I(N__8800));
    Sp12to4 I__1678 (
            .O(N__8800),
            .I(N__8797));
    Span12Mux_h I__1677 (
            .O(N__8797),
            .I(N__8793));
    CascadeMux I__1676 (
            .O(N__8796),
            .I(N__8790));
    Span12Mux_v I__1675 (
            .O(N__8793),
            .I(N__8787));
    InMux I__1674 (
            .O(N__8790),
            .I(N__8784));
    Odrv12 I__1673 (
            .O(N__8787),
            .I(P1A7_c));
    LocalMux I__1672 (
            .O(N__8784),
            .I(P1A7_c));
    InMux I__1671 (
            .O(N__8779),
            .I(N__8776));
    LocalMux I__1670 (
            .O(N__8776),
            .I(\DUT.uart_inst0.N_6 ));
    InMux I__1669 (
            .O(N__8773),
            .I(N__8770));
    LocalMux I__1668 (
            .O(N__8770),
            .I(N__8767));
    Odrv4 I__1667 (
            .O(N__8767),
            .I(\DUT.uart_inst0.un1_tx_bits_remaining_axbxc2_N_4L5_1_0 ));
    InMux I__1666 (
            .O(N__8764),
            .I(N__8761));
    LocalMux I__1665 (
            .O(N__8761),
            .I(N__8758));
    Odrv4 I__1664 (
            .O(N__8758),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1 ));
    CascadeMux I__1663 (
            .O(N__8755),
            .I(N__8752));
    InMux I__1662 (
            .O(N__8752),
            .I(N__8749));
    LocalMux I__1661 (
            .O(N__8749),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_1 ));
    CascadeMux I__1660 (
            .O(N__8746),
            .I(N__8743));
    InMux I__1659 (
            .O(N__8743),
            .I(N__8740));
    LocalMux I__1658 (
            .O(N__8740),
            .I(N__8736));
    InMux I__1657 (
            .O(N__8739),
            .I(N__8733));
    Odrv4 I__1656 (
            .O(N__8736),
            .I(\DUT.uart_inst0.tx_dataZ0Z_2 ));
    LocalMux I__1655 (
            .O(N__8733),
            .I(\DUT.uart_inst0.tx_dataZ0Z_2 ));
    CascadeMux I__1654 (
            .O(N__8728),
            .I(\DUT.rFifoDatarx_1_cascade_ ));
    CascadeMux I__1653 (
            .O(N__8725),
            .I(\DUT.uart_inst0.tx_data_RNO_0Z0Z_1_cascade_ ));
    InMux I__1652 (
            .O(N__8722),
            .I(N__8719));
    LocalMux I__1651 (
            .O(N__8719),
            .I(N__8715));
    InMux I__1650 (
            .O(N__8718),
            .I(N__8712));
    Odrv4 I__1649 (
            .O(N__8715),
            .I(\DUT.uart_inst0.tx_dataZ0Z_1 ));
    LocalMux I__1648 (
            .O(N__8712),
            .I(\DUT.uart_inst0.tx_dataZ0Z_1 ));
    InMux I__1647 (
            .O(N__8707),
            .I(N__8704));
    LocalMux I__1646 (
            .O(N__8704),
            .I(\DUT.uart_inst0.tx_data_RNO_0Z0Z_0 ));
    CascadeMux I__1645 (
            .O(N__8701),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_6_cascade_ ));
    InMux I__1644 (
            .O(N__8698),
            .I(N__8695));
    LocalMux I__1643 (
            .O(N__8695),
            .I(\DUT.uart_inst0.un1_tx_bits_remaining_axbxc2_N_4L5_1_1 ));
    CascadeMux I__1642 (
            .O(N__8692),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_0_cascade_ ));
    InMux I__1641 (
            .O(N__8689),
            .I(N__8686));
    LocalMux I__1640 (
            .O(N__8686),
            .I(\DUT.uart_inst0.un1_tx_bits_remaining_axbxc2_N_4L5_1 ));
    InMux I__1639 (
            .O(N__8683),
            .I(N__8677));
    InMux I__1638 (
            .O(N__8682),
            .I(N__8670));
    CascadeMux I__1637 (
            .O(N__8681),
            .I(N__8667));
    CascadeMux I__1636 (
            .O(N__8680),
            .I(N__8664));
    LocalMux I__1635 (
            .O(N__8677),
            .I(N__8661));
    InMux I__1634 (
            .O(N__8676),
            .I(N__8658));
    InMux I__1633 (
            .O(N__8675),
            .I(N__8651));
    InMux I__1632 (
            .O(N__8674),
            .I(N__8651));
    InMux I__1631 (
            .O(N__8673),
            .I(N__8651));
    LocalMux I__1630 (
            .O(N__8670),
            .I(N__8648));
    InMux I__1629 (
            .O(N__8667),
            .I(N__8643));
    InMux I__1628 (
            .O(N__8664),
            .I(N__8643));
    Span4Mux_h I__1627 (
            .O(N__8661),
            .I(N__8636));
    LocalMux I__1626 (
            .O(N__8658),
            .I(N__8636));
    LocalMux I__1625 (
            .O(N__8651),
            .I(N__8636));
    Odrv4 I__1624 (
            .O(N__8648),
            .I(rRxReadZ0));
    LocalMux I__1623 (
            .O(N__8643),
            .I(rRxReadZ0));
    Odrv4 I__1622 (
            .O(N__8636),
            .I(rRxReadZ0));
    CascadeMux I__1621 (
            .O(N__8629),
            .I(N__8626));
    InMux I__1620 (
            .O(N__8626),
            .I(N__8623));
    LocalMux I__1619 (
            .O(N__8623),
            .I(N__8617));
    InMux I__1618 (
            .O(N__8622),
            .I(N__8614));
    InMux I__1617 (
            .O(N__8621),
            .I(N__8609));
    InMux I__1616 (
            .O(N__8620),
            .I(N__8609));
    Odrv4 I__1615 (
            .O(N__8617),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_1 ));
    LocalMux I__1614 (
            .O(N__8614),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_1 ));
    LocalMux I__1613 (
            .O(N__8609),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_1 ));
    CascadeMux I__1612 (
            .O(N__8602),
            .I(N__8599));
    InMux I__1611 (
            .O(N__8599),
            .I(N__8596));
    LocalMux I__1610 (
            .O(N__8596),
            .I(N__8593));
    Odrv4 I__1609 (
            .O(N__8593),
            .I(\DUT.fifo_tx_inst.rFifoCount_RNIBPFMZ0Z_1 ));
    CascadeMux I__1608 (
            .O(N__8590),
            .I(\DUT.uart_inst0.g0_0_0_a3_3_cascade_ ));
    CascadeMux I__1607 (
            .O(N__8587),
            .I(\DUT.uart_inst0.g0_0_0_a3_5_cascade_ ));
    InMux I__1606 (
            .O(N__8584),
            .I(N__8581));
    LocalMux I__1605 (
            .O(N__8581),
            .I(\DUT.uart_inst0.N_159_0_0 ));
    InMux I__1604 (
            .O(N__8578),
            .I(N__8570));
    InMux I__1603 (
            .O(N__8577),
            .I(N__8570));
    InMux I__1602 (
            .O(N__8576),
            .I(N__8565));
    InMux I__1601 (
            .O(N__8575),
            .I(N__8565));
    LocalMux I__1600 (
            .O(N__8570),
            .I(N__8562));
    LocalMux I__1599 (
            .O(N__8565),
            .I(N__8559));
    Odrv12 I__1598 (
            .O(N__8562),
            .I(\DUT.N_37 ));
    Odrv4 I__1597 (
            .O(N__8559),
            .I(\DUT.N_37 ));
    InMux I__1596 (
            .O(N__8554),
            .I(N__8551));
    LocalMux I__1595 (
            .O(N__8551),
            .I(N__8548));
    Odrv4 I__1594 (
            .O(N__8548),
            .I(\DUT.uart_inst0.N_105 ));
    InMux I__1593 (
            .O(N__8545),
            .I(N__8541));
    CascadeMux I__1592 (
            .O(N__8544),
            .I(N__8537));
    LocalMux I__1591 (
            .O(N__8541),
            .I(N__8534));
    InMux I__1590 (
            .O(N__8540),
            .I(N__8531));
    InMux I__1589 (
            .O(N__8537),
            .I(N__8528));
    Odrv4 I__1588 (
            .O(N__8534),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_1 ));
    LocalMux I__1587 (
            .O(N__8531),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_1 ));
    LocalMux I__1586 (
            .O(N__8528),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_1 ));
    InMux I__1585 (
            .O(N__8521),
            .I(N__8518));
    LocalMux I__1584 (
            .O(N__8518),
            .I(N__8515));
    Odrv4 I__1583 (
            .O(N__8515),
            .I(\DUT.uart_inst0.N_102 ));
    CascadeMux I__1582 (
            .O(N__8512),
            .I(N__8509));
    InMux I__1581 (
            .O(N__8509),
            .I(N__8505));
    CascadeMux I__1580 (
            .O(N__8508),
            .I(N__8501));
    LocalMux I__1579 (
            .O(N__8505),
            .I(N__8498));
    InMux I__1578 (
            .O(N__8504),
            .I(N__8495));
    InMux I__1577 (
            .O(N__8501),
            .I(N__8492));
    Odrv4 I__1576 (
            .O(N__8498),
            .I(\DUT.uart_inst0.rx_countdownZ1Z_3 ));
    LocalMux I__1575 (
            .O(N__8495),
            .I(\DUT.uart_inst0.rx_countdownZ1Z_3 ));
    LocalMux I__1574 (
            .O(N__8492),
            .I(\DUT.uart_inst0.rx_countdownZ1Z_3 ));
    InMux I__1573 (
            .O(N__8485),
            .I(N__8482));
    LocalMux I__1572 (
            .O(N__8482),
            .I(N__8479));
    Odrv4 I__1571 (
            .O(N__8479),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_1_1_2 ));
    InMux I__1570 (
            .O(N__8476),
            .I(N__8472));
    InMux I__1569 (
            .O(N__8475),
            .I(N__8469));
    LocalMux I__1568 (
            .O(N__8472),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_4 ));
    LocalMux I__1567 (
            .O(N__8469),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_4 ));
    CascadeMux I__1566 (
            .O(N__8464),
            .I(N__8460));
    CascadeMux I__1565 (
            .O(N__8463),
            .I(N__8456));
    InMux I__1564 (
            .O(N__8460),
            .I(N__8451));
    InMux I__1563 (
            .O(N__8459),
            .I(N__8451));
    InMux I__1562 (
            .O(N__8456),
            .I(N__8448));
    LocalMux I__1561 (
            .O(N__8451),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_4 ));
    LocalMux I__1560 (
            .O(N__8448),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_4 ));
    InMux I__1559 (
            .O(N__8443),
            .I(N__8440));
    LocalMux I__1558 (
            .O(N__8440),
            .I(N__8437));
    Span4Mux_h I__1557 (
            .O(N__8437),
            .I(N__8434));
    Odrv4 I__1556 (
            .O(N__8434),
            .I(\DUT.uart_inst0.rx_countdown_RNO_0Z0Z_2 ));
    InMux I__1555 (
            .O(N__8431),
            .I(N__8427));
    InMux I__1554 (
            .O(N__8430),
            .I(N__8423));
    LocalMux I__1553 (
            .O(N__8427),
            .I(N__8420));
    InMux I__1552 (
            .O(N__8426),
            .I(N__8412));
    LocalMux I__1551 (
            .O(N__8423),
            .I(N__8409));
    Span4Mux_h I__1550 (
            .O(N__8420),
            .I(N__8406));
    InMux I__1549 (
            .O(N__8419),
            .I(N__8401));
    InMux I__1548 (
            .O(N__8418),
            .I(N__8401));
    InMux I__1547 (
            .O(N__8417),
            .I(N__8394));
    InMux I__1546 (
            .O(N__8416),
            .I(N__8394));
    InMux I__1545 (
            .O(N__8415),
            .I(N__8394));
    LocalMux I__1544 (
            .O(N__8412),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_1_2 ));
    Odrv4 I__1543 (
            .O(N__8409),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_1_2 ));
    Odrv4 I__1542 (
            .O(N__8406),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_1_2 ));
    LocalMux I__1541 (
            .O(N__8401),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_1_2 ));
    LocalMux I__1540 (
            .O(N__8394),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_1_2 ));
    CascadeMux I__1539 (
            .O(N__8383),
            .I(N__8380));
    InMux I__1538 (
            .O(N__8380),
            .I(N__8377));
    LocalMux I__1537 (
            .O(N__8377),
            .I(N__8374));
    Odrv4 I__1536 (
            .O(N__8374),
            .I(\DUT.uart_inst0.rx_countdown_RNO_1Z0Z_2 ));
    InMux I__1535 (
            .O(N__8371),
            .I(N__8363));
    InMux I__1534 (
            .O(N__8370),
            .I(N__8360));
    CascadeMux I__1533 (
            .O(N__8369),
            .I(N__8356));
    CascadeMux I__1532 (
            .O(N__8368),
            .I(N__8352));
    CascadeMux I__1531 (
            .O(N__8367),
            .I(N__8349));
    InMux I__1530 (
            .O(N__8366),
            .I(N__8346));
    LocalMux I__1529 (
            .O(N__8363),
            .I(N__8343));
    LocalMux I__1528 (
            .O(N__8360),
            .I(N__8340));
    InMux I__1527 (
            .O(N__8359),
            .I(N__8337));
    InMux I__1526 (
            .O(N__8356),
            .I(N__8332));
    InMux I__1525 (
            .O(N__8355),
            .I(N__8332));
    InMux I__1524 (
            .O(N__8352),
            .I(N__8327));
    InMux I__1523 (
            .O(N__8349),
            .I(N__8327));
    LocalMux I__1522 (
            .O(N__8346),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_2_2 ));
    Odrv4 I__1521 (
            .O(N__8343),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_2_2 ));
    Odrv4 I__1520 (
            .O(N__8340),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_2_2 ));
    LocalMux I__1519 (
            .O(N__8337),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_2_2 ));
    LocalMux I__1518 (
            .O(N__8332),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_2_2 ));
    LocalMux I__1517 (
            .O(N__8327),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_2_2 ));
    InMux I__1516 (
            .O(N__8314),
            .I(N__8310));
    CascadeMux I__1515 (
            .O(N__8313),
            .I(N__8307));
    LocalMux I__1514 (
            .O(N__8310),
            .I(N__8304));
    InMux I__1513 (
            .O(N__8307),
            .I(N__8301));
    Span4Mux_h I__1512 (
            .O(N__8304),
            .I(N__8296));
    LocalMux I__1511 (
            .O(N__8301),
            .I(N__8296));
    Odrv4 I__1510 (
            .O(N__8296),
            .I(\DUT.uart_inst0.rx_countdownZ0Z_2 ));
    CascadeMux I__1509 (
            .O(N__8293),
            .I(N__8285));
    InMux I__1508 (
            .O(N__8292),
            .I(N__8280));
    InMux I__1507 (
            .O(N__8291),
            .I(N__8280));
    InMux I__1506 (
            .O(N__8290),
            .I(N__8275));
    InMux I__1505 (
            .O(N__8289),
            .I(N__8275));
    InMux I__1504 (
            .O(N__8288),
            .I(N__8270));
    InMux I__1503 (
            .O(N__8285),
            .I(N__8270));
    LocalMux I__1502 (
            .O(N__8280),
            .I(\DUT.uart_inst0.recv_stateZ0Z_5 ));
    LocalMux I__1501 (
            .O(N__8275),
            .I(\DUT.uart_inst0.recv_stateZ0Z_5 ));
    LocalMux I__1500 (
            .O(N__8270),
            .I(\DUT.uart_inst0.recv_stateZ0Z_5 ));
    InMux I__1499 (
            .O(N__8263),
            .I(N__8258));
    InMux I__1498 (
            .O(N__8262),
            .I(N__8255));
    InMux I__1497 (
            .O(N__8261),
            .I(N__8252));
    LocalMux I__1496 (
            .O(N__8258),
            .I(N__8249));
    LocalMux I__1495 (
            .O(N__8255),
            .I(\DUT.uart_inst0.recv_stateZ0Z_3 ));
    LocalMux I__1494 (
            .O(N__8252),
            .I(\DUT.uart_inst0.recv_stateZ0Z_3 ));
    Odrv4 I__1493 (
            .O(N__8249),
            .I(\DUT.uart_inst0.recv_stateZ0Z_3 ));
    InMux I__1492 (
            .O(N__8242),
            .I(N__8233));
    InMux I__1491 (
            .O(N__8241),
            .I(N__8233));
    CascadeMux I__1490 (
            .O(N__8240),
            .I(N__8230));
    CascadeMux I__1489 (
            .O(N__8239),
            .I(N__8225));
    InMux I__1488 (
            .O(N__8238),
            .I(N__8220));
    LocalMux I__1487 (
            .O(N__8233),
            .I(N__8217));
    InMux I__1486 (
            .O(N__8230),
            .I(N__8214));
    InMux I__1485 (
            .O(N__8229),
            .I(N__8211));
    InMux I__1484 (
            .O(N__8228),
            .I(N__8206));
    InMux I__1483 (
            .O(N__8225),
            .I(N__8206));
    InMux I__1482 (
            .O(N__8224),
            .I(N__8203));
    InMux I__1481 (
            .O(N__8223),
            .I(N__8200));
    LocalMux I__1480 (
            .O(N__8220),
            .I(N__8197));
    Span4Mux_h I__1479 (
            .O(N__8217),
            .I(N__8184));
    LocalMux I__1478 (
            .O(N__8214),
            .I(N__8184));
    LocalMux I__1477 (
            .O(N__8211),
            .I(N__8184));
    LocalMux I__1476 (
            .O(N__8206),
            .I(N__8184));
    LocalMux I__1475 (
            .O(N__8203),
            .I(N__8184));
    LocalMux I__1474 (
            .O(N__8200),
            .I(N__8184));
    Span4Mux_v I__1473 (
            .O(N__8197),
            .I(N__8180));
    Span4Mux_v I__1472 (
            .O(N__8184),
            .I(N__8177));
    InMux I__1471 (
            .O(N__8183),
            .I(N__8174));
    Sp12to4 I__1470 (
            .O(N__8180),
            .I(N__8167));
    Sp12to4 I__1469 (
            .O(N__8177),
            .I(N__8167));
    LocalMux I__1468 (
            .O(N__8174),
            .I(N__8167));
    Span12Mux_h I__1467 (
            .O(N__8167),
            .I(N__8164));
    Span12Mux_v I__1466 (
            .O(N__8164),
            .I(N__8161));
    Odrv12 I__1465 (
            .O(N__8161),
            .I(P1A1_c));
    InMux I__1464 (
            .O(N__8158),
            .I(N__8147));
    InMux I__1463 (
            .O(N__8157),
            .I(N__8142));
    InMux I__1462 (
            .O(N__8156),
            .I(N__8142));
    InMux I__1461 (
            .O(N__8155),
            .I(N__8139));
    InMux I__1460 (
            .O(N__8154),
            .I(N__8132));
    InMux I__1459 (
            .O(N__8153),
            .I(N__8132));
    InMux I__1458 (
            .O(N__8152),
            .I(N__8132));
    InMux I__1457 (
            .O(N__8151),
            .I(N__8127));
    InMux I__1456 (
            .O(N__8150),
            .I(N__8127));
    LocalMux I__1455 (
            .O(N__8147),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    LocalMux I__1454 (
            .O(N__8142),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    LocalMux I__1453 (
            .O(N__8139),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    LocalMux I__1452 (
            .O(N__8132),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    LocalMux I__1451 (
            .O(N__8127),
            .I(\DUT.uart_inst0.recv_stateZ0Z_1 ));
    InMux I__1450 (
            .O(N__8116),
            .I(N__8113));
    LocalMux I__1449 (
            .O(N__8113),
            .I(N__8110));
    Odrv4 I__1448 (
            .O(N__8110),
            .I(\DUT.uart_inst0.recv_state_srsts_1_5 ));
    InMux I__1447 (
            .O(N__8107),
            .I(N__8104));
    LocalMux I__1446 (
            .O(N__8104),
            .I(N__8100));
    InMux I__1445 (
            .O(N__8103),
            .I(N__8097));
    Odrv4 I__1444 (
            .O(N__8100),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_1 ));
    LocalMux I__1443 (
            .O(N__8097),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_1 ));
    InMux I__1442 (
            .O(N__8092),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_0_s1 ));
    InMux I__1441 (
            .O(N__8089),
            .I(N__8086));
    LocalMux I__1440 (
            .O(N__8086),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_1_s1_THRU_CO ));
    InMux I__1439 (
            .O(N__8083),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_1_s1 ));
    InMux I__1438 (
            .O(N__8080),
            .I(N__8074));
    InMux I__1437 (
            .O(N__8079),
            .I(N__8074));
    LocalMux I__1436 (
            .O(N__8074),
            .I(\DUT.uart_inst0.rx_countdown_3_s1_3 ));
    InMux I__1435 (
            .O(N__8071),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_2_s1 ));
    InMux I__1434 (
            .O(N__8068),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_3_s1 ));
    InMux I__1433 (
            .O(N__8065),
            .I(\DUT.uart_inst0.rx_countdown_3_cry_4_s1 ));
    CascadeMux I__1432 (
            .O(N__8062),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_10_cascade_ ));
    CascadeMux I__1431 (
            .O(N__8059),
            .I(N__8056));
    InMux I__1430 (
            .O(N__8056),
            .I(N__8053));
    LocalMux I__1429 (
            .O(N__8053),
            .I(\DUT.uart_inst0.rx_clk_divider_RNIKU472Z0Z_10 ));
    InMux I__1428 (
            .O(N__8050),
            .I(N__8047));
    LocalMux I__1427 (
            .O(N__8047),
            .I(\DUT.uart_inst0.recv_state_RNO_0Z0Z_0 ));
    CascadeMux I__1426 (
            .O(N__8044),
            .I(\DUT.uart_inst0.recv_state_RNO_1Z0Z_0_cascade_ ));
    InMux I__1425 (
            .O(N__8041),
            .I(N__8031));
    InMux I__1424 (
            .O(N__8040),
            .I(N__8031));
    InMux I__1423 (
            .O(N__8039),
            .I(N__8031));
    InMux I__1422 (
            .O(N__8038),
            .I(N__8028));
    LocalMux I__1421 (
            .O(N__8031),
            .I(\DUT.uart_inst0.recv_stateZ0Z_0 ));
    LocalMux I__1420 (
            .O(N__8028),
            .I(\DUT.uart_inst0.recv_stateZ0Z_0 ));
    InMux I__1419 (
            .O(N__8023),
            .I(N__8020));
    LocalMux I__1418 (
            .O(N__8020),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_a_10 ));
    CascadeMux I__1417 (
            .O(N__8017),
            .I(\DUT.uart_inst0.un2_rx_clk_divider_0_cascade_ ));
    InMux I__1416 (
            .O(N__8014),
            .I(N__8004));
    InMux I__1415 (
            .O(N__8013),
            .I(N__8001));
    InMux I__1414 (
            .O(N__8012),
            .I(N__7998));
    InMux I__1413 (
            .O(N__8011),
            .I(N__7993));
    InMux I__1412 (
            .O(N__8010),
            .I(N__7993));
    InMux I__1411 (
            .O(N__8009),
            .I(N__7986));
    InMux I__1410 (
            .O(N__8008),
            .I(N__7986));
    InMux I__1409 (
            .O(N__8007),
            .I(N__7986));
    LocalMux I__1408 (
            .O(N__8004),
            .I(\DUT.uart_inst0.rx_countdown_3_2 ));
    LocalMux I__1407 (
            .O(N__8001),
            .I(\DUT.uart_inst0.rx_countdown_3_2 ));
    LocalMux I__1406 (
            .O(N__7998),
            .I(\DUT.uart_inst0.rx_countdown_3_2 ));
    LocalMux I__1405 (
            .O(N__7993),
            .I(\DUT.uart_inst0.rx_countdown_3_2 ));
    LocalMux I__1404 (
            .O(N__7986),
            .I(\DUT.uart_inst0.rx_countdown_3_2 ));
    CascadeMux I__1403 (
            .O(N__7975),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_1_2_cascade_ ));
    CascadeMux I__1402 (
            .O(N__7972),
            .I(\DUT.uart_inst0.recv_state_RNO_0Z0Z_4_cascade_ ));
    InMux I__1401 (
            .O(N__7969),
            .I(N__7966));
    LocalMux I__1400 (
            .O(N__7966),
            .I(N__7962));
    InMux I__1399 (
            .O(N__7965),
            .I(N__7959));
    Odrv4 I__1398 (
            .O(N__7962),
            .I(\DUT.uart_inst0.recv_stateZ0Z_4 ));
    LocalMux I__1397 (
            .O(N__7959),
            .I(\DUT.uart_inst0.recv_stateZ0Z_4 ));
    InMux I__1396 (
            .O(N__7954),
            .I(N__7951));
    LocalMux I__1395 (
            .O(N__7951),
            .I(N__7948));
    Odrv4 I__1394 (
            .O(N__7948),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_6 ));
    InMux I__1393 (
            .O(N__7945),
            .I(N__7941));
    InMux I__1392 (
            .O(N__7944),
            .I(N__7938));
    LocalMux I__1391 (
            .O(N__7941),
            .I(N__7933));
    LocalMux I__1390 (
            .O(N__7938),
            .I(N__7930));
    InMux I__1389 (
            .O(N__7937),
            .I(N__7927));
    InMux I__1388 (
            .O(N__7936),
            .I(N__7924));
    Span4Mux_h I__1387 (
            .O(N__7933),
            .I(N__7915));
    Span4Mux_h I__1386 (
            .O(N__7930),
            .I(N__7915));
    LocalMux I__1385 (
            .O(N__7927),
            .I(N__7915));
    LocalMux I__1384 (
            .O(N__7924),
            .I(N__7915));
    Sp12to4 I__1383 (
            .O(N__7915),
            .I(N__7912));
    Odrv12 I__1382 (
            .O(N__7912),
            .I(rTxByteZ0Z_7));
    InMux I__1381 (
            .O(N__7909),
            .I(N__7906));
    LocalMux I__1380 (
            .O(N__7906),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_7 ));
    CEMux I__1379 (
            .O(N__7903),
            .I(N__7900));
    LocalMux I__1378 (
            .O(N__7900),
            .I(N__7897));
    Span4Mux_h I__1377 (
            .O(N__7897),
            .I(N__7893));
    InMux I__1376 (
            .O(N__7896),
            .I(N__7890));
    Odrv4 I__1375 (
            .O(N__7893),
            .I(\DUT.fifo_tx_inst.rFifoData_awe3 ));
    LocalMux I__1374 (
            .O(N__7890),
            .I(\DUT.fifo_tx_inst.rFifoData_awe3 ));
    InMux I__1373 (
            .O(N__7885),
            .I(N__7882));
    LocalMux I__1372 (
            .O(N__7882),
            .I(\DUT.rFifoDatarx_7 ));
    CascadeMux I__1371 (
            .O(N__7879),
            .I(G_152_cascade_));
    CascadeMux I__1370 (
            .O(N__7876),
            .I(N__7873));
    InMux I__1369 (
            .O(N__7873),
            .I(N__7870));
    LocalMux I__1368 (
            .O(N__7870),
            .I(N__7865));
    InMux I__1367 (
            .O(N__7869),
            .I(N__7860));
    InMux I__1366 (
            .O(N__7868),
            .I(N__7860));
    Odrv12 I__1365 (
            .O(N__7865),
            .I(G_151));
    LocalMux I__1364 (
            .O(N__7860),
            .I(G_151));
    CascadeMux I__1363 (
            .O(N__7855),
            .I(N__7852));
    InMux I__1362 (
            .O(N__7852),
            .I(N__7849));
    LocalMux I__1361 (
            .O(N__7849),
            .I(N__7844));
    InMux I__1360 (
            .O(N__7848),
            .I(N__7839));
    InMux I__1359 (
            .O(N__7847),
            .I(N__7839));
    Odrv12 I__1358 (
            .O(N__7844),
            .I(G_150));
    LocalMux I__1357 (
            .O(N__7839),
            .I(G_150));
    InMux I__1356 (
            .O(N__7834),
            .I(N__7829));
    InMux I__1355 (
            .O(N__7833),
            .I(N__7824));
    InMux I__1354 (
            .O(N__7832),
            .I(N__7824));
    LocalMux I__1353 (
            .O(N__7829),
            .I(\fifo_inst.ftdi_input_inst.un1_rWrStateZ0Z_1 ));
    LocalMux I__1352 (
            .O(N__7824),
            .I(\fifo_inst.ftdi_input_inst.un1_rWrStateZ0Z_1 ));
    CascadeMux I__1351 (
            .O(N__7819),
            .I(N__7816));
    InMux I__1350 (
            .O(N__7816),
            .I(N__7813));
    LocalMux I__1349 (
            .O(N__7813),
            .I(N__7807));
    InMux I__1348 (
            .O(N__7812),
            .I(N__7800));
    InMux I__1347 (
            .O(N__7811),
            .I(N__7800));
    InMux I__1346 (
            .O(N__7810),
            .I(N__7800));
    Odrv12 I__1345 (
            .O(N__7807),
            .I(G_149));
    LocalMux I__1344 (
            .O(N__7800),
            .I(G_149));
    InMux I__1343 (
            .O(N__7795),
            .I(N__7792));
    LocalMux I__1342 (
            .O(N__7792),
            .I(\fifo_inst.ftdi_input_inst.un2_oPacketAvail_iZ0 ));
    CascadeMux I__1341 (
            .O(N__7789),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_ ));
    InMux I__1340 (
            .O(N__7786),
            .I(N__7783));
    LocalMux I__1339 (
            .O(N__7783),
            .I(\DUT.uart_inst0.tx_data_RNO_0Z0Z_2 ));
    InMux I__1338 (
            .O(N__7780),
            .I(N__7777));
    LocalMux I__1337 (
            .O(N__7777),
            .I(N__7774));
    Odrv4 I__1336 (
            .O(N__7774),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_0 ));
    InMux I__1335 (
            .O(N__7771),
            .I(N__7768));
    LocalMux I__1334 (
            .O(N__7768),
            .I(N__7763));
    InMux I__1333 (
            .O(N__7767),
            .I(N__7760));
    InMux I__1332 (
            .O(N__7766),
            .I(N__7757));
    Span4Mux_h I__1331 (
            .O(N__7763),
            .I(N__7751));
    LocalMux I__1330 (
            .O(N__7760),
            .I(N__7751));
    LocalMux I__1329 (
            .O(N__7757),
            .I(N__7748));
    InMux I__1328 (
            .O(N__7756),
            .I(N__7745));
    Span4Mux_v I__1327 (
            .O(N__7751),
            .I(N__7742));
    Span4Mux_v I__1326 (
            .O(N__7748),
            .I(N__7737));
    LocalMux I__1325 (
            .O(N__7745),
            .I(N__7737));
    Span4Mux_v I__1324 (
            .O(N__7742),
            .I(N__7734));
    Span4Mux_v I__1323 (
            .O(N__7737),
            .I(N__7731));
    Odrv4 I__1322 (
            .O(N__7734),
            .I(rTxByteZ0Z_2));
    Odrv4 I__1321 (
            .O(N__7731),
            .I(rTxByteZ0Z_2));
    InMux I__1320 (
            .O(N__7726),
            .I(N__7723));
    LocalMux I__1319 (
            .O(N__7723),
            .I(N__7720));
    Odrv4 I__1318 (
            .O(N__7720),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_2 ));
    InMux I__1317 (
            .O(N__7717),
            .I(N__7712));
    InMux I__1316 (
            .O(N__7716),
            .I(N__7709));
    InMux I__1315 (
            .O(N__7715),
            .I(N__7706));
    LocalMux I__1314 (
            .O(N__7712),
            .I(N__7702));
    LocalMux I__1313 (
            .O(N__7709),
            .I(N__7697));
    LocalMux I__1312 (
            .O(N__7706),
            .I(N__7697));
    InMux I__1311 (
            .O(N__7705),
            .I(N__7694));
    Span4Mux_v I__1310 (
            .O(N__7702),
            .I(N__7691));
    Span4Mux_v I__1309 (
            .O(N__7697),
            .I(N__7686));
    LocalMux I__1308 (
            .O(N__7694),
            .I(N__7686));
    Span4Mux_v I__1307 (
            .O(N__7691),
            .I(N__7683));
    Span4Mux_v I__1306 (
            .O(N__7686),
            .I(N__7680));
    Odrv4 I__1305 (
            .O(N__7683),
            .I(rTxByteZ0Z_4));
    Odrv4 I__1304 (
            .O(N__7680),
            .I(rTxByteZ0Z_4));
    CascadeMux I__1303 (
            .O(N__7675),
            .I(N__7672));
    InMux I__1302 (
            .O(N__7672),
            .I(N__7669));
    LocalMux I__1301 (
            .O(N__7669),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_4 ));
    InMux I__1300 (
            .O(N__7666),
            .I(N__7663));
    LocalMux I__1299 (
            .O(N__7663),
            .I(N__7657));
    InMux I__1298 (
            .O(N__7662),
            .I(N__7654));
    InMux I__1297 (
            .O(N__7661),
            .I(N__7651));
    InMux I__1296 (
            .O(N__7660),
            .I(N__7648));
    Span4Mux_h I__1295 (
            .O(N__7657),
            .I(N__7639));
    LocalMux I__1294 (
            .O(N__7654),
            .I(N__7639));
    LocalMux I__1293 (
            .O(N__7651),
            .I(N__7639));
    LocalMux I__1292 (
            .O(N__7648),
            .I(N__7639));
    Span4Mux_v I__1291 (
            .O(N__7639),
            .I(N__7636));
    Odrv4 I__1290 (
            .O(N__7636),
            .I(rTxByteZ0Z_5));
    InMux I__1289 (
            .O(N__7633),
            .I(N__7630));
    LocalMux I__1288 (
            .O(N__7630),
            .I(N__7627));
    Odrv4 I__1287 (
            .O(N__7627),
            .I(\DUT.fifo_tx_inst.rFifoData_ram3_5 ));
    CascadeMux I__1286 (
            .O(N__7624),
            .I(\DUT.uart_inst0.g0_i_o4_0_4_cascade_ ));
    CascadeMux I__1285 (
            .O(N__7621),
            .I(N__7616));
    InMux I__1284 (
            .O(N__7620),
            .I(N__7613));
    InMux I__1283 (
            .O(N__7619),
            .I(N__7605));
    InMux I__1282 (
            .O(N__7616),
            .I(N__7602));
    LocalMux I__1281 (
            .O(N__7613),
            .I(N__7599));
    InMux I__1280 (
            .O(N__7612),
            .I(N__7596));
    InMux I__1279 (
            .O(N__7611),
            .I(N__7591));
    InMux I__1278 (
            .O(N__7610),
            .I(N__7591));
    InMux I__1277 (
            .O(N__7609),
            .I(N__7588));
    InMux I__1276 (
            .O(N__7608),
            .I(N__7585));
    LocalMux I__1275 (
            .O(N__7605),
            .I(N__7582));
    LocalMux I__1274 (
            .O(N__7602),
            .I(N__7575));
    Span4Mux_v I__1273 (
            .O(N__7599),
            .I(N__7575));
    LocalMux I__1272 (
            .O(N__7596),
            .I(N__7575));
    LocalMux I__1271 (
            .O(N__7591),
            .I(N__7569));
    LocalMux I__1270 (
            .O(N__7588),
            .I(N__7569));
    LocalMux I__1269 (
            .O(N__7585),
            .I(N__7564));
    Span4Mux_v I__1268 (
            .O(N__7582),
            .I(N__7564));
    Span4Mux_v I__1267 (
            .O(N__7575),
            .I(N__7561));
    InMux I__1266 (
            .O(N__7574),
            .I(N__7558));
    Odrv12 I__1265 (
            .O(N__7569),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_1 ));
    Odrv4 I__1264 (
            .O(N__7564),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_1 ));
    Odrv4 I__1263 (
            .O(N__7561),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_1 ));
    LocalMux I__1262 (
            .O(N__7558),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_1 ));
    CascadeMux I__1261 (
            .O(N__7549),
            .I(N__7542));
    InMux I__1260 (
            .O(N__7548),
            .I(N__7538));
    CascadeMux I__1259 (
            .O(N__7547),
            .I(N__7535));
    CascadeMux I__1258 (
            .O(N__7546),
            .I(N__7532));
    InMux I__1257 (
            .O(N__7545),
            .I(N__7529));
    InMux I__1256 (
            .O(N__7542),
            .I(N__7525));
    InMux I__1255 (
            .O(N__7541),
            .I(N__7522));
    LocalMux I__1254 (
            .O(N__7538),
            .I(N__7519));
    InMux I__1253 (
            .O(N__7535),
            .I(N__7514));
    InMux I__1252 (
            .O(N__7532),
            .I(N__7514));
    LocalMux I__1251 (
            .O(N__7529),
            .I(N__7511));
    InMux I__1250 (
            .O(N__7528),
            .I(N__7508));
    LocalMux I__1249 (
            .O(N__7525),
            .I(N__7505));
    LocalMux I__1248 (
            .O(N__7522),
            .I(N__7497));
    Span4Mux_v I__1247 (
            .O(N__7519),
            .I(N__7497));
    LocalMux I__1246 (
            .O(N__7514),
            .I(N__7488));
    Span4Mux_v I__1245 (
            .O(N__7511),
            .I(N__7488));
    LocalMux I__1244 (
            .O(N__7508),
            .I(N__7488));
    Span4Mux_h I__1243 (
            .O(N__7505),
            .I(N__7488));
    InMux I__1242 (
            .O(N__7504),
            .I(N__7481));
    InMux I__1241 (
            .O(N__7503),
            .I(N__7481));
    InMux I__1240 (
            .O(N__7502),
            .I(N__7481));
    Odrv4 I__1239 (
            .O(N__7497),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_0 ));
    Odrv4 I__1238 (
            .O(N__7488),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_0 ));
    LocalMux I__1237 (
            .O(N__7481),
            .I(\DUT.fifo_tx_inst.rWritePtrZ0Z_0 ));
    InMux I__1236 (
            .O(N__7474),
            .I(N__7467));
    InMux I__1235 (
            .O(N__7473),
            .I(N__7464));
    InMux I__1234 (
            .O(N__7472),
            .I(N__7457));
    InMux I__1233 (
            .O(N__7471),
            .I(N__7457));
    InMux I__1232 (
            .O(N__7470),
            .I(N__7457));
    LocalMux I__1231 (
            .O(N__7467),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_2 ));
    LocalMux I__1230 (
            .O(N__7464),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_2 ));
    LocalMux I__1229 (
            .O(N__7457),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_2 ));
    InMux I__1228 (
            .O(N__7450),
            .I(N__7447));
    LocalMux I__1227 (
            .O(N__7447),
            .I(\DUT.rFifoDatarxZ0Z_0 ));
    InMux I__1226 (
            .O(N__7444),
            .I(N__7441));
    LocalMux I__1225 (
            .O(N__7441),
            .I(N__7438));
    Span4Mux_h I__1224 (
            .O(N__7438),
            .I(N__7435));
    Odrv4 I__1223 (
            .O(N__7435),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_4 ));
    InMux I__1222 (
            .O(N__7432),
            .I(N__7429));
    LocalMux I__1221 (
            .O(N__7429),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4 ));
    CascadeMux I__1220 (
            .O(N__7426),
            .I(\DUT.rFifoDatarx_4_cascade_ ));
    InMux I__1219 (
            .O(N__7423),
            .I(N__7420));
    LocalMux I__1218 (
            .O(N__7420),
            .I(\DUT.uart_inst0.tx_data_RNO_0Z0Z_4 ));
    InMux I__1217 (
            .O(N__7417),
            .I(N__7414));
    LocalMux I__1216 (
            .O(N__7414),
            .I(N__7411));
    Span4Mux_v I__1215 (
            .O(N__7411),
            .I(N__7408));
    Odrv4 I__1214 (
            .O(N__7408),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_6 ));
    CascadeMux I__1213 (
            .O(N__7405),
            .I(N__7402));
    InMux I__1212 (
            .O(N__7402),
            .I(N__7399));
    LocalMux I__1211 (
            .O(N__7399),
            .I(N__7396));
    Odrv4 I__1210 (
            .O(N__7396),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_6 ));
    CascadeMux I__1209 (
            .O(N__7393),
            .I(N__7387));
    InMux I__1208 (
            .O(N__7392),
            .I(N__7377));
    InMux I__1207 (
            .O(N__7391),
            .I(N__7374));
    InMux I__1206 (
            .O(N__7390),
            .I(N__7367));
    InMux I__1205 (
            .O(N__7387),
            .I(N__7367));
    InMux I__1204 (
            .O(N__7386),
            .I(N__7367));
    InMux I__1203 (
            .O(N__7385),
            .I(N__7362));
    InMux I__1202 (
            .O(N__7384),
            .I(N__7362));
    InMux I__1201 (
            .O(N__7383),
            .I(N__7353));
    InMux I__1200 (
            .O(N__7382),
            .I(N__7353));
    InMux I__1199 (
            .O(N__7381),
            .I(N__7353));
    InMux I__1198 (
            .O(N__7380),
            .I(N__7353));
    LocalMux I__1197 (
            .O(N__7377),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__1196 (
            .O(N__7374),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__1195 (
            .O(N__7367),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__1194 (
            .O(N__7362),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__1193 (
            .O(N__7353),
            .I(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ));
    InMux I__1192 (
            .O(N__7342),
            .I(N__7339));
    LocalMux I__1191 (
            .O(N__7339),
            .I(\DUT.uart_inst0.tx_countdown_0_c3 ));
    InMux I__1190 (
            .O(N__7336),
            .I(N__7333));
    LocalMux I__1189 (
            .O(N__7333),
            .I(\DUT.uart_inst0.un1_m7_3 ));
    CascadeMux I__1188 (
            .O(N__7330),
            .I(\DUT.uart_inst0.un1_tx_state_0_a4_1_cascade_ ));
    CascadeMux I__1187 (
            .O(N__7327),
            .I(\DUT.uart_inst0.un1_tx_clk_divider_s1_sn_0_cascade_ ));
    InMux I__1186 (
            .O(N__7324),
            .I(N__7321));
    LocalMux I__1185 (
            .O(N__7321),
            .I(\DUT.uart_inst0.tx_countdown_7_1_0_3 ));
    CascadeMux I__1184 (
            .O(N__7318),
            .I(\DUT.uart_inst0.tx_countdown_RNO_0Z0Z_1_cascade_ ));
    CascadeMux I__1183 (
            .O(N__7315),
            .I(\DUT.uart_inst0.N_98_4_cascade_ ));
    InMux I__1182 (
            .O(N__7312),
            .I(N__7308));
    InMux I__1181 (
            .O(N__7311),
            .I(N__7305));
    LocalMux I__1180 (
            .O(N__7308),
            .I(N__7302));
    LocalMux I__1179 (
            .O(N__7305),
            .I(\DUT.uart_inst0.rx_m2_e_0 ));
    Odrv4 I__1178 (
            .O(N__7302),
            .I(\DUT.uart_inst0.rx_m2_e_0 ));
    CascadeMux I__1177 (
            .O(N__7297),
            .I(\DUT.uart_inst0.r_N_5_mux_cascade_ ));
    InMux I__1176 (
            .O(N__7294),
            .I(N__7281));
    InMux I__1175 (
            .O(N__7293),
            .I(N__7281));
    InMux I__1174 (
            .O(N__7292),
            .I(N__7281));
    InMux I__1173 (
            .O(N__7291),
            .I(N__7281));
    InMux I__1172 (
            .O(N__7290),
            .I(N__7278));
    LocalMux I__1171 (
            .O(N__7281),
            .I(\DUT.uart_inst0.recv_stateZ0Z_2 ));
    LocalMux I__1170 (
            .O(N__7278),
            .I(\DUT.uart_inst0.recv_stateZ0Z_2 ));
    InMux I__1169 (
            .O(N__7273),
            .I(N__7270));
    LocalMux I__1168 (
            .O(N__7270),
            .I(\DUT.uart_inst0.N_98_4 ));
    CascadeMux I__1167 (
            .O(N__7267),
            .I(\DUT.uart_inst0.r_N_3_mux_cascade_ ));
    InMux I__1166 (
            .O(N__7264),
            .I(N__7258));
    InMux I__1165 (
            .O(N__7263),
            .I(N__7258));
    LocalMux I__1164 (
            .O(N__7258),
            .I(\DUT.uart_inst0.recv_N_5_mux ));
    CascadeMux I__1163 (
            .O(N__7255),
            .I(\DUT.uart_inst0.g3_cascade_ ));
    CascadeMux I__1162 (
            .O(N__7252),
            .I(N__7249));
    InMux I__1161 (
            .O(N__7249),
            .I(N__7246));
    LocalMux I__1160 (
            .O(N__7246),
            .I(\DUT.uart_inst0.g3_1 ));
    CascadeMux I__1159 (
            .O(N__7243),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_2_2_cascade_ ));
    CascadeMux I__1158 (
            .O(N__7240),
            .I(\DUT.uart_inst0.recv_state_RNO_0Z0Z_1_cascade_ ));
    CascadeMux I__1157 (
            .O(N__7237),
            .I(\DUT.uart_inst0.un1_m2_e_0_cascade_ ));
    CascadeMux I__1156 (
            .O(N__7234),
            .I(N__7230));
    InMux I__1155 (
            .O(N__7233),
            .I(N__7227));
    InMux I__1154 (
            .O(N__7230),
            .I(N__7224));
    LocalMux I__1153 (
            .O(N__7227),
            .I(N__7221));
    LocalMux I__1152 (
            .O(N__7224),
            .I(\DUT.uart_inst0.N_69 ));
    Odrv4 I__1151 (
            .O(N__7221),
            .I(\DUT.uart_inst0.N_69 ));
    CascadeMux I__1150 (
            .O(N__7216),
            .I(\DUT.uart_inst0.recv_state_RNITN8GJZ0Z_2_cascade_ ));
    CEMux I__1149 (
            .O(N__7213),
            .I(N__7210));
    LocalMux I__1148 (
            .O(N__7210),
            .I(N__7207));
    Span4Mux_h I__1147 (
            .O(N__7207),
            .I(N__7203));
    InMux I__1146 (
            .O(N__7206),
            .I(N__7200));
    Odrv4 I__1145 (
            .O(N__7203),
            .I(\DUT.uart_inst0.recv_state_RNITN8GJZ0Z_2 ));
    LocalMux I__1144 (
            .O(N__7200),
            .I(\DUT.uart_inst0.recv_state_RNITN8GJZ0Z_2 ));
    InMux I__1143 (
            .O(N__7195),
            .I(N__7190));
    InMux I__1142 (
            .O(N__7194),
            .I(N__7187));
    InMux I__1141 (
            .O(N__7193),
            .I(N__7184));
    LocalMux I__1140 (
            .O(N__7190),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_2 ));
    LocalMux I__1139 (
            .O(N__7187),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_2 ));
    LocalMux I__1138 (
            .O(N__7184),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_2 ));
    InMux I__1137 (
            .O(N__7177),
            .I(N__7173));
    CascadeMux I__1136 (
            .O(N__7176),
            .I(N__7170));
    LocalMux I__1135 (
            .O(N__7173),
            .I(N__7166));
    InMux I__1134 (
            .O(N__7170),
            .I(N__7161));
    InMux I__1133 (
            .O(N__7169),
            .I(N__7161));
    Odrv4 I__1132 (
            .O(N__7166),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_1 ));
    LocalMux I__1131 (
            .O(N__7161),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_1 ));
    CascadeMux I__1130 (
            .O(N__7156),
            .I(N__7153));
    InMux I__1129 (
            .O(N__7153),
            .I(N__7149));
    InMux I__1128 (
            .O(N__7152),
            .I(N__7146));
    LocalMux I__1127 (
            .O(N__7149),
            .I(N__7143));
    LocalMux I__1126 (
            .O(N__7146),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_3 ));
    Odrv4 I__1125 (
            .O(N__7143),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_3 ));
    InMux I__1124 (
            .O(N__7138),
            .I(N__7132));
    InMux I__1123 (
            .O(N__7137),
            .I(N__7127));
    InMux I__1122 (
            .O(N__7136),
            .I(N__7127));
    InMux I__1121 (
            .O(N__7135),
            .I(N__7124));
    LocalMux I__1120 (
            .O(N__7132),
            .I(N__7119));
    LocalMux I__1119 (
            .O(N__7127),
            .I(N__7119));
    LocalMux I__1118 (
            .O(N__7124),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_0 ));
    Odrv4 I__1117 (
            .O(N__7119),
            .I(\DUT.uart_inst0.rx_bits_remainingZ0Z_0 ));
    CEMux I__1116 (
            .O(N__7114),
            .I(N__7111));
    LocalMux I__1115 (
            .O(N__7111),
            .I(N__7108));
    Odrv12 I__1114 (
            .O(N__7108),
            .I(\DUT.uart_inst0.rx_bits_remaining_2_sqmuxa ));
    CascadeMux I__1113 (
            .O(N__7105),
            .I(\DUT.uart_inst0.rx_countdown_3_2_cascade_ ));
    CascadeMux I__1112 (
            .O(N__7102),
            .I(N__7097));
    InMux I__1111 (
            .O(N__7101),
            .I(N__7094));
    InMux I__1110 (
            .O(N__7100),
            .I(N__7088));
    InMux I__1109 (
            .O(N__7097),
            .I(N__7085));
    LocalMux I__1108 (
            .O(N__7094),
            .I(N__7082));
    InMux I__1107 (
            .O(N__7093),
            .I(N__7079));
    InMux I__1106 (
            .O(N__7092),
            .I(N__7074));
    InMux I__1105 (
            .O(N__7091),
            .I(N__7074));
    LocalMux I__1104 (
            .O(N__7088),
            .I(\DUT.wRcvd ));
    LocalMux I__1103 (
            .O(N__7085),
            .I(\DUT.wRcvd ));
    Odrv4 I__1102 (
            .O(N__7082),
            .I(\DUT.wRcvd ));
    LocalMux I__1101 (
            .O(N__7079),
            .I(\DUT.wRcvd ));
    LocalMux I__1100 (
            .O(N__7074),
            .I(\DUT.wRcvd ));
    CascadeMux I__1099 (
            .O(N__7063),
            .I(\DUT.uart_inst0.rx_countdown_8_i_o2_2_1_2_cascade_ ));
    CascadeMux I__1098 (
            .O(N__7060),
            .I(N__7057));
    InMux I__1097 (
            .O(N__7057),
            .I(N__7054));
    LocalMux I__1096 (
            .O(N__7054),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_7 ));
    CEMux I__1095 (
            .O(N__7051),
            .I(N__7048));
    LocalMux I__1094 (
            .O(N__7048),
            .I(N__7045));
    Span4Mux_h I__1093 (
            .O(N__7045),
            .I(N__7042));
    Span4Mux_h I__1092 (
            .O(N__7042),
            .I(N__7039));
    Odrv4 I__1091 (
            .O(N__7039),
            .I(\DUT.fifo_rx_inst.rFifoData_awe1 ));
    InMux I__1090 (
            .O(N__7036),
            .I(N__7033));
    LocalMux I__1089 (
            .O(N__7033),
            .I(N__7028));
    InMux I__1088 (
            .O(N__7032),
            .I(N__7025));
    InMux I__1087 (
            .O(N__7031),
            .I(N__7021));
    Span4Mux_v I__1086 (
            .O(N__7028),
            .I(N__7016));
    LocalMux I__1085 (
            .O(N__7025),
            .I(N__7016));
    InMux I__1084 (
            .O(N__7024),
            .I(N__7013));
    LocalMux I__1083 (
            .O(N__7021),
            .I(\DUT.wRxByte_0 ));
    Odrv4 I__1082 (
            .O(N__7016),
            .I(\DUT.wRxByte_0 ));
    LocalMux I__1081 (
            .O(N__7013),
            .I(\DUT.wRxByte_0 ));
    InMux I__1080 (
            .O(N__7006),
            .I(N__7003));
    LocalMux I__1079 (
            .O(N__7003),
            .I(N__6998));
    InMux I__1078 (
            .O(N__7002),
            .I(N__6995));
    InMux I__1077 (
            .O(N__7001),
            .I(N__6990));
    Span4Mux_v I__1076 (
            .O(N__6998),
            .I(N__6985));
    LocalMux I__1075 (
            .O(N__6995),
            .I(N__6985));
    InMux I__1074 (
            .O(N__6994),
            .I(N__6982));
    InMux I__1073 (
            .O(N__6993),
            .I(N__6979));
    LocalMux I__1072 (
            .O(N__6990),
            .I(\DUT.wRxByte_1 ));
    Odrv4 I__1071 (
            .O(N__6985),
            .I(\DUT.wRxByte_1 ));
    LocalMux I__1070 (
            .O(N__6982),
            .I(\DUT.wRxByte_1 ));
    LocalMux I__1069 (
            .O(N__6979),
            .I(\DUT.wRxByte_1 ));
    InMux I__1068 (
            .O(N__6970),
            .I(N__6967));
    LocalMux I__1067 (
            .O(N__6967),
            .I(N__6962));
    InMux I__1066 (
            .O(N__6966),
            .I(N__6959));
    InMux I__1065 (
            .O(N__6965),
            .I(N__6956));
    Span4Mux_h I__1064 (
            .O(N__6962),
            .I(N__6951));
    LocalMux I__1063 (
            .O(N__6959),
            .I(N__6946));
    LocalMux I__1062 (
            .O(N__6956),
            .I(N__6946));
    InMux I__1061 (
            .O(N__6955),
            .I(N__6943));
    InMux I__1060 (
            .O(N__6954),
            .I(N__6940));
    Odrv4 I__1059 (
            .O(N__6951),
            .I(\DUT.wRxByte_2 ));
    Odrv4 I__1058 (
            .O(N__6946),
            .I(\DUT.wRxByte_2 ));
    LocalMux I__1057 (
            .O(N__6943),
            .I(\DUT.wRxByte_2 ));
    LocalMux I__1056 (
            .O(N__6940),
            .I(\DUT.wRxByte_2 ));
    InMux I__1055 (
            .O(N__6931),
            .I(N__6927));
    InMux I__1054 (
            .O(N__6930),
            .I(N__6924));
    LocalMux I__1053 (
            .O(N__6927),
            .I(N__6920));
    LocalMux I__1052 (
            .O(N__6924),
            .I(N__6917));
    InMux I__1051 (
            .O(N__6923),
            .I(N__6914));
    Span4Mux_h I__1050 (
            .O(N__6920),
            .I(N__6909));
    Span4Mux_v I__1049 (
            .O(N__6917),
            .I(N__6904));
    LocalMux I__1048 (
            .O(N__6914),
            .I(N__6904));
    InMux I__1047 (
            .O(N__6913),
            .I(N__6901));
    InMux I__1046 (
            .O(N__6912),
            .I(N__6898));
    Odrv4 I__1045 (
            .O(N__6909),
            .I(\DUT.wRxByte_3 ));
    Odrv4 I__1044 (
            .O(N__6904),
            .I(\DUT.wRxByte_3 ));
    LocalMux I__1043 (
            .O(N__6901),
            .I(\DUT.wRxByte_3 ));
    LocalMux I__1042 (
            .O(N__6898),
            .I(\DUT.wRxByte_3 ));
    InMux I__1041 (
            .O(N__6889),
            .I(N__6885));
    InMux I__1040 (
            .O(N__6888),
            .I(N__6882));
    LocalMux I__1039 (
            .O(N__6885),
            .I(N__6878));
    LocalMux I__1038 (
            .O(N__6882),
            .I(N__6875));
    InMux I__1037 (
            .O(N__6881),
            .I(N__6872));
    Span4Mux_v I__1036 (
            .O(N__6878),
            .I(N__6863));
    Span4Mux_v I__1035 (
            .O(N__6875),
            .I(N__6863));
    LocalMux I__1034 (
            .O(N__6872),
            .I(N__6863));
    InMux I__1033 (
            .O(N__6871),
            .I(N__6860));
    InMux I__1032 (
            .O(N__6870),
            .I(N__6857));
    Odrv4 I__1031 (
            .O(N__6863),
            .I(\DUT.wRxByte_4 ));
    LocalMux I__1030 (
            .O(N__6860),
            .I(\DUT.wRxByte_4 ));
    LocalMux I__1029 (
            .O(N__6857),
            .I(\DUT.wRxByte_4 ));
    InMux I__1028 (
            .O(N__6850),
            .I(N__6846));
    InMux I__1027 (
            .O(N__6849),
            .I(N__6843));
    LocalMux I__1026 (
            .O(N__6846),
            .I(N__6839));
    LocalMux I__1025 (
            .O(N__6843),
            .I(N__6836));
    InMux I__1024 (
            .O(N__6842),
            .I(N__6833));
    Span4Mux_v I__1023 (
            .O(N__6839),
            .I(N__6824));
    Span4Mux_v I__1022 (
            .O(N__6836),
            .I(N__6824));
    LocalMux I__1021 (
            .O(N__6833),
            .I(N__6824));
    InMux I__1020 (
            .O(N__6832),
            .I(N__6821));
    InMux I__1019 (
            .O(N__6831),
            .I(N__6818));
    Odrv4 I__1018 (
            .O(N__6824),
            .I(\DUT.wRxByte_5 ));
    LocalMux I__1017 (
            .O(N__6821),
            .I(\DUT.wRxByte_5 ));
    LocalMux I__1016 (
            .O(N__6818),
            .I(\DUT.wRxByte_5 ));
    InMux I__1015 (
            .O(N__6811),
            .I(N__6807));
    InMux I__1014 (
            .O(N__6810),
            .I(N__6804));
    LocalMux I__1013 (
            .O(N__6807),
            .I(N__6800));
    LocalMux I__1012 (
            .O(N__6804),
            .I(N__6797));
    InMux I__1011 (
            .O(N__6803),
            .I(N__6794));
    Span4Mux_v I__1010 (
            .O(N__6800),
            .I(N__6785));
    Span4Mux_v I__1009 (
            .O(N__6797),
            .I(N__6785));
    LocalMux I__1008 (
            .O(N__6794),
            .I(N__6785));
    InMux I__1007 (
            .O(N__6793),
            .I(N__6782));
    InMux I__1006 (
            .O(N__6792),
            .I(N__6779));
    Odrv4 I__1005 (
            .O(N__6785),
            .I(\DUT.wRxByte_6 ));
    LocalMux I__1004 (
            .O(N__6782),
            .I(\DUT.wRxByte_6 ));
    LocalMux I__1003 (
            .O(N__6779),
            .I(\DUT.wRxByte_6 ));
    InMux I__1002 (
            .O(N__6772),
            .I(N__6769));
    LocalMux I__1001 (
            .O(N__6769),
            .I(N__6765));
    InMux I__1000 (
            .O(N__6768),
            .I(N__6761));
    Span4Mux_h I__999 (
            .O(N__6765),
            .I(N__6756));
    InMux I__998 (
            .O(N__6764),
            .I(N__6753));
    LocalMux I__997 (
            .O(N__6761),
            .I(N__6750));
    InMux I__996 (
            .O(N__6760),
            .I(N__6747));
    InMux I__995 (
            .O(N__6759),
            .I(N__6744));
    Odrv4 I__994 (
            .O(N__6756),
            .I(\DUT.wRxByte_7 ));
    LocalMux I__993 (
            .O(N__6753),
            .I(\DUT.wRxByte_7 ));
    Odrv4 I__992 (
            .O(N__6750),
            .I(\DUT.wRxByte_7 ));
    LocalMux I__991 (
            .O(N__6747),
            .I(\DUT.wRxByte_7 ));
    LocalMux I__990 (
            .O(N__6744),
            .I(\DUT.wRxByte_7 ));
    CascadeMux I__989 (
            .O(N__6733),
            .I(G_141_cascade_));
    CascadeMux I__988 (
            .O(N__6730),
            .I(N__6726));
    CascadeMux I__987 (
            .O(N__6729),
            .I(N__6722));
    InMux I__986 (
            .O(N__6726),
            .I(N__6715));
    InMux I__985 (
            .O(N__6725),
            .I(N__6715));
    InMux I__984 (
            .O(N__6722),
            .I(N__6708));
    InMux I__983 (
            .O(N__6721),
            .I(N__6708));
    InMux I__982 (
            .O(N__6720),
            .I(N__6708));
    LocalMux I__981 (
            .O(N__6715),
            .I(G_140));
    LocalMux I__980 (
            .O(N__6708),
            .I(G_140));
    InMux I__979 (
            .O(N__6703),
            .I(N__6700));
    LocalMux I__978 (
            .O(N__6700),
            .I(fifo_inst_ftdi_input_inst_oTxFull_0));
    CascadeMux I__977 (
            .O(N__6697),
            .I(G_140_cascade_));
    InMux I__976 (
            .O(N__6694),
            .I(N__6684));
    InMux I__975 (
            .O(N__6693),
            .I(N__6684));
    InMux I__974 (
            .O(N__6692),
            .I(N__6684));
    InMux I__973 (
            .O(N__6691),
            .I(N__6681));
    LocalMux I__972 (
            .O(N__6684),
            .I(G_143));
    LocalMux I__971 (
            .O(N__6681),
            .I(G_143));
    InMux I__970 (
            .O(N__6676),
            .I(N__6667));
    InMux I__969 (
            .O(N__6675),
            .I(N__6667));
    InMux I__968 (
            .O(N__6674),
            .I(N__6667));
    LocalMux I__967 (
            .O(N__6667),
            .I(G_146));
    InMux I__966 (
            .O(N__6664),
            .I(N__6661));
    LocalMux I__965 (
            .O(N__6661),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_0 ));
    CascadeMux I__964 (
            .O(N__6658),
            .I(N__6655));
    InMux I__963 (
            .O(N__6655),
            .I(N__6652));
    LocalMux I__962 (
            .O(N__6652),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_1 ));
    CascadeMux I__961 (
            .O(N__6649),
            .I(N__6646));
    InMux I__960 (
            .O(N__6646),
            .I(N__6643));
    LocalMux I__959 (
            .O(N__6643),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_2 ));
    CascadeMux I__958 (
            .O(N__6640),
            .I(N__6637));
    InMux I__957 (
            .O(N__6637),
            .I(N__6634));
    LocalMux I__956 (
            .O(N__6634),
            .I(N__6631));
    Span4Mux_v I__955 (
            .O(N__6631),
            .I(N__6628));
    Odrv4 I__954 (
            .O(N__6628),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_3 ));
    CascadeMux I__953 (
            .O(N__6625),
            .I(N__6622));
    InMux I__952 (
            .O(N__6622),
            .I(N__6619));
    LocalMux I__951 (
            .O(N__6619),
            .I(N__6616));
    Span4Mux_h I__950 (
            .O(N__6616),
            .I(N__6613));
    Odrv4 I__949 (
            .O(N__6613),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_4 ));
    CascadeMux I__948 (
            .O(N__6610),
            .I(N__6607));
    InMux I__947 (
            .O(N__6607),
            .I(N__6604));
    LocalMux I__946 (
            .O(N__6604),
            .I(N__6601));
    Span4Mux_h I__945 (
            .O(N__6601),
            .I(N__6598));
    Odrv4 I__944 (
            .O(N__6598),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_5 ));
    CascadeMux I__943 (
            .O(N__6595),
            .I(N__6592));
    InMux I__942 (
            .O(N__6592),
            .I(N__6589));
    LocalMux I__941 (
            .O(N__6589),
            .I(N__6586));
    Span4Mux_h I__940 (
            .O(N__6586),
            .I(N__6583));
    Odrv4 I__939 (
            .O(N__6583),
            .I(\DUT.fifo_rx_inst.rFifoData_ram1_6 ));
    CEMux I__938 (
            .O(N__6580),
            .I(N__6576));
    CEMux I__937 (
            .O(N__6579),
            .I(N__6573));
    LocalMux I__936 (
            .O(N__6576),
            .I(\DUT.fifo_tx_inst.N_40 ));
    LocalMux I__935 (
            .O(N__6573),
            .I(\DUT.fifo_tx_inst.N_40 ));
    CascadeMux I__934 (
            .O(N__6568),
            .I(G_145_cascade_));
    InMux I__933 (
            .O(N__6565),
            .I(N__6559));
    InMux I__932 (
            .O(N__6564),
            .I(N__6559));
    LocalMux I__931 (
            .O(N__6559),
            .I(G_145));
    CascadeMux I__930 (
            .O(N__6556),
            .I(G_142_cascade_));
    InMux I__929 (
            .O(N__6553),
            .I(N__6542));
    InMux I__928 (
            .O(N__6552),
            .I(N__6542));
    InMux I__927 (
            .O(N__6551),
            .I(N__6542));
    InMux I__926 (
            .O(N__6550),
            .I(N__6539));
    InMux I__925 (
            .O(N__6549),
            .I(N__6536));
    LocalMux I__924 (
            .O(N__6542),
            .I(G_144));
    LocalMux I__923 (
            .O(N__6539),
            .I(G_144));
    LocalMux I__922 (
            .O(N__6536),
            .I(G_144));
    InMux I__921 (
            .O(N__6529),
            .I(N__6526));
    LocalMux I__920 (
            .O(N__6526),
            .I(\fifo_inst.ftdi_input_inst.SUMZ0Z_3 ));
    SRMux I__919 (
            .O(N__6523),
            .I(N__6520));
    LocalMux I__918 (
            .O(N__6520),
            .I(N__6517));
    Span4Mux_h I__917 (
            .O(N__6517),
            .I(N__6512));
    InMux I__916 (
            .O(N__6516),
            .I(N__6509));
    InMux I__915 (
            .O(N__6515),
            .I(N__6506));
    Odrv4 I__914 (
            .O(N__6512),
            .I(G_147));
    LocalMux I__913 (
            .O(N__6509),
            .I(G_147));
    LocalMux I__912 (
            .O(N__6506),
            .I(G_147));
    CascadeMux I__911 (
            .O(N__6499),
            .I(N__6493));
    InMux I__910 (
            .O(N__6498),
            .I(N__6484));
    InMux I__909 (
            .O(N__6497),
            .I(N__6484));
    InMux I__908 (
            .O(N__6496),
            .I(N__6484));
    InMux I__907 (
            .O(N__6493),
            .I(N__6484));
    LocalMux I__906 (
            .O(N__6484),
            .I(G_142));
    InMux I__905 (
            .O(N__6481),
            .I(N__6474));
    InMux I__904 (
            .O(N__6480),
            .I(N__6474));
    InMux I__903 (
            .O(N__6479),
            .I(N__6471));
    LocalMux I__902 (
            .O(N__6474),
            .I(G_141));
    LocalMux I__901 (
            .O(N__6471),
            .I(G_141));
    InMux I__900 (
            .O(N__6466),
            .I(N__6463));
    LocalMux I__899 (
            .O(N__6463),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_5 ));
    CascadeMux I__898 (
            .O(N__6460),
            .I(N__6457));
    InMux I__897 (
            .O(N__6457),
            .I(N__6454));
    LocalMux I__896 (
            .O(N__6454),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_5 ));
    CascadeMux I__895 (
            .O(N__6451),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ));
    InMux I__894 (
            .O(N__6448),
            .I(N__6445));
    LocalMux I__893 (
            .O(N__6445),
            .I(N__6442));
    Odrv4 I__892 (
            .O(N__6442),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_5 ));
    InMux I__891 (
            .O(N__6439),
            .I(N__6436));
    LocalMux I__890 (
            .O(N__6436),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_7 ));
    InMux I__889 (
            .O(N__6433),
            .I(N__6430));
    LocalMux I__888 (
            .O(N__6430),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_7 ));
    CascadeMux I__887 (
            .O(N__6427),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_ ));
    InMux I__886 (
            .O(N__6424),
            .I(N__6421));
    LocalMux I__885 (
            .O(N__6421),
            .I(N__6418));
    Odrv4 I__884 (
            .O(N__6418),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_7 ));
    InMux I__883 (
            .O(N__6415),
            .I(N__6404));
    InMux I__882 (
            .O(N__6414),
            .I(N__6401));
    InMux I__881 (
            .O(N__6413),
            .I(N__6393));
    InMux I__880 (
            .O(N__6412),
            .I(N__6393));
    InMux I__879 (
            .O(N__6411),
            .I(N__6393));
    InMux I__878 (
            .O(N__6410),
            .I(N__6389));
    InMux I__877 (
            .O(N__6409),
            .I(N__6386));
    InMux I__876 (
            .O(N__6408),
            .I(N__6381));
    InMux I__875 (
            .O(N__6407),
            .I(N__6381));
    LocalMux I__874 (
            .O(N__6404),
            .I(N__6378));
    LocalMux I__873 (
            .O(N__6401),
            .I(N__6375));
    InMux I__872 (
            .O(N__6400),
            .I(N__6372));
    LocalMux I__871 (
            .O(N__6393),
            .I(N__6369));
    InMux I__870 (
            .O(N__6392),
            .I(N__6366));
    LocalMux I__869 (
            .O(N__6389),
            .I(\DUT.fifo_tx_inst.N_33 ));
    LocalMux I__868 (
            .O(N__6386),
            .I(\DUT.fifo_tx_inst.N_33 ));
    LocalMux I__867 (
            .O(N__6381),
            .I(\DUT.fifo_tx_inst.N_33 ));
    Odrv4 I__866 (
            .O(N__6378),
            .I(\DUT.fifo_tx_inst.N_33 ));
    Odrv12 I__865 (
            .O(N__6375),
            .I(\DUT.fifo_tx_inst.N_33 ));
    LocalMux I__864 (
            .O(N__6372),
            .I(\DUT.fifo_tx_inst.N_33 ));
    Odrv4 I__863 (
            .O(N__6369),
            .I(\DUT.fifo_tx_inst.N_33 ));
    LocalMux I__862 (
            .O(N__6366),
            .I(\DUT.fifo_tx_inst.N_33 ));
    CEMux I__861 (
            .O(N__6349),
            .I(N__6346));
    LocalMux I__860 (
            .O(N__6346),
            .I(\DUT.fifo_tx_inst.N_41 ));
    InMux I__859 (
            .O(N__6343),
            .I(N__6340));
    LocalMux I__858 (
            .O(N__6340),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_4 ));
    InMux I__857 (
            .O(N__6337),
            .I(N__6334));
    LocalMux I__856 (
            .O(N__6334),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_4 ));
    InMux I__855 (
            .O(N__6331),
            .I(N__6328));
    LocalMux I__854 (
            .O(N__6328),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_2 ));
    InMux I__853 (
            .O(N__6325),
            .I(N__6322));
    LocalMux I__852 (
            .O(N__6322),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_2 ));
    CascadeMux I__851 (
            .O(N__6319),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_ ));
    InMux I__850 (
            .O(N__6316),
            .I(N__6313));
    LocalMux I__849 (
            .O(N__6313),
            .I(N__6310));
    Odrv4 I__848 (
            .O(N__6310),
            .I(\DUT.fifo_tx_inst.rFifoData_ram2_2 ));
    CascadeMux I__847 (
            .O(N__6307),
            .I(\DUT.rFifoDatarx_2_cascade_ ));
    InMux I__846 (
            .O(N__6304),
            .I(N__6300));
    InMux I__845 (
            .O(N__6303),
            .I(N__6297));
    LocalMux I__844 (
            .O(N__6300),
            .I(\DUT.fifo_tx_inst.rFifoDataro_1 ));
    LocalMux I__843 (
            .O(N__6297),
            .I(\DUT.fifo_tx_inst.rFifoDataro_1 ));
    InMux I__842 (
            .O(N__6292),
            .I(N__6288));
    InMux I__841 (
            .O(N__6291),
            .I(N__6285));
    LocalMux I__840 (
            .O(N__6288),
            .I(\DUT.fifo_tx_inst.rFifoDataro_0 ));
    LocalMux I__839 (
            .O(N__6285),
            .I(\DUT.fifo_tx_inst.rFifoDataro_0 ));
    CascadeMux I__838 (
            .O(N__6280),
            .I(\DUT.fifo_tx_inst.rFifoDataror_1_0_cascade_ ));
    InMux I__837 (
            .O(N__6277),
            .I(N__6274));
    LocalMux I__836 (
            .O(N__6274),
            .I(N__6271));
    Odrv4 I__835 (
            .O(N__6271),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_0 ));
    InMux I__834 (
            .O(N__6268),
            .I(N__6265));
    LocalMux I__833 (
            .O(N__6265),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_0 ));
    CascadeMux I__832 (
            .O(N__6262),
            .I(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ));
    CascadeMux I__831 (
            .O(N__6259),
            .I(\DUT.fifo_tx_inst.un1_i11_2_i_cascade_ ));
    InMux I__830 (
            .O(N__6256),
            .I(N__6253));
    LocalMux I__829 (
            .O(N__6253),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_1 ));
    CascadeMux I__828 (
            .O(N__6250),
            .I(N__6247));
    InMux I__827 (
            .O(N__6247),
            .I(N__6244));
    LocalMux I__826 (
            .O(N__6244),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_1 ));
    InMux I__825 (
            .O(N__6241),
            .I(N__6238));
    LocalMux I__824 (
            .O(N__6238),
            .I(\DUT.fifo_tx_inst.rFifoData_ram1_3 ));
    InMux I__823 (
            .O(N__6235),
            .I(N__6232));
    LocalMux I__822 (
            .O(N__6232),
            .I(\DUT.fifo_tx_inst.rFifoData_ram0_3 ));
    InMux I__821 (
            .O(N__6229),
            .I(N__6226));
    LocalMux I__820 (
            .O(N__6226),
            .I(\DUT.fifo_tx_inst.CO0 ));
    CascadeMux I__819 (
            .O(N__6223),
            .I(\DUT.fifo_tx_inst.CO0_cascade_ ));
    InMux I__818 (
            .O(N__6220),
            .I(N__6217));
    LocalMux I__817 (
            .O(N__6217),
            .I(\DUT.fifo_tx_inst.un1_i11_2_i ));
    IoInMux I__816 (
            .O(N__6214),
            .I(N__6211));
    LocalMux I__815 (
            .O(N__6211),
            .I(N__6208));
    Span4Mux_s1_v I__814 (
            .O(N__6208),
            .I(N__6205));
    Span4Mux_v I__813 (
            .O(N__6205),
            .I(N__6201));
    InMux I__812 (
            .O(N__6204),
            .I(N__6198));
    Span4Mux_v I__811 (
            .O(N__6201),
            .I(N__6193));
    LocalMux I__810 (
            .O(N__6198),
            .I(N__6193));
    Span4Mux_v I__809 (
            .O(N__6193),
            .I(N__6189));
    InMux I__808 (
            .O(N__6192),
            .I(N__6186));
    Odrv4 I__807 (
            .O(N__6189),
            .I(oTx_n_c));
    LocalMux I__806 (
            .O(N__6186),
            .I(oTx_n_c));
    IoInMux I__805 (
            .O(N__6181),
            .I(N__6178));
    LocalMux I__804 (
            .O(N__6178),
            .I(N__6175));
    Span4Mux_s3_v I__803 (
            .O(N__6175),
            .I(N__6172));
    Span4Mux_h I__802 (
            .O(N__6172),
            .I(N__6169));
    Sp12to4 I__801 (
            .O(N__6169),
            .I(N__6166));
    Span12Mux_v I__800 (
            .O(N__6166),
            .I(N__6162));
    InMux I__799 (
            .O(N__6165),
            .I(N__6159));
    Odrv12 I__798 (
            .O(N__6162),
            .I(P1A2_c));
    LocalMux I__797 (
            .O(N__6159),
            .I(P1A2_c));
    InMux I__796 (
            .O(N__6154),
            .I(N__6150));
    InMux I__795 (
            .O(N__6153),
            .I(N__6147));
    LocalMux I__794 (
            .O(N__6150),
            .I(N__6139));
    LocalMux I__793 (
            .O(N__6147),
            .I(N__6139));
    InMux I__792 (
            .O(N__6146),
            .I(N__6132));
    InMux I__791 (
            .O(N__6145),
            .I(N__6132));
    InMux I__790 (
            .O(N__6144),
            .I(N__6132));
    Odrv4 I__789 (
            .O(N__6139),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_0 ));
    LocalMux I__788 (
            .O(N__6132),
            .I(\DUT.fifo_tx_inst.rFifoCountZ0Z_0 ));
    CascadeMux I__787 (
            .O(N__6127),
            .I(N__6124));
    InMux I__786 (
            .O(N__6124),
            .I(N__6121));
    LocalMux I__785 (
            .O(N__6121),
            .I(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0 ));
    InMux I__784 (
            .O(N__6118),
            .I(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0 ));
    CascadeMux I__783 (
            .O(N__6115),
            .I(N__6111));
    CascadeMux I__782 (
            .O(N__6114),
            .I(N__6108));
    InMux I__781 (
            .O(N__6111),
            .I(N__6105));
    InMux I__780 (
            .O(N__6108),
            .I(N__6102));
    LocalMux I__779 (
            .O(N__6105),
            .I(\DUT.fifo_tx_inst.N_35 ));
    LocalMux I__778 (
            .O(N__6102),
            .I(\DUT.fifo_tx_inst.N_35 ));
    InMux I__777 (
            .O(N__6097),
            .I(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1 ));
    InMux I__776 (
            .O(N__6094),
            .I(N__6088));
    InMux I__775 (
            .O(N__6093),
            .I(N__6088));
    LocalMux I__774 (
            .O(N__6088),
            .I(\DUT.fifo_tx_inst.rFifoDataro_3 ));
    InMux I__773 (
            .O(N__6085),
            .I(N__6079));
    InMux I__772 (
            .O(N__6084),
            .I(N__6079));
    LocalMux I__771 (
            .O(N__6079),
            .I(\DUT.fifo_tx_inst.rFifoDataro_2 ));
    InMux I__770 (
            .O(N__6076),
            .I(N__6073));
    LocalMux I__769 (
            .O(N__6073),
            .I(\DUT.fifo_rx_inst.rTxByte_42_0 ));
    CascadeMux I__768 (
            .O(N__6070),
            .I(\DUT.fifo_rx_inst.rTxByte_42_1_cascade_ ));
    InMux I__767 (
            .O(N__6067),
            .I(N__6063));
    CascadeMux I__766 (
            .O(N__6066),
            .I(N__6059));
    LocalMux I__765 (
            .O(N__6063),
            .I(N__6055));
    InMux I__764 (
            .O(N__6062),
            .I(N__6050));
    InMux I__763 (
            .O(N__6059),
            .I(N__6050));
    InMux I__762 (
            .O(N__6058),
            .I(N__6047));
    Odrv4 I__761 (
            .O(N__6055),
            .I(wRxBufferEmpty_i_0));
    LocalMux I__760 (
            .O(N__6050),
            .I(wRxBufferEmpty_i_0));
    LocalMux I__759 (
            .O(N__6047),
            .I(wRxBufferEmpty_i_0));
    SRMux I__758 (
            .O(N__6040),
            .I(N__6037));
    LocalMux I__757 (
            .O(N__6037),
            .I(N__6033));
    SRMux I__756 (
            .O(N__6036),
            .I(N__6030));
    Span4Mux_v I__755 (
            .O(N__6033),
            .I(N__6025));
    LocalMux I__754 (
            .O(N__6030),
            .I(N__6025));
    Sp12to4 I__753 (
            .O(N__6025),
            .I(N__6021));
    InMux I__752 (
            .O(N__6024),
            .I(N__6018));
    Odrv12 I__751 (
            .O(N__6021),
            .I(rFifoDatarff_0_RNIHJV05));
    LocalMux I__750 (
            .O(N__6018),
            .I(rFifoDatarff_0_RNIHJV05));
    CascadeMux I__749 (
            .O(N__6013),
            .I(N__6004));
    InMux I__748 (
            .O(N__6012),
            .I(N__5976));
    InMux I__747 (
            .O(N__6011),
            .I(N__5976));
    InMux I__746 (
            .O(N__6010),
            .I(N__5976));
    InMux I__745 (
            .O(N__6009),
            .I(N__5976));
    InMux I__744 (
            .O(N__6008),
            .I(N__5976));
    InMux I__743 (
            .O(N__6007),
            .I(N__5976));
    InMux I__742 (
            .O(N__6004),
            .I(N__5976));
    InMux I__741 (
            .O(N__6003),
            .I(N__5976));
    CascadeMux I__740 (
            .O(N__6002),
            .I(N__5971));
    CascadeMux I__739 (
            .O(N__6001),
            .I(N__5968));
    InMux I__738 (
            .O(N__6000),
            .I(N__5951));
    InMux I__737 (
            .O(N__5999),
            .I(N__5951));
    InMux I__736 (
            .O(N__5998),
            .I(N__5951));
    InMux I__735 (
            .O(N__5997),
            .I(N__5951));
    InMux I__734 (
            .O(N__5996),
            .I(N__5951));
    InMux I__733 (
            .O(N__5995),
            .I(N__5951));
    InMux I__732 (
            .O(N__5994),
            .I(N__5951));
    InMux I__731 (
            .O(N__5993),
            .I(N__5951));
    LocalMux I__730 (
            .O(N__5976),
            .I(N__5948));
    InMux I__729 (
            .O(N__5975),
            .I(N__5941));
    InMux I__728 (
            .O(N__5974),
            .I(N__5941));
    InMux I__727 (
            .O(N__5971),
            .I(N__5941));
    InMux I__726 (
            .O(N__5968),
            .I(N__5938));
    LocalMux I__725 (
            .O(N__5951),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    Odrv4 I__724 (
            .O(N__5948),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__723 (
            .O(N__5941),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    LocalMux I__722 (
            .O(N__5938),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ));
    InMux I__721 (
            .O(N__5929),
            .I(N__5926));
    LocalMux I__720 (
            .O(N__5926),
            .I(\DUT.fifo_rx_inst.rReadPtr_RNI4NC92Z0Z_0 ));
    CascadeMux I__719 (
            .O(N__5923),
            .I(N__5920));
    InMux I__718 (
            .O(N__5920),
            .I(N__5911));
    InMux I__717 (
            .O(N__5919),
            .I(N__5911));
    InMux I__716 (
            .O(N__5918),
            .I(N__5911));
    LocalMux I__715 (
            .O(N__5911),
            .I(\DUT.fifo_rx_inst.N_73 ));
    CascadeMux I__714 (
            .O(N__5908),
            .I(\DUT.fifo_rx_inst.rReadPtr_RNI4NC92Z0Z_0_cascade_ ));
    InMux I__713 (
            .O(N__5905),
            .I(N__5889));
    InMux I__712 (
            .O(N__5904),
            .I(N__5889));
    InMux I__711 (
            .O(N__5903),
            .I(N__5889));
    InMux I__710 (
            .O(N__5902),
            .I(N__5889));
    InMux I__709 (
            .O(N__5901),
            .I(N__5875));
    InMux I__708 (
            .O(N__5900),
            .I(N__5875));
    InMux I__707 (
            .O(N__5899),
            .I(N__5875));
    InMux I__706 (
            .O(N__5898),
            .I(N__5875));
    LocalMux I__705 (
            .O(N__5889),
            .I(N__5872));
    InMux I__704 (
            .O(N__5888),
            .I(N__5863));
    InMux I__703 (
            .O(N__5887),
            .I(N__5863));
    InMux I__702 (
            .O(N__5886),
            .I(N__5863));
    InMux I__701 (
            .O(N__5885),
            .I(N__5863));
    InMux I__700 (
            .O(N__5884),
            .I(N__5860));
    LocalMux I__699 (
            .O(N__5875),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    Odrv4 I__698 (
            .O(N__5872),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__697 (
            .O(N__5863),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    LocalMux I__696 (
            .O(N__5860),
            .I(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ));
    CascadeMux I__695 (
            .O(N__5851),
            .I(\DUT.uart_inst0.recv_state_srsts_1_0_6_cascade_ ));
    InMux I__694 (
            .O(N__5848),
            .I(N__5844));
    InMux I__693 (
            .O(N__5847),
            .I(N__5841));
    LocalMux I__692 (
            .O(N__5844),
            .I(\DUT.fifo_rx_inst.un1_rFifoCount16_0_0 ));
    LocalMux I__691 (
            .O(N__5841),
            .I(\DUT.fifo_rx_inst.un1_rFifoCount16_0_0 ));
    InMux I__690 (
            .O(N__5836),
            .I(N__5833));
    LocalMux I__689 (
            .O(N__5833),
            .I(N__5828));
    CascadeMux I__688 (
            .O(N__5832),
            .I(N__5825));
    InMux I__687 (
            .O(N__5831),
            .I(N__5820));
    Span4Mux_h I__686 (
            .O(N__5828),
            .I(N__5817));
    InMux I__685 (
            .O(N__5825),
            .I(N__5814));
    InMux I__684 (
            .O(N__5824),
            .I(N__5809));
    InMux I__683 (
            .O(N__5823),
            .I(N__5809));
    LocalMux I__682 (
            .O(N__5820),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_0 ));
    Odrv4 I__681 (
            .O(N__5817),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_0 ));
    LocalMux I__680 (
            .O(N__5814),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_0 ));
    LocalMux I__679 (
            .O(N__5809),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_0 ));
    CEMux I__678 (
            .O(N__5800),
            .I(N__5797));
    LocalMux I__677 (
            .O(N__5797),
            .I(N__5794));
    Sp12to4 I__676 (
            .O(N__5794),
            .I(N__5790));
    InMux I__675 (
            .O(N__5793),
            .I(N__5787));
    Odrv12 I__674 (
            .O(N__5790),
            .I(\DUT.fifo_rx_inst.rFifoData_awe0 ));
    LocalMux I__673 (
            .O(N__5787),
            .I(\DUT.fifo_rx_inst.rFifoData_awe0 ));
    InMux I__672 (
            .O(N__5782),
            .I(N__5778));
    InMux I__671 (
            .O(N__5781),
            .I(N__5775));
    LocalMux I__670 (
            .O(N__5778),
            .I(\DUT.fifo_rx_inst.rFifoDataro_0 ));
    LocalMux I__669 (
            .O(N__5775),
            .I(\DUT.fifo_rx_inst.rFifoDataro_0 ));
    InMux I__668 (
            .O(N__5770),
            .I(N__5767));
    LocalMux I__667 (
            .O(N__5767),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_1 ));
    InMux I__666 (
            .O(N__5764),
            .I(N__5761));
    LocalMux I__665 (
            .O(N__5761),
            .I(N__5758));
    Odrv4 I__664 (
            .O(N__5758),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_1 ));
    CascadeMux I__663 (
            .O(N__5755),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1_cascade_ ));
    InMux I__662 (
            .O(N__5752),
            .I(N__5749));
    LocalMux I__661 (
            .O(N__5749),
            .I(N__5746));
    Odrv4 I__660 (
            .O(N__5746),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_1 ));
    InMux I__659 (
            .O(N__5743),
            .I(N__5740));
    LocalMux I__658 (
            .O(N__5740),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_7 ));
    InMux I__657 (
            .O(N__5737),
            .I(N__5734));
    LocalMux I__656 (
            .O(N__5734),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7 ));
    InMux I__655 (
            .O(N__5731),
            .I(N__5728));
    LocalMux I__654 (
            .O(N__5728),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_0 ));
    InMux I__653 (
            .O(N__5725),
            .I(N__5722));
    LocalMux I__652 (
            .O(N__5722),
            .I(N__5719));
    Odrv4 I__651 (
            .O(N__5719),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_0 ));
    InMux I__650 (
            .O(N__5716),
            .I(N__5713));
    LocalMux I__649 (
            .O(N__5713),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_0 ));
    CascadeMux I__648 (
            .O(N__5710),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ));
    CEMux I__647 (
            .O(N__5707),
            .I(N__5703));
    CEMux I__646 (
            .O(N__5706),
            .I(N__5700));
    LocalMux I__645 (
            .O(N__5703),
            .I(N__5697));
    LocalMux I__644 (
            .O(N__5700),
            .I(N__5694));
    Odrv4 I__643 (
            .O(N__5697),
            .I(wRxBufferEmpty_i_0_0));
    Odrv4 I__642 (
            .O(N__5694),
            .I(wRxBufferEmpty_i_0_0));
    InMux I__641 (
            .O(N__5689),
            .I(N__5685));
    InMux I__640 (
            .O(N__5688),
            .I(N__5682));
    LocalMux I__639 (
            .O(N__5685),
            .I(\DUT.fifo_rx_inst.rFifoDataro_1 ));
    LocalMux I__638 (
            .O(N__5682),
            .I(\DUT.fifo_rx_inst.rFifoDataro_1 ));
    CascadeMux I__637 (
            .O(N__5677),
            .I(G_143_cascade_));
    CascadeMux I__636 (
            .O(N__5674),
            .I(\fifo_inst.ftdi_input_inst.SUMZ0Z_2_cascade_ ));
    CEMux I__635 (
            .O(N__5671),
            .I(N__5667));
    CEMux I__634 (
            .O(N__5670),
            .I(N__5664));
    LocalMux I__633 (
            .O(N__5667),
            .I(N__5660));
    LocalMux I__632 (
            .O(N__5664),
            .I(N__5657));
    CEMux I__631 (
            .O(N__5663),
            .I(N__5654));
    Span4Mux_v I__630 (
            .O(N__5660),
            .I(N__5651));
    Span4Mux_h I__629 (
            .O(N__5657),
            .I(N__5647));
    LocalMux I__628 (
            .O(N__5654),
            .I(N__5642));
    Span4Mux_h I__627 (
            .O(N__5651),
            .I(N__5642));
    InMux I__626 (
            .O(N__5650),
            .I(N__5639));
    Odrv4 I__625 (
            .O(N__5647),
            .I(\DUT.fifo_rx_inst.N_86 ));
    Odrv4 I__624 (
            .O(N__5642),
            .I(\DUT.fifo_rx_inst.N_86 ));
    LocalMux I__623 (
            .O(N__5639),
            .I(\DUT.fifo_rx_inst.N_86 ));
    InMux I__622 (
            .O(N__5632),
            .I(N__5629));
    LocalMux I__621 (
            .O(N__5629),
            .I(N__5626));
    Odrv4 I__620 (
            .O(N__5626),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_7 ));
    CascadeMux I__619 (
            .O(N__5623),
            .I(N__5620));
    InMux I__618 (
            .O(N__5620),
            .I(N__5617));
    LocalMux I__617 (
            .O(N__5617),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_7 ));
    InMux I__616 (
            .O(N__5614),
            .I(N__5611));
    LocalMux I__615 (
            .O(N__5611),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_2 ));
    InMux I__614 (
            .O(N__5608),
            .I(N__5605));
    LocalMux I__613 (
            .O(N__5605),
            .I(N__5602));
    Odrv12 I__612 (
            .O(N__5602),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_2 ));
    CascadeMux I__611 (
            .O(N__5599),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2_cascade_ ));
    InMux I__610 (
            .O(N__5596),
            .I(N__5593));
    LocalMux I__609 (
            .O(N__5593),
            .I(N__5590));
    Odrv4 I__608 (
            .O(N__5590),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_2 ));
    CascadeMux I__607 (
            .O(N__5587),
            .I(wRxBufferEmpty_i_0_cascade_));
    InMux I__606 (
            .O(N__5584),
            .I(N__5581));
    LocalMux I__605 (
            .O(N__5581),
            .I(\DUT.fifo_rx_inst.un1_rFifoCount16_0_i_0 ));
    CascadeMux I__604 (
            .O(N__5578),
            .I(N__5575));
    InMux I__603 (
            .O(N__5575),
            .I(N__5572));
    LocalMux I__602 (
            .O(N__5572),
            .I(\DUT.fifo_rx_inst.rFifoCount_RNIK3G92Z0Z_1 ));
    InMux I__601 (
            .O(N__5569),
            .I(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0 ));
    InMux I__600 (
            .O(N__5566),
            .I(N__5563));
    LocalMux I__599 (
            .O(N__5563),
            .I(\DUT.fifo_rx_inst.un1_rFifoCount_1_axb_2 ));
    InMux I__598 (
            .O(N__5560),
            .I(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1 ));
    InMux I__597 (
            .O(N__5557),
            .I(N__5552));
    InMux I__596 (
            .O(N__5556),
            .I(N__5549));
    InMux I__595 (
            .O(N__5555),
            .I(N__5542));
    LocalMux I__594 (
            .O(N__5552),
            .I(N__5537));
    LocalMux I__593 (
            .O(N__5549),
            .I(N__5537));
    InMux I__592 (
            .O(N__5548),
            .I(N__5528));
    InMux I__591 (
            .O(N__5547),
            .I(N__5528));
    InMux I__590 (
            .O(N__5546),
            .I(N__5528));
    InMux I__589 (
            .O(N__5545),
            .I(N__5528));
    LocalMux I__588 (
            .O(N__5542),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ));
    Odrv4 I__587 (
            .O(N__5537),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ));
    LocalMux I__586 (
            .O(N__5528),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ));
    CascadeMux I__585 (
            .O(N__5521),
            .I(N__5515));
    InMux I__584 (
            .O(N__5520),
            .I(N__5511));
    InMux I__583 (
            .O(N__5519),
            .I(N__5508));
    InMux I__582 (
            .O(N__5518),
            .I(N__5501));
    InMux I__581 (
            .O(N__5515),
            .I(N__5501));
    InMux I__580 (
            .O(N__5514),
            .I(N__5501));
    LocalMux I__579 (
            .O(N__5511),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_1 ));
    LocalMux I__578 (
            .O(N__5508),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_1 ));
    LocalMux I__577 (
            .O(N__5501),
            .I(\DUT.fifo_rx_inst.rFifoCountZ0Z_1 ));
    CascadeMux I__576 (
            .O(N__5494),
            .I(\DUT.fifo_tx_inst.N_35_cascade_ ));
    InMux I__575 (
            .O(N__5491),
            .I(N__5485));
    InMux I__574 (
            .O(N__5490),
            .I(N__5485));
    LocalMux I__573 (
            .O(N__5485),
            .I(\DUT.fifo_rx_inst.rFifoDataro_3 ));
    InMux I__572 (
            .O(N__5482),
            .I(N__5476));
    InMux I__571 (
            .O(N__5481),
            .I(N__5476));
    LocalMux I__570 (
            .O(N__5476),
            .I(\DUT.fifo_rx_inst.rFifoDataro_2 ));
    InMux I__569 (
            .O(N__5473),
            .I(N__5465));
    InMux I__568 (
            .O(N__5472),
            .I(N__5465));
    InMux I__567 (
            .O(N__5471),
            .I(N__5460));
    InMux I__566 (
            .O(N__5470),
            .I(N__5460));
    LocalMux I__565 (
            .O(N__5465),
            .I(\DUT.fifo_rx_inst.N_42 ));
    LocalMux I__564 (
            .O(N__5460),
            .I(\DUT.fifo_rx_inst.N_42 ));
    CascadeMux I__563 (
            .O(N__5455),
            .I(N__5447));
    InMux I__562 (
            .O(N__5454),
            .I(N__5440));
    InMux I__561 (
            .O(N__5453),
            .I(N__5440));
    InMux I__560 (
            .O(N__5452),
            .I(N__5440));
    InMux I__559 (
            .O(N__5451),
            .I(N__5433));
    InMux I__558 (
            .O(N__5450),
            .I(N__5433));
    InMux I__557 (
            .O(N__5447),
            .I(N__5433));
    LocalMux I__556 (
            .O(N__5440),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_0 ));
    LocalMux I__555 (
            .O(N__5433),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_0 ));
    CascadeMux I__554 (
            .O(N__5428),
            .I(\DUT.fifo_rx_inst.N_42_cascade_ ));
    CascadeMux I__553 (
            .O(N__5425),
            .I(N__5419));
    InMux I__552 (
            .O(N__5424),
            .I(N__5411));
    InMux I__551 (
            .O(N__5423),
            .I(N__5411));
    InMux I__550 (
            .O(N__5422),
            .I(N__5411));
    InMux I__549 (
            .O(N__5419),
            .I(N__5406));
    InMux I__548 (
            .O(N__5418),
            .I(N__5406));
    LocalMux I__547 (
            .O(N__5411),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_1 ));
    LocalMux I__546 (
            .O(N__5406),
            .I(\DUT.fifo_rx_inst.rWritePtrZ0Z_1 ));
    CascadeMux I__545 (
            .O(N__5401),
            .I(\DUT.fifo_rx_inst.rFifoData_awe1_cascade_ ));
    CascadeMux I__544 (
            .O(N__5398),
            .I(N__5395));
    InMux I__543 (
            .O(N__5395),
            .I(N__5392));
    LocalMux I__542 (
            .O(N__5392),
            .I(\DUT.fifo_tx_inst.un1_i11_i ));
    CascadeMux I__541 (
            .O(N__5389),
            .I(\DUT.fifo_tx_inst.un1_i11_i_cascade_ ));
    InMux I__540 (
            .O(N__5386),
            .I(N__5383));
    LocalMux I__539 (
            .O(N__5383),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_5 ));
    InMux I__538 (
            .O(N__5380),
            .I(N__5377));
    LocalMux I__537 (
            .O(N__5377),
            .I(N__5374));
    Odrv4 I__536 (
            .O(N__5374),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_6 ));
    InMux I__535 (
            .O(N__5371),
            .I(N__5368));
    LocalMux I__534 (
            .O(N__5368),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_6 ));
    CascadeMux I__533 (
            .O(N__5365),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6_cascade_ ));
    InMux I__532 (
            .O(N__5362),
            .I(N__5359));
    LocalMux I__531 (
            .O(N__5359),
            .I(N__5356));
    Odrv4 I__530 (
            .O(N__5356),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_6 ));
    InMux I__529 (
            .O(N__5353),
            .I(N__5350));
    LocalMux I__528 (
            .O(N__5350),
            .I(N__5347));
    Odrv4 I__527 (
            .O(N__5347),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_4 ));
    InMux I__526 (
            .O(N__5344),
            .I(N__5341));
    LocalMux I__525 (
            .O(N__5341),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4 ));
    InMux I__524 (
            .O(N__5338),
            .I(N__5335));
    LocalMux I__523 (
            .O(N__5335),
            .I(N__5332));
    Odrv4 I__522 (
            .O(N__5332),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_3 ));
    InMux I__521 (
            .O(N__5329),
            .I(N__5326));
    LocalMux I__520 (
            .O(N__5326),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_3 ));
    InMux I__519 (
            .O(N__5323),
            .I(N__5320));
    LocalMux I__518 (
            .O(N__5320),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_3 ));
    CascadeMux I__517 (
            .O(N__5317),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ));
    CEMux I__516 (
            .O(N__5314),
            .I(N__5311));
    LocalMux I__515 (
            .O(N__5311),
            .I(N__5308));
    Span4Mux_v I__514 (
            .O(N__5308),
            .I(N__5305));
    Odrv4 I__513 (
            .O(N__5305),
            .I(\DUT.fifo_rx_inst.rFifoData_awe2 ));
    CascadeMux I__512 (
            .O(N__5302),
            .I(\DUT.fifo_rx_inst.rFifoData_awe2_cascade_ ));
    InMux I__511 (
            .O(N__5299),
            .I(N__5296));
    LocalMux I__510 (
            .O(N__5296),
            .I(\DUT.fifo_rx_inst.rFifoData_ram2_4 ));
    CascadeMux I__509 (
            .O(N__5293),
            .I(N__5290));
    InMux I__508 (
            .O(N__5290),
            .I(N__5287));
    LocalMux I__507 (
            .O(N__5287),
            .I(N__5284));
    Odrv4 I__506 (
            .O(N__5284),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_4 ));
    InMux I__505 (
            .O(N__5281),
            .I(N__5278));
    LocalMux I__504 (
            .O(N__5278),
            .I(N__5275));
    Odrv4 I__503 (
            .O(N__5275),
            .I(\DUT.fifo_rx_inst.rFifoData_ram0_5 ));
    InMux I__502 (
            .O(N__5272),
            .I(N__5269));
    LocalMux I__501 (
            .O(N__5269),
            .I(\DUT.fifo_rx_inst.rFifoData_ram3_5 ));
    CascadeMux I__500 (
            .O(N__5266),
            .I(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ));
    CascadeMux I__499 (
            .O(N__5263),
            .I(\DUT.fifo_rx_inst.N_86_cascade_ ));
    InMux I__498 (
            .O(N__5260),
            .I(N__5257));
    LocalMux I__497 (
            .O(N__5257),
            .I(\DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1 ));
    CascadeMux I__496 (
            .O(N__5254),
            .I(\DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1_cascade_ ));
    IoInMux I__495 (
            .O(N__5251),
            .I(N__5247));
    IoInMux I__494 (
            .O(N__5250),
            .I(N__5244));
    LocalMux I__493 (
            .O(N__5247),
            .I(N__5239));
    LocalMux I__492 (
            .O(N__5244),
            .I(N__5236));
    IoInMux I__491 (
            .O(N__5243),
            .I(N__5233));
    IoInMux I__490 (
            .O(N__5242),
            .I(N__5230));
    IoSpan4Mux I__489 (
            .O(N__5239),
            .I(N__5220));
    IoSpan4Mux I__488 (
            .O(N__5236),
            .I(N__5220));
    LocalMux I__487 (
            .O(N__5233),
            .I(N__5220));
    LocalMux I__486 (
            .O(N__5230),
            .I(N__5220));
    IoInMux I__485 (
            .O(N__5229),
            .I(N__5217));
    IoSpan4Mux I__484 (
            .O(N__5220),
            .I(N__5209));
    LocalMux I__483 (
            .O(N__5217),
            .I(N__5209));
    IoInMux I__482 (
            .O(N__5216),
            .I(N__5206));
    IoInMux I__481 (
            .O(N__5215),
            .I(N__5203));
    IoInMux I__480 (
            .O(N__5214),
            .I(N__5200));
    IoSpan4Mux I__479 (
            .O(N__5209),
            .I(N__5197));
    LocalMux I__478 (
            .O(N__5206),
            .I(N__5194));
    LocalMux I__477 (
            .O(N__5203),
            .I(N__5189));
    LocalMux I__476 (
            .O(N__5200),
            .I(N__5189));
    Span4Mux_s2_v I__475 (
            .O(N__5197),
            .I(N__5184));
    Span4Mux_s2_v I__474 (
            .O(N__5194),
            .I(N__5184));
    IoSpan4Mux I__473 (
            .O(N__5189),
            .I(N__5181));
    Span4Mux_v I__472 (
            .O(N__5184),
            .I(N__5178));
    Sp12to4 I__471 (
            .O(N__5181),
            .I(N__5175));
    Span4Mux_v I__470 (
            .O(N__5178),
            .I(N__5172));
    Span12Mux_v I__469 (
            .O(N__5175),
            .I(N__5169));
    Span4Mux_v I__468 (
            .O(N__5172),
            .I(N__5166));
    Odrv12 I__467 (
            .O(N__5169),
            .I(oTx_n_c_i));
    Odrv4 I__466 (
            .O(N__5166),
            .I(oTx_n_c_i));
    IoInMux I__465 (
            .O(N__5161),
            .I(N__5158));
    LocalMux I__464 (
            .O(N__5158),
            .I(N__5155));
    Span4Mux_s3_v I__463 (
            .O(N__5155),
            .I(N__5152));
    Span4Mux_v I__462 (
            .O(N__5152),
            .I(N__5149));
    Span4Mux_h I__461 (
            .O(N__5149),
            .I(N__5146));
    Odrv4 I__460 (
            .O(N__5146),
            .I(wRamRdData_1));
    InMux I__459 (
            .O(N__5143),
            .I(N__5140));
    LocalMux I__458 (
            .O(N__5140),
            .I(\PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO ));
    IoInMux I__457 (
            .O(N__5137),
            .I(N__5134));
    LocalMux I__456 (
            .O(N__5134),
            .I(N__5131));
    Span12Mux_s9_v I__455 (
            .O(N__5131),
            .I(N__5128));
    Span12Mux_v I__454 (
            .O(N__5128),
            .I(N__5125));
    Odrv12 I__453 (
            .O(N__5125),
            .I(BTN_N_c));
    IoInMux I__452 (
            .O(N__5122),
            .I(N__5119));
    LocalMux I__451 (
            .O(N__5119),
            .I(N__5116));
    Sp12to4 I__450 (
            .O(N__5116),
            .I(N__5113));
    Span12Mux_v I__449 (
            .O(N__5113),
            .I(N__5110));
    Odrv12 I__448 (
            .O(N__5110),
            .I(wRamRdData_7));
    IoInMux I__447 (
            .O(N__5107),
            .I(N__5104));
    LocalMux I__446 (
            .O(N__5104),
            .I(N__5101));
    Span4Mux_s1_v I__445 (
            .O(N__5101),
            .I(N__5098));
    Span4Mux_v I__444 (
            .O(N__5098),
            .I(N__5095));
    Span4Mux_v I__443 (
            .O(N__5095),
            .I(N__5092));
    Span4Mux_h I__442 (
            .O(N__5092),
            .I(N__5089));
    Odrv4 I__441 (
            .O(N__5089),
            .I(wRamRdData_0));
    IoInMux I__440 (
            .O(N__5086),
            .I(N__5083));
    LocalMux I__439 (
            .O(N__5083),
            .I(N__5080));
    Span12Mux_s3_v I__438 (
            .O(N__5080),
            .I(N__5077));
    Odrv12 I__437 (
            .O(N__5077),
            .I(wRamRdData_4));
    IoInMux I__436 (
            .O(N__5074),
            .I(N__5071));
    LocalMux I__435 (
            .O(N__5071),
            .I(N__5068));
    Span12Mux_s10_v I__434 (
            .O(N__5068),
            .I(N__5065));
    Odrv12 I__433 (
            .O(N__5065),
            .I(wRamRdData_6));
    IoInMux I__432 (
            .O(N__5062),
            .I(N__5059));
    LocalMux I__431 (
            .O(N__5059),
            .I(N__5056));
    Span4Mux_s1_v I__430 (
            .O(N__5056),
            .I(N__5053));
    Span4Mux_v I__429 (
            .O(N__5053),
            .I(N__5050));
    Span4Mux_v I__428 (
            .O(N__5050),
            .I(N__5047));
    Odrv4 I__427 (
            .O(N__5047),
            .I(wRamRdData_2));
    IoInMux I__426 (
            .O(N__5044),
            .I(N__5041));
    LocalMux I__425 (
            .O(N__5041),
            .I(N__5038));
    Span4Mux_s1_v I__424 (
            .O(N__5038),
            .I(N__5035));
    Span4Mux_v I__423 (
            .O(N__5035),
            .I(N__5032));
    Span4Mux_v I__422 (
            .O(N__5032),
            .I(N__5029));
    Odrv4 I__421 (
            .O(N__5029),
            .I(wRamRdData_3));
    IoInMux I__420 (
            .O(N__5026),
            .I(N__5023));
    LocalMux I__419 (
            .O(N__5023),
            .I(N__5020));
    Span12Mux_s8_v I__418 (
            .O(N__5020),
            .I(N__5017));
    Odrv12 I__417 (
            .O(N__5017),
            .I(wRamRdData_5));
    defparam IN_MUX_bfv_18_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_19_0_));
    defparam IN_MUX_bfv_18_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_20_0_ (
            .carryinitin(\DUT.uart_inst0.tx_clk_divider_cry_7 ),
            .carryinitout(bfn_18_20_0_));
    defparam IN_MUX_bfv_16_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_16_0_));
    defparam IN_MUX_bfv_18_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_13_0_));
    defparam IN_MUX_bfv_18_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_14_0_ (
            .carryinitin(\DUT.uart_inst0.rx_clk_divider_1_cry_7 ),
            .carryinitout(bfn_18_14_0_));
    defparam IN_MUX_bfv_18_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_15_0_ (
            .carryinitin(\DUT.uart_inst0.rx_clk_divider_1_cry_15 ),
            .carryinitout(bfn_18_15_0_));
    defparam IN_MUX_bfv_14_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_19_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_18_0_));
    ICE_GB \top_pll_inst.top_pll_inst_RNISDA2_1  (
            .USERSIGNALTOGLOBALBUFFER(N__10830),
            .GLOBALBUFFEROUTPUT(wPllLocked_iso_i_g));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB \top_pll_inst.top_pll_inst_RNISDA2  (
            .USERSIGNALTOGLOBALBUFFER(N__11536),
            .GLOBALBUFFEROUTPUT(wPllLocked_g));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0 .C_ON=1'b0;
    defparam \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0 .SEQ_MODE=4'b0000;
    defparam \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5143),
            .lcout(wPllLocked),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_12_14_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_12_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__2_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6966),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12109),
            .ce(N__5663),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_12_15_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_12_15_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_12_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__5_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6850),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12102),
            .ce(N__5671),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_12_15_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_12_15_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_12_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__4_LC_12_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6889),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12102),
            .ce(N__5671),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_12_15_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_12_15_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_12_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__3_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6930),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12102),
            .ce(N__5671),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_12_15_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_12_15_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_12_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__6_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6811),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12102),
            .ce(N__5671),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_1_LC_12_16_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_1_LC_12_16_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rWritePtr_1_LC_12_16_0 .LUT_INIT=16'b0000000010110100;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_1_LC_12_16_0  (
            .in0(N__5473),
            .in1(N__5451),
            .in2(N__5425),
            .in3(N__5260),
            .lcout(\DUT.fifo_rx_inst.rWritePtrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12097),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_2_1_LC_12_16_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_2_1_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_2_1_LC_12_16_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI96D91_2_1_LC_12_16_1  (
            .in0(N__5557),
            .in1(N__5418),
            .in2(N__5455),
            .in3(N__7101),
            .lcout(\DUT.fifo_rx_inst.N_86 ),
            .ltout(\DUT.fifo_rx_inst.N_86_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1_1_LC_12_16_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1_1_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1_1_LC_12_16_2 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI5KNB1_1_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5263),
            .in3(N__11506),
            .lcout(\DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1 ),
            .ltout(\DUT.fifo_rx_inst.rWritePtr_RNI5KNB1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_0_LC_12_16_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_0_LC_12_16_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rWritePtr_0_LC_12_16_3 .LUT_INIT=16'b0000101000000101;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_0_LC_12_16_3  (
            .in0(N__5450),
            .in1(_gnd_net_),
            .in2(N__5254),
            .in3(N__5472),
            .lcout(\DUT.fifo_rx_inst.rWritePtrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12097),
            .ce(),
            .sr(_gnd_net_));
    defparam oTx_n_c_sbtinv_LC_12_18_3.C_ON=1'b0;
    defparam oTx_n_c_sbtinv_LC_12_18_3.SEQ_MODE=4'b0000;
    defparam oTx_n_c_sbtinv_LC_12_18_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 oTx_n_c_sbtinv_LC_12_18_3 (
            .in0(N__6204),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(oTx_n_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_0_LC_12_19_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_0_LC_12_19_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoCount_0_LC_12_19_1 .LUT_INIT=16'b1110010000011011;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_0_LC_12_19_1  (
            .in0(N__11619),
            .in1(N__6410),
            .in2(N__6115),
            .in3(N__6154),
            .lcout(\DUT.fifo_tx_inst.rFifoCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12080),
            .ce(),
            .sr(N__12484));
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_LC_12_20_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_LC_12_20_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_LC_12_20_2  (
            .in0(N__7528),
            .in1(N__7619),
            .in2(_gnd_net_),
            .in3(N__6400),
            .lcout(\DUT.fifo_tx_inst.N_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \top_pll_inst.top_pll_inst_RNISDA2_0_LC_12_20_4 .C_ON=1'b0;
    defparam \top_pll_inst.top_pll_inst_RNISDA2_0_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \top_pll_inst.top_pll_inst_RNISDA2_0_LC_12_20_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \top_pll_inst.top_pll_inst_RNISDA2_0_LC_12_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11924),
            .lcout(wPllLocked_iso_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_12_21_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_12_21_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_12_21_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__5_LC_12_21_7  (
            .in0(N__7662),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12076),
            .ce(N__10211),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_12_22_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_12_22_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_12_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__7_LC_12_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7945),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12075),
            .ce(N__10229),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_12_22_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_12_22_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_12_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__4_LC_12_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7716),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12075),
            .ce(N__10229),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_12_22_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_12_22_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_12_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__2_LC_12_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7771),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12075),
            .ce(N__10229),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_13_13_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_13_13_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_13_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__0_LC_13_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7036),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12121),
            .ce(N__5800),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_13_13_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_13_13_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_13_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__1_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7006),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12121),
            .ce(N__5800),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_13_13_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_13_13_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_13_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__2_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6970),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12121),
            .ce(N__5800),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_13_13_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_13_13_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_13_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__3_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6931),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12121),
            .ce(N__5800),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_13_13_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_13_13_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_13_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__4_LC_13_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6888),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12121),
            .ce(N__5800),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_13_13_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_13_13_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_13_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__5_LC_13_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6849),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12121),
            .ce(N__5800),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_13_13_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_13_13_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_13_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__6_LC_13_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6810),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12121),
            .ce(N__5800),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_13_13_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_13_13_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_13_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__7_LC_13_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6772),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12121),
            .ce(N__5800),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_13_14_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_13_14_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_13_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__0_LC_13_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7032),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12115),
            .ce(N__5314),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_13_14_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_13_14_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_13_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__1_LC_13_14_1  (
            .in0(N__7002),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12115),
            .ce(N__5314),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_13_14_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_13_14_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_13_14_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__2_LC_13_14_2  (
            .in0(N__6965),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12115),
            .ce(N__5314),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_13_14_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_13_14_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_13_14_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__3_LC_13_14_3  (
            .in0(N__6923),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12115),
            .ce(N__5314),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_13_14_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_13_14_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_13_14_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__4_LC_13_14_4  (
            .in0(N__6881),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12115),
            .ce(N__5314),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_13_14_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_13_14_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_13_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__5_LC_13_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6842),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12115),
            .ce(N__5314),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_13_14_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_13_14_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_13_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__6_LC_13_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6803),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12115),
            .ce(N__5314),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_13_14_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_13_14_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_13_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram2__7_LC_13_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6768),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12115),
            .ce(N__5314),
            .sr(_gnd_net_));
    defparam rTxByte_esr_4_LC_13_15_0.C_ON=1'b0;
    defparam rTxByte_esr_4_LC_13_15_0.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_4_LC_13_15_0.LUT_INIT=16'b1000100011110101;
    LogicCell40 rTxByte_esr_4_LC_13_15_0 (
            .in0(N__5998),
            .in1(N__5299),
            .in2(N__5293),
            .in3(N__5344),
            .lcout(rTxByteZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12110),
            .ce(N__5706),
            .sr(N__6040));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_13_15_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_13_15_1 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIQ7AF1_5_LC_13_15_1  (
            .in0(N__5900),
            .in1(N__5281),
            .in2(N__6610),
            .in3(N__5995),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rTxByte_esr_5_LC_13_15_2.C_ON=1'b0;
    defparam rTxByte_esr_5_LC_13_15_2.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_5_LC_13_15_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 rTxByte_esr_5_LC_13_15_2 (
            .in0(N__5999),
            .in1(N__5272),
            .in2(N__5266),
            .in3(N__5386),
            .lcout(rTxByteZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12110),
            .ce(N__5706),
            .sr(N__6040));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_13_15_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_13_15_3 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIS9AF1_6_LC_13_15_3  (
            .in0(N__5901),
            .in1(N__5380),
            .in2(N__6595),
            .in3(N__5996),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rTxByte_esr_6_LC_13_15_4.C_ON=1'b0;
    defparam rTxByte_esr_6_LC_13_15_4.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_6_LC_13_15_4.LUT_INIT=16'b1010110100001101;
    LogicCell40 rTxByte_esr_6_LC_13_15_4 (
            .in0(N__6000),
            .in1(N__5371),
            .in2(N__5365),
            .in3(N__5362),
            .lcout(rTxByteZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12110),
            .ce(N__5706),
            .sr(N__6040));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_13_15_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_13_15_5 .LUT_INIT=16'b0101010100011011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIO5AF1_4_LC_13_15_5  (
            .in0(N__5898),
            .in1(N__5353),
            .in2(N__6625),
            .in3(N__5993),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_13_15_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_13_15_6 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIM3AF1_3_LC_13_15_6  (
            .in0(N__5994),
            .in1(N__5338),
            .in2(N__6640),
            .in3(N__5899),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rTxByte_esr_3_LC_13_15_7.C_ON=1'b0;
    defparam rTxByte_esr_3_LC_13_15_7.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_3_LC_13_15_7.LUT_INIT=16'b1010110000001111;
    LogicCell40 rTxByte_esr_3_LC_13_15_7 (
            .in0(N__5329),
            .in1(N__5323),
            .in2(N__5317),
            .in3(N__5997),
            .lcout(rTxByteZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12110),
            .ce(N__5706),
            .sr(N__6040));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_13_16_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_13_16_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_LC_13_16_0  (
            .in0(N__5454),
            .in1(N__5424),
            .in2(_gnd_net_),
            .in3(N__5471),
            .lcout(\DUT.fifo_rx_inst.rFifoData_awe2 ),
            .ltout(\DUT.fifo_rx_inst.rFifoData_awe2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_LC_13_16_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_LC_13_16_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_LC_13_16_1 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_2_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5302),
            .in3(N__5482),
            .lcout(\DUT.fifo_rx_inst.rFifoDataro_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12103),
            .ce(),
            .sr(N__12491));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_3_LC_13_16_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_3_LC_13_16_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_3_LC_13_16_2 .LUT_INIT=16'b1110111011101110;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_3_LC_13_16_2  (
            .in0(N__5491),
            .in1(N__5650),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_rx_inst.rFifoDataro_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12103),
            .ce(),
            .sr(N__12491));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_13_16_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_13_16_3 .LUT_INIT=16'b0010111101111111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_2_RNI4AQO1_LC_13_16_3  (
            .in0(N__5884),
            .in1(N__5490),
            .in2(N__6001),
            .in3(N__5481),
            .lcout(\DUT.fifo_rx_inst.rTxByte_42_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_13_16_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_13_16_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_13_16_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI96D91_1_1_LC_13_16_4  (
            .in0(N__5452),
            .in1(N__5422),
            .in2(_gnd_net_),
            .in3(N__5470),
            .lcout(\DUT.fifo_rx_inst.rFifoData_awe0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_13_16_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_13_16_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNICMVR_2_LC_13_16_5  (
            .in0(_gnd_net_),
            .in1(N__7093),
            .in2(_gnd_net_),
            .in3(N__5556),
            .lcout(\DUT.fifo_rx_inst.N_42 ),
            .ltout(\DUT.fifo_rx_inst.N_42_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_13_16_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_13_16_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_13_16_6 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \DUT.fifo_rx_inst.rWritePtr_RNI96D91_0_1_LC_13_16_6  (
            .in0(N__5453),
            .in1(_gnd_net_),
            .in2(N__5428),
            .in3(N__5423),
            .lcout(\DUT.fifo_rx_inst.rFifoData_awe1 ),
            .ltout(\DUT.fifo_rx_inst.rFifoData_awe1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_1_LC_13_16_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_1_LC_13_16_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_1_LC_13_16_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_1_LC_13_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5401),
            .in3(N__5689),
            .lcout(\DUT.fifo_rx_inst.rFifoDataro_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12103),
            .ce(),
            .sr(N__12491));
    defparam \DUT.fifo_tx_inst.rWritePtr_1_LC_13_17_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_1_LC_13_17_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rWritePtr_1_LC_13_17_0 .LUT_INIT=16'b0000101100000100;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_1_LC_13_17_0  (
            .in0(N__6413),
            .in1(N__7504),
            .in2(N__5398),
            .in3(N__7608),
            .lcout(\DUT.fifo_tx_inst.rWritePtrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12098),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIJLJC_1_LC_13_17_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIJLJC_1_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIJLJC_1_LC_13_17_1 .LUT_INIT=16'b0000111110001111;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_RNIJLJC_1_LC_13_17_1  (
            .in0(N__7502),
            .in1(N__7574),
            .in2(N__11520),
            .in3(N__6411),
            .lcout(\DUT.fifo_tx_inst.un1_i11_i ),
            .ltout(\DUT.fifo_tx_inst.un1_i11_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_0_LC_13_17_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_0_LC_13_17_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rWritePtr_0_LC_13_17_2 .LUT_INIT=16'b0000101000000101;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_0_LC_13_17_2  (
            .in0(N__6412),
            .in1(_gnd_net_),
            .in2(N__5389),
            .in3(N__7503),
            .lcout(\DUT.fifo_tx_inst.rWritePtrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12098),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI9EGD1_0_LC_13_17_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI9EGD1_0_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI9EGD1_0_LC_13_17_3 .LUT_INIT=16'b0011001100110111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNI9EGD1_0_LC_13_17_3  (
            .in0(N__5824),
            .in1(N__8676),
            .in2(N__5521),
            .in3(N__5547),
            .lcout(\DUT.fifo_rx_inst.N_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIK3G92_1_LC_13_17_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIK3G92_1_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIK3G92_1_LC_13_17_4 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNIK3G92_1_LC_13_17_4  (
            .in0(N__7092),
            .in1(N__5518),
            .in2(N__6066),
            .in3(N__8674),
            .lcout(\DUT.fifo_rx_inst.rFifoCount_RNIK3G92Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNO_0_2_LC_13_17_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNO_0_2_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNO_0_2_LC_13_17_5 .LUT_INIT=16'b1100011011001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNO_0_2_LC_13_17_5  (
            .in0(N__8675),
            .in1(N__5548),
            .in2(N__7102),
            .in3(N__6062),
            .lcout(\DUT.fifo_rx_inst.un1_rFifoCount_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_LC_13_17_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_LC_13_17_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNIHH0D1_0_LC_13_17_6  (
            .in0(N__5545),
            .in1(N__5514),
            .in2(_gnd_net_),
            .in3(N__5823),
            .lcout(wRxBufferEmpty_i_0),
            .ltout(wRxBufferEmpty_i_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIL4G92_2_LC_13_17_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIL4G92_2_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNIL4G92_2_LC_13_17_7 .LUT_INIT=16'b1101111110011011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNIL4G92_2_LC_13_17_7  (
            .in0(N__8673),
            .in1(N__7091),
            .in2(N__5587),
            .in3(N__5546),
            .lcout(\DUT.fifo_rx_inst.un1_rFifoCount16_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_inv_LC_13_18_0 .C_ON=1'b1;
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_inv_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_inv_LC_13_18_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0_c_inv_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(N__5584),
            .in2(N__5832),
            .in3(N__5847),
            .lcout(\DUT.fifo_rx_inst.un1_rFifoCount16_0_i_0 ),
            .ltout(),
            .carryin(bfn_13_18_0_),
            .carryout(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_1_LC_13_18_1 .C_ON=1'b1;
    defparam \DUT.fifo_rx_inst.rFifoCount_1_LC_13_18_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoCount_1_LC_13_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_1_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(N__5519),
            .in2(N__5578),
            .in3(N__5569),
            .lcout(\DUT.fifo_rx_inst.rFifoCountZ0Z_1 ),
            .ltout(),
            .carryin(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_0 ),
            .carryout(\DUT.fifo_rx_inst.un1_rFifoCount_1_cry_1 ),
            .clk(N__12091),
            .ce(),
            .sr(N__12488));
    defparam \DUT.fifo_rx_inst.rFifoCount_2_LC_13_18_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_2_LC_13_18_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoCount_2_LC_13_18_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_2_LC_13_18_2  (
            .in0(_gnd_net_),
            .in1(N__5566),
            .in2(_gnd_net_),
            .in3(N__5560),
            .lcout(\DUT.fifo_rx_inst.rFifoCountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12091),
            .ce(),
            .sr(N__12488));
    defparam rRxRead_LC_13_19_1.C_ON=1'b0;
    defparam rRxRead_LC_13_19_1.SEQ_MODE=4'b1000;
    defparam rRxRead_LC_13_19_1.LUT_INIT=16'b1111111111101110;
    LogicCell40 rRxRead_LC_13_19_1 (
            .in0(N__5555),
            .in1(N__5520),
            .in2(_gnd_net_),
            .in3(N__5836),
            .lcout(rRxReadZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12086),
            .ce(),
            .sr(N__12486));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIF689_0_LC_13_19_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIF689_0_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIF689_0_LC_13_19_2 .LUT_INIT=16'b1111000011110001;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNIF689_0_LC_13_19_2  (
            .in0(N__7472),
            .in1(N__6145),
            .in2(N__8681),
            .in3(N__8621),
            .lcout(\DUT.fifo_tx_inst.N_35 ),
            .ltout(\DUT.fifo_tx_inst.N_35_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_13_19_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_13_19_3 .LUT_INIT=16'b0000110000111111;
    LogicCell40 \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNO_LC_13_19_3  (
            .in0(N__6146),
            .in1(N__11617),
            .in2(N__5494),
            .in3(N__6392),
            .lcout(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIMBD3_2_LC_13_19_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIMBD3_2_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIMBD3_2_LC_13_19_4 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNIMBD3_2_LC_13_19_4  (
            .in0(N__7471),
            .in1(_gnd_net_),
            .in2(N__8680),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_tx_inst.N_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIN9O8_0_LC_13_19_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIN9O8_0_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIN9O8_0_LC_13_19_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNIN9O8_0_LC_13_19_6  (
            .in0(N__7470),
            .in1(N__6144),
            .in2(_gnd_net_),
            .in3(N__8620),
            .lcout(\DUT.N_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_1_LC_13_20_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_1_LC_13_20_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_1_LC_13_20_3 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_1_LC_13_20_3  (
            .in0(N__7611),
            .in1(N__6304),
            .in2(N__7547),
            .in3(N__6408),
            .lcout(\DUT.fifo_tx_inst.rFifoDataro_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12081),
            .ce(),
            .sr(N__12485));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_LC_13_20_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_LC_13_20_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_LC_13_20_7 .LUT_INIT=16'b1100110011001101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_0_LC_13_20_7  (
            .in0(N__7610),
            .in1(N__6292),
            .in2(N__7546),
            .in3(N__6407),
            .lcout(\DUT.fifo_tx_inst.rFifoDataro_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12081),
            .ce(),
            .sr(N__12485));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_13_21_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_13_21_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_13_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__0_LC_13_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8929),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12079),
            .ce(N__6349),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_13_21_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_13_21_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_13_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__1_LC_13_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8983),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12079),
            .ce(N__6349),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_13_21_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_13_21_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_13_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__2_LC_13_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7756),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12079),
            .ce(N__6349),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_13_21_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_13_21_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_13_21_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__3_LC_13_21_3  (
            .in0(N__10267),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12079),
            .ce(N__6349),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_13_21_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_13_21_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_13_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__4_LC_13_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7705),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12079),
            .ce(N__6349),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_13_21_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_13_21_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_13_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__5_LC_13_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7660),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12079),
            .ce(N__6349),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_13_21_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_13_21_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_13_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__6_LC_13_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8866),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12079),
            .ce(N__6349),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_13_21_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_13_21_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_13_21_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__7_LC_13_21_7  (
            .in0(N__7936),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12079),
            .ce(N__6349),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_13_22_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_13_22_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_13_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__7_LC_13_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7937),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12077),
            .ce(N__6579),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_13_22_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_13_22_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_13_22_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__2_LC_13_22_1  (
            .in0(N__7766),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12077),
            .ce(N__6579),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_13_22_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_13_22_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_13_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__3_LC_13_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10268),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12077),
            .ce(N__6579),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_13_22_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_13_22_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_13_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__0_LC_13_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8937),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12077),
            .ce(N__6579),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_13_22_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_13_22_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_13_22_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__5_LC_13_22_4  (
            .in0(_gnd_net_),
            .in1(N__7661),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12077),
            .ce(N__6579),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_13_22_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_13_22_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_13_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__1_LC_13_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8984),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12077),
            .ce(N__6579),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_13_22_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_13_22_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_13_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__4_LC_13_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7715),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12077),
            .ce(N__6579),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_0_1_LC_13_23_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_0_1_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_0_1_LC_13_23_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_RNIN79A_0_1_LC_13_23_2  (
            .in0(N__7545),
            .in1(N__7609),
            .in2(_gnd_net_),
            .in3(N__6414),
            .lcout(\DUT.fifo_tx_inst.N_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_1_LC_14_11_4 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_1_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_1_LC_14_11_4 .LUT_INIT=16'b0001010001000100;
    LogicCell40 \fifo_inst.ftdi_input_inst.rPacketCount_latch_1_LC_14_11_4  (
            .in0(N__12528),
            .in1(N__6691),
            .in2(N__6730),
            .in3(N__6480),
            .lcout(G_143),
            .ltout(G_143_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.SUM_2_LC_14_11_5 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.SUM_2_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.SUM_2_LC_14_11_5 .LUT_INIT=16'b0011110011001100;
    LogicCell40 \fifo_inst.ftdi_input_inst.SUM_2_LC_14_11_5  (
            .in0(_gnd_net_),
            .in1(N__6549),
            .in2(N__5677),
            .in3(N__6725),
            .lcout(),
            .ltout(\fifo_inst.ftdi_input_inst.SUMZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_2_LC_14_11_6 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_2_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_2_LC_14_11_6 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \fifo_inst.ftdi_input_inst.rPacketCount_latch_2_LC_14_11_6  (
            .in0(N__12529),
            .in1(N__6550),
            .in2(N__5674),
            .in3(N__6481),
            .lcout(G_144),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_14_13_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_14_13_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_14_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__0_LC_14_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7031),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12127),
            .ce(N__5670),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_14_13_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_14_13_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_14_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__1_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7001),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12127),
            .ce(N__5670),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_14_13_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_14_13_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_14_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram3__7_LC_14_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6764),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12127),
            .ce(N__5670),
            .sr(_gnd_net_));
    defparam rTxByte_esr_7_LC_14_14_0.C_ON=1'b0;
    defparam rTxByte_esr_7_LC_14_14_0.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_7_LC_14_14_0.LUT_INIT=16'b1010000011011101;
    LogicCell40 rTxByte_esr_7_LC_14_14_0 (
            .in0(N__6012),
            .in1(N__5632),
            .in2(N__5623),
            .in3(N__5737),
            .lcout(rTxByteZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12122),
            .ce(N__5707),
            .sr(N__6036));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_14_14_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_14_14_1 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIK1AF1_2_LC_14_14_1  (
            .in0(N__5614),
            .in1(N__6008),
            .in2(N__6649),
            .in3(N__5905),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rTxByte_esr_2_LC_14_14_2.C_ON=1'b0;
    defparam rTxByte_esr_2_LC_14_14_2.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_2_LC_14_14_2.LUT_INIT=16'b1010110100001101;
    LogicCell40 rTxByte_esr_2_LC_14_14_2 (
            .in0(N__6011),
            .in1(N__5608),
            .in2(N__5599),
            .in3(N__5596),
            .lcout(rTxByteZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12122),
            .ce(N__5707),
            .sr(N__6036));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_14_14_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_14_14_3 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIIV9F1_1_LC_14_14_3  (
            .in0(N__5770),
            .in1(N__6007),
            .in2(N__6658),
            .in3(N__5904),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rTxByte_esr_1_LC_14_14_4.C_ON=1'b0;
    defparam rTxByte_esr_1_LC_14_14_4.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_1_LC_14_14_4.LUT_INIT=16'b1010110100001101;
    LogicCell40 rTxByte_esr_1_LC_14_14_4 (
            .in0(N__6010),
            .in1(N__5764),
            .in2(N__5755),
            .in3(N__5752),
            .lcout(rTxByteZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12122),
            .ce(N__5707),
            .sr(N__6036));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_14_14_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_14_14_5 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIUBAF1_7_LC_14_14_5  (
            .in0(N__5743),
            .in1(N__6003),
            .in2(N__7060),
            .in3(N__5902),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_14_14_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_14_14_6 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram0__RNIGT9F1_0_LC_14_14_6  (
            .in0(N__5903),
            .in1(N__6664),
            .in2(N__6013),
            .in3(N__5731),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rTxByte_esr_0_LC_14_14_7.C_ON=1'b0;
    defparam rTxByte_esr_0_LC_14_14_7.SEQ_MODE=4'b1000;
    defparam rTxByte_esr_0_LC_14_14_7.LUT_INIT=16'b1100101000001111;
    LogicCell40 rTxByte_esr_0_LC_14_14_7 (
            .in0(N__5725),
            .in1(N__5716),
            .in2(N__5710),
            .in3(N__6009),
            .lcout(rTxByteZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12122),
            .ce(N__5707),
            .sr(N__6036));
    defparam \DUT.uart_inst0.rx_bits_remaining_3_LC_14_15_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_3_LC_14_15_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_bits_remaining_3_LC_14_15_0 .LUT_INIT=16'b1110111011101101;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_3_LC_14_15_0  (
            .in0(N__7152),
            .in1(N__8157),
            .in2(N__7234),
            .in3(N__7194),
            .lcout(\DUT.uart_inst0.rx_bits_remainingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12116),
            .ce(N__7213),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_0_LC_14_15_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_0_LC_14_15_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_bits_remaining_0_LC_14_15_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_0_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__8156),
            .in2(_gnd_net_),
            .in3(N__7135),
            .lcout(\DUT.uart_inst0.rx_bits_remainingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12116),
            .ce(N__7213),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI250E6_0_LC_14_15_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI250E6_0_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoCount_RNI250E6_0_LC_14_15_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_RNI250E6_0_LC_14_15_7  (
            .in0(_gnd_net_),
            .in1(N__6067),
            .in2(_gnd_net_),
            .in3(N__6024),
            .lcout(wRxBufferEmpty_i_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNI0AQO1_LC_14_16_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNI0AQO1_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNI0AQO1_LC_14_16_0 .LUT_INIT=16'b1111010111110011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_0_RNI0AQO1_LC_14_16_0  (
            .in0(N__5688),
            .in1(N__5781),
            .in2(N__6002),
            .in3(N__5885),
            .lcout(),
            .ltout(\DUT.fifo_rx_inst.rTxByte_42_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNIHJV05_LC_14_16_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNIHJV05_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_RNIHJV05_LC_14_16_1 .LUT_INIT=16'b1101010101010101;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_0_RNIHJV05_LC_14_16_1  (
            .in0(N__11502),
            .in1(N__6076),
            .in2(N__6070),
            .in3(N__6058),
            .lcout(rFifoDatarff_0_RNIHJV05),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rReadPtr_1_LC_14_16_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rReadPtr_1_LC_14_16_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rReadPtr_1_LC_14_16_2 .LUT_INIT=16'b0010000100100010;
    LogicCell40 \DUT.fifo_rx_inst.rReadPtr_1_LC_14_16_2  (
            .in0(N__5975),
            .in1(N__5929),
            .in2(N__5923),
            .in3(N__5888),
            .lcout(\DUT.fifo_rx_inst.rReadPtrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12111),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rReadPtr_RNI4NC92_0_LC_14_16_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rReadPtr_RNI4NC92_0_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_rx_inst.rReadPtr_RNI4NC92_0_LC_14_16_3 .LUT_INIT=16'b0010111100001111;
    LogicCell40 \DUT.fifo_rx_inst.rReadPtr_RNI4NC92_0_LC_14_16_3  (
            .in0(N__5886),
            .in1(N__5918),
            .in2(N__11524),
            .in3(N__5974),
            .lcout(\DUT.fifo_rx_inst.rReadPtr_RNI4NC92Z0Z_0 ),
            .ltout(\DUT.fifo_rx_inst.rReadPtr_RNI4NC92Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rReadPtr_0_LC_14_16_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rReadPtr_0_LC_14_16_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rReadPtr_0_LC_14_16_4 .LUT_INIT=16'b0000101000000101;
    LogicCell40 \DUT.fifo_rx_inst.rReadPtr_0_LC_14_16_4  (
            .in0(N__5919),
            .in1(_gnd_net_),
            .in2(N__5908),
            .in3(N__5887),
            .lcout(\DUT.fifo_rx_inst.rReadPtrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12111),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_6_LC_14_16_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_6_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_6_LC_14_16_6 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_6_LC_14_16_6  (
            .in0(N__8238),
            .in1(N__11922),
            .in2(_gnd_net_),
            .in3(N__8261),
            .lcout(),
            .ltout(\DUT.uart_inst0.recv_state_srsts_1_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_6_LC_14_16_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_6_LC_14_16_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_6_LC_14_16_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.recv_state_6_LC_14_16_7  (
            .in0(N__8014),
            .in1(N__8431),
            .in2(N__5851),
            .in3(N__8366),
            .lcout(\DUT.wRcvd ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12111),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoCount_0_LC_14_17_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoCount_0_LC_14_17_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoCount_0_LC_14_17_1 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \DUT.fifo_rx_inst.rFifoCount_0_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(N__5831),
            .in2(_gnd_net_),
            .in3(N__5848),
            .lcout(\DUT.fifo_rx_inst.rFifoCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12104),
            .ce(),
            .sr(N__12492));
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_LC_14_17_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_LC_14_17_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoDatarff_0_LC_14_17_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_rx_inst.rFifoDatarff_0_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(N__5793),
            .in2(_gnd_net_),
            .in3(N__5782),
            .lcout(\DUT.fifo_rx_inst.rFifoDataro_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12104),
            .ce(),
            .sr(N__12492));
    defparam \fifo_inst.ftdi_output_inst.oTx_n_LC_14_17_3 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.oTx_n_LC_14_17_3 .SEQ_MODE=4'b1001;
    defparam \fifo_inst.ftdi_output_inst.oTx_n_LC_14_17_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \fifo_inst.ftdi_output_inst.oTx_n_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(N__6192),
            .in2(_gnd_net_),
            .in3(N__9250),
            .lcout(oTx_n_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12104),
            .ce(),
            .sr(N__12492));
    defparam \fifo_inst.ftdi_output_inst.rWrDelay_LC_14_17_4 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rWrDelay_LC_14_17_4 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rWrDelay_LC_14_17_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \fifo_inst.ftdi_output_inst.rWrDelay_LC_14_17_4  (
            .in0(_gnd_net_),
            .in1(N__11044),
            .in2(_gnd_net_),
            .in3(N__11005),
            .lcout(\fifo_inst.ftdi_output_inst.rWrDelayZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12104),
            .ce(),
            .sr(N__12492));
    defparam \fifo_inst.ftdi_output_inst.oRxFlag_LC_14_18_6 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.oRxFlag_LC_14_18_6 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.oRxFlag_LC_14_18_6 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \fifo_inst.ftdi_output_inst.oRxFlag_LC_14_18_6  (
            .in0(N__6165),
            .in1(N__11296),
            .in2(_gnd_net_),
            .in3(N__9235),
            .lcout(P1A2_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12099),
            .ce(),
            .sr(N__12490));
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_14_19_0 .C_ON=1'b1;
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_14_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0_c_LC_14_19_0  (
            .in0(_gnd_net_),
            .in1(N__6153),
            .in2(N__6127),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_19_0_),
            .carryout(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_1_LC_14_19_1 .C_ON=1'b1;
    defparam \DUT.fifo_tx_inst.rFifoCount_1_LC_14_19_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoCount_1_LC_14_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_1_LC_14_19_1  (
            .in0(_gnd_net_),
            .in1(N__8622),
            .in2(N__8602),
            .in3(N__6118),
            .lcout(\DUT.fifo_tx_inst.rFifoCountZ0Z_1 ),
            .ltout(),
            .carryin(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_0 ),
            .carryout(\DUT.fifo_tx_inst.un1_rFifoCount_1_cry_1 ),
            .clk(N__12092),
            .ce(),
            .sr(N__12489));
    defparam \DUT.fifo_tx_inst.rFifoCount_2_LC_14_19_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_2_LC_14_19_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoCount_2_LC_14_19_2 .LUT_INIT=16'b0011100111000110;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_2_LC_14_19_2  (
            .in0(N__11618),
            .in1(N__7474),
            .in2(N__6114),
            .in3(N__6097),
            .lcout(\DUT.fifo_tx_inst.rFifoCountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12092),
            .ce(),
            .sr(N__12489));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_3_LC_14_20_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_3_LC_14_20_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_3_LC_14_20_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_3_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(N__7896),
            .in2(_gnd_net_),
            .in3(N__6094),
            .lcout(\DUT.fifo_tx_inst.rFifoDataro_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12087),
            .ce(),
            .sr(N__12487));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_LC_14_20_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_LC_14_20_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_LC_14_20_2 .LUT_INIT=16'b1010101010111010;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_2_LC_14_20_2  (
            .in0(N__6085),
            .in1(N__7541),
            .in2(N__7621),
            .in3(N__6409),
            .lcout(\DUT.fifo_tx_inst.rFifoDataro_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12087),
            .ce(),
            .sr(N__12487));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_14_20_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_14_20_3 .LUT_INIT=16'b0010010101110101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_2_RNIC6BE_LC_14_20_3  (
            .in0(N__7384),
            .in1(N__6093),
            .in2(N__9670),
            .in3(N__6084),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoDataror_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_RNIJBAM_LC_14_20_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_RNIJBAM_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoDatarff_0_RNIJBAM_LC_14_20_4 .LUT_INIT=16'b1111000000110101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoDatarff_0_RNIJBAM_LC_14_20_4  (
            .in0(N__6303),
            .in1(N__6291),
            .in2(N__6280),
            .in3(N__9642),
            .lcout(\DUT.rFifoDataror_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_14_20_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_14_20_5 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIOH0H_0_LC_14_20_5  (
            .in0(N__7385),
            .in1(N__6277),
            .in2(N__9671),
            .in3(N__6268),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_14_20_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_14_20_6 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIJIDC1_0_LC_14_20_6  (
            .in0(N__7780),
            .in1(N__8890),
            .in2(N__6262),
            .in3(N__9643),
            .lcout(\DUT.rFifoDatarxZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rReadPtr_RNILV421_1_LC_14_21_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rReadPtr_RNILV421_1_LC_14_21_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rReadPtr_RNILV421_1_LC_14_21_0 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \DUT.fifo_tx_inst.rReadPtr_RNILV421_1_LC_14_21_0  (
            .in0(N__11501),
            .in1(N__9650),
            .in2(_gnd_net_),
            .in3(N__6229),
            .lcout(\DUT.fifo_tx_inst.un1_i11_2_i ),
            .ltout(\DUT.fifo_tx_inst.un1_i11_2_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rReadPtr_0_LC_14_21_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rReadPtr_0_LC_14_21_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rReadPtr_0_LC_14_21_1 .LUT_INIT=16'b0000101100000100;
    LogicCell40 \DUT.fifo_tx_inst.rReadPtr_0_LC_14_21_1  (
            .in0(N__8576),
            .in1(N__11621),
            .in2(N__6259),
            .in3(N__7392),
            .lcout(\DUT.fifo_tx_inst.rReadPtrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12082),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_14_21_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_14_21_2 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIQJ0H_1_LC_14_21_2  (
            .in0(N__6256),
            .in1(N__9647),
            .in2(N__6250),
            .in3(N__7382),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_14_21_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_14_21_3 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNIUN0H_3_LC_14_21_3  (
            .in0(N__7380),
            .in1(N__6241),
            .in2(N__9672),
            .in3(N__6235),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rReadPtr_RNINFEP_0_LC_14_21_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rReadPtr_RNINFEP_0_LC_14_21_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rReadPtr_RNINFEP_0_LC_14_21_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \DUT.fifo_tx_inst.rReadPtr_RNINFEP_0_LC_14_21_4  (
            .in0(N__11620),
            .in1(N__7383),
            .in2(_gnd_net_),
            .in3(N__8575),
            .lcout(\DUT.fifo_tx_inst.CO0 ),
            .ltout(\DUT.fifo_tx_inst.CO0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rReadPtr_1_LC_14_21_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rReadPtr_1_LC_14_21_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rReadPtr_1_LC_14_21_5 .LUT_INIT=16'b0000000001011010;
    LogicCell40 \DUT.fifo_tx_inst.rReadPtr_1_LC_14_21_5  (
            .in0(N__9651),
            .in1(_gnd_net_),
            .in2(N__6223),
            .in3(N__6220),
            .lcout(\DUT.fifo_tx_inst.rReadPtrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12082),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_14_21_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_14_21_6 .LUT_INIT=16'b0000001111011101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI2S0H_5_LC_14_21_6  (
            .in0(N__6466),
            .in1(N__9648),
            .in2(N__6460),
            .in3(N__7381),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_14_21_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_14_21_7 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_14_21_7 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI77EC1_5_LC_14_21_7  (
            .in0(N__9649),
            .in1(N__7633),
            .in2(N__6451),
            .in3(N__6448),
            .lcout(\DUT.rFifoDatarx_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_14_22_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_14_22_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_14_22_0 .LUT_INIT=16'b0001110000011111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI601H_7_LC_14_22_0  (
            .in0(N__6439),
            .in1(N__9652),
            .in2(N__7393),
            .in3(N__6433),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_14_22_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_14_22_1 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_14_22_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIFFEC1_7_LC_14_22_1  (
            .in0(N__9656),
            .in1(N__7909),
            .in2(N__6427),
            .in3(N__6424),
            .lcout(\DUT.rFifoDatarx_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_1_LC_14_22_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_1_LC_14_22_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_1_LC_14_22_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DUT.fifo_tx_inst.rWritePtr_RNIN79A_1_1_LC_14_22_2  (
            .in0(N__7548),
            .in1(N__7620),
            .in2(_gnd_net_),
            .in3(N__6415),
            .lcout(\DUT.fifo_tx_inst.N_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_14_22_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_14_22_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_14_22_3 .LUT_INIT=16'b0011010000110111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI0Q0H_4_LC_14_22_3  (
            .in0(N__6343),
            .in1(N__7386),
            .in2(N__9673),
            .in3(N__6337),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_14_22_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_14_22_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_14_22_4 .LUT_INIT=16'b0101001001010111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNISL0H_2_LC_14_22_4  (
            .in0(N__7390),
            .in1(N__6331),
            .in2(N__9674),
            .in3(N__6325),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_14_22_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_14_22_5 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_14_22_5 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIRQDC1_2_LC_14_22_5  (
            .in0(N__9657),
            .in1(N__7726),
            .in2(N__6319),
            .in3(N__6316),
            .lcout(),
            .ltout(\DUT.rFifoDatarx_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_RNO_0_2_LC_14_22_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_RNO_0_2_LC_14_22_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_data_RNO_0_2_LC_14_22_6 .LUT_INIT=16'b1000100010111000;
    LogicCell40 \DUT.uart_inst0.tx_data_RNO_0_2_LC_14_22_6  (
            .in0(N__9910),
            .in1(N__12674),
            .in2(N__6307),
            .in3(N__10041),
            .lcout(\DUT.uart_inst0.tx_data_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_14_23_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_14_23_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_14_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram1__6_LC_14_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8878),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12078),
            .ce(N__6580),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.rWrState_latch_1_LC_15_10_3 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.rWrState_latch_1_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.rWrState_latch_1_LC_15_10_3 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \fifo_inst.ftdi_input_inst.rWrState_latch_1_LC_15_10_3  (
            .in0(N__11918),
            .in1(N__6675),
            .in2(_gnd_net_),
            .in3(N__6564),
            .lcout(G_145),
            .ltout(G_145_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.rRamWrEn_latch_LC_15_10_4 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.rRamWrEn_latch_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.rRamWrEn_latch_LC_15_10_4 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \fifo_inst.ftdi_input_inst.rRamWrEn_latch_LC_15_10_4  (
            .in0(N__6674),
            .in1(N__6515),
            .in2(N__6568),
            .in3(N__12534),
            .lcout(G_147),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.un1_rWrState_1_LC_15_10_7 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.un1_rWrState_1_LC_15_10_7 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.un1_rWrState_1_LC_15_10_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \fifo_inst.ftdi_input_inst.un1_rWrState_1_LC_15_10_7  (
            .in0(_gnd_net_),
            .in1(N__6676),
            .in2(_gnd_net_),
            .in3(N__6565),
            .lcout(\fifo_inst.ftdi_input_inst.un1_rWrStateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.un2_oPacketAvail_i_LC_15_11_0 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.un2_oPacketAvail_i_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.un2_oPacketAvail_i_LC_15_11_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \fifo_inst.ftdi_input_inst.un2_oPacketAvail_i_LC_15_11_0  (
            .in0(N__6553),
            .in1(N__6498),
            .in2(N__6729),
            .in3(N__6694),
            .lcout(\fifo_inst.ftdi_input_inst.un2_oPacketAvail_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_3_LC_15_11_1 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_3_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_3_LC_15_11_1 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \fifo_inst.ftdi_input_inst.rPacketCount_latch_3_LC_15_11_1  (
            .in0(N__6497),
            .in1(N__6479),
            .in2(N__12540),
            .in3(N__6529),
            .lcout(G_142),
            .ltout(G_142_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.oTxFull_0_LC_15_11_2 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.oTxFull_0_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.oTxFull_0_LC_15_11_2 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \fifo_inst.ftdi_input_inst.oTxFull_0_LC_15_11_2  (
            .in0(N__6552),
            .in1(_gnd_net_),
            .in2(N__6556),
            .in3(_gnd_net_),
            .lcout(fifo_inst_ftdi_input_inst_oTxFull_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.SUM_3_LC_15_11_3 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.SUM_3_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.SUM_3_LC_15_11_3 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \fifo_inst.ftdi_input_inst.SUM_3_LC_15_11_3  (
            .in0(N__6693),
            .in1(N__6551),
            .in2(N__6499),
            .in3(N__6720),
            .lcout(\fifo_inst.ftdi_input_inst.SUMZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.rPacketCount15_LC_15_11_4 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.rPacketCount15_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.rPacketCount15_LC_15_11_4 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \fifo_inst.ftdi_input_inst.rPacketCount15_LC_15_11_4  (
            .in0(N__6516),
            .in1(N__6496),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(G_141),
            .ltout(G_141_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_0_LC_15_11_5 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_0_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.rPacketCount_latch_0_LC_15_11_5 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \fifo_inst.ftdi_input_inst.rPacketCount_latch_0_LC_15_11_5  (
            .in0(N__12530),
            .in1(_gnd_net_),
            .in2(N__6733),
            .in3(N__6721),
            .lcout(G_140),
            .ltout(G_140_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.wTxEn_1_LC_15_11_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.wTxEn_1_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.wTxEn_1_LC_15_11_6 .LUT_INIT=16'b1100110011000100;
    LogicCell40 \DUT.uart_inst0.wTxEn_1_LC_15_11_6  (
            .in0(N__6703),
            .in1(N__11919),
            .in2(N__6697),
            .in3(N__6692),
            .lcout(G_146),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_15_13_0 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_15_13_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_15_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__0_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7024),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12132),
            .ce(N__7051),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_15_13_1 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_15_13_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_15_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__1_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6994),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12132),
            .ce(N__7051),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_15_13_2 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_15_13_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_15_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__2_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6955),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12132),
            .ce(N__7051),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_15_13_3 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_15_13_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_15_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__3_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6913),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12132),
            .ce(N__7051),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_15_13_4 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_15_13_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_15_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__4_LC_15_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6871),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12132),
            .ce(N__7051),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_15_13_5 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_15_13_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_15_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__5_LC_15_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6832),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12132),
            .ce(N__7051),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_15_13_6 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_15_13_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_15_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__6_LC_15_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6793),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12132),
            .ce(N__7051),
            .sr(_gnd_net_));
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_15_13_7 .C_ON=1'b0;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_15_13_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_15_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_rx_inst.rFifoData_rFifoData_ram1__7_LC_15_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6760),
            .lcout(\DUT.fifo_rx_inst.rFifoData_ram1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12132),
            .ce(N__7051),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_0_LC_15_14_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_0_LC_15_14_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_0_LC_15_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_0_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6993),
            .lcout(\DUT.wRxByte_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12128),
            .ce(N__7114),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_1_LC_15_14_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_1_LC_15_14_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_1_LC_15_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_1_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6954),
            .lcout(\DUT.wRxByte_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12128),
            .ce(N__7114),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_2_LC_15_14_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_2_LC_15_14_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_2_LC_15_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_2_LC_15_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6912),
            .lcout(\DUT.wRxByte_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12128),
            .ce(N__7114),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_3_LC_15_14_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_3_LC_15_14_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_3_LC_15_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_3_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6870),
            .lcout(\DUT.wRxByte_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12128),
            .ce(N__7114),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_4_LC_15_14_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_4_LC_15_14_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_4_LC_15_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_4_LC_15_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6831),
            .lcout(\DUT.wRxByte_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12128),
            .ce(N__7114),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_5_LC_15_14_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_5_LC_15_14_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_5_LC_15_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_5_LC_15_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6792),
            .lcout(\DUT.wRxByte_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12128),
            .ce(N__7114),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_6_LC_15_14_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_6_LC_15_14_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_6_LC_15_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_data_6_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6759),
            .lcout(\DUT.wRxByte_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12128),
            .ce(N__7114),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_data_7_LC_15_14_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_data_7_LC_15_14_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_data_7_LC_15_14_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DUT.uart_inst0.rx_data_7_LC_15_14_7  (
            .in0(N__8223),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DUT.wRxByte_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12128),
            .ce(N__7114),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNIQJ1OI_2_LC_15_15_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNIQJ1OI_2_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNIQJ1OI_2_LC_15_15_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \DUT.uart_inst0.recv_state_RNIQJ1OI_2_LC_15_15_0  (
            .in0(N__7312),
            .in1(N__8418),
            .in2(N__8367),
            .in3(N__8010),
            .lcout(\DUT.uart_inst0.rx_bits_remaining_2_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNITG1J4_LC_15_15_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNITG1J4_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNITG1J4_LC_15_15_1 .LUT_INIT=16'b1001101010101010;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNITG1J4_LC_15_15_1  (
            .in0(N__8314),
            .in1(N__8089),
            .in2(N__8059),
            .in3(N__9196),
            .lcout(\DUT.uart_inst0.rx_countdown_3_2 ),
            .ltout(\DUT.uart_inst0.rx_countdown_3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_15_15_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_15_15_2 .LUT_INIT=16'b0000000011010000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_1_2_LC_15_15_2  (
            .in0(N__8041),
            .in1(N__8228),
            .in2(N__7105),
            .in3(N__8289),
            .lcout(\DUT.uart_inst0.rx_countdown_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_0_LC_15_15_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_0_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_0_LC_15_15_3 .LUT_INIT=16'b0000000000101010;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_0_LC_15_15_3  (
            .in0(N__11921),
            .in1(N__8039),
            .in2(N__8239),
            .in3(N__7100),
            .lcout(\DUT.uart_inst0.recv_state_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIT7PG_1_LC_15_15_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIT7PG_1_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIT7PG_1_LC_15_15_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNIT7PG_1_LC_15_15_4  (
            .in0(N__7138),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7177),
            .lcout(\DUT.uart_inst0.N_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_5_LC_15_15_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_5_LC_15_15_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_5_LC_15_15_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.recv_state_5_LC_15_15_6  (
            .in0(N__8116),
            .in1(N__8011),
            .in2(N__8368),
            .in3(N__8419),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12123),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNIHH651_0_LC_15_15_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNIHH651_0_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNIHH651_0_LC_15_15_7 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \DUT.uart_inst0.recv_state_RNIHH651_0_LC_15_15_7  (
            .in0(N__8290),
            .in1(N__8224),
            .in2(_gnd_net_),
            .in3(N__8040),
            .lcout(\DUT.uart_inst0.N_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNIEMU42_5_LC_15_16_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNIEMU42_5_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNIEMU42_5_LC_15_16_0 .LUT_INIT=16'b0000000111001101;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNIEMU42_5_LC_15_16_0  (
            .in0(N__8540),
            .in1(N__9069),
            .in2(N__9169),
            .in3(N__9180),
            .lcout(),
            .ltout(\DUT.uart_inst0.rx_countdown_8_i_o2_2_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNIDB3D7_0_LC_15_16_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNIDB3D7_0_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNIDB3D7_0_LC_15_16_1 .LUT_INIT=16'b1101111110101111;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNIDB3D7_0_LC_15_16_1  (
            .in0(N__9070),
            .in1(N__8103),
            .in2(N__7063),
            .in3(N__9127),
            .lcout(\DUT.uart_inst0.rx_countdown_8_i_o2_2_2 ),
            .ltout(\DUT.uart_inst0.rx_countdown_8_i_o2_2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNIIQN8I_LC_15_16_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNIIQN8I_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNIIQN8I_LC_15_16_2 .LUT_INIT=16'b0000000100000001;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_1_s1_c_RNIIQN8I_LC_15_16_2  (
            .in0(N__8416),
            .in1(N__8008),
            .in2(N__7243),
            .in3(_gnd_net_),
            .lcout(\DUT.uart_inst0.recv_N_5_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_1_LC_15_16_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_1_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_1_LC_15_16_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_1_LC_15_16_3  (
            .in0(N__8009),
            .in1(N__8417),
            .in2(N__8369),
            .in3(N__11194),
            .lcout(),
            .ltout(\DUT.uart_inst0.recv_state_RNO_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_1_LC_15_16_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_1_LC_15_16_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_1_LC_15_16_4 .LUT_INIT=16'b0000110000000100;
    LogicCell40 \DUT.uart_inst0.recv_state_1_LC_15_16_4  (
            .in0(N__11195),
            .in1(N__11527),
            .in2(N__7240),
            .in3(N__8158),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12117),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNIBTG71_2_LC_15_16_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNIBTG71_2_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNIBTG71_2_LC_15_16_5 .LUT_INIT=16'b1111000001000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNIBTG71_2_LC_15_16_5  (
            .in0(N__8229),
            .in1(N__8150),
            .in2(N__11535),
            .in3(N__7290),
            .lcout(),
            .ltout(\DUT.uart_inst0.un1_m2_e_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNITN8GJ_2_LC_15_16_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNITN8GJ_2_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNITN8GJ_2_LC_15_16_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNITN8GJ_2_LC_15_16_6  (
            .in0(N__8415),
            .in1(N__8007),
            .in2(N__7237),
            .in3(N__8355),
            .lcout(\DUT.uart_inst0.recv_state_RNITN8GJZ0Z_2 ),
            .ltout(\DUT.uart_inst0.recv_state_RNITN8GJZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_2_LC_15_16_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_2_LC_15_16_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_bits_remaining_2_LC_15_16_7 .LUT_INIT=16'b0010111100010000;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_2_LC_15_16_7  (
            .in0(N__7233),
            .in1(N__8151),
            .in2(N__7216),
            .in3(N__7195),
            .lcout(\DUT.uart_inst0.rx_bits_remainingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12117),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_15_17_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_15_17_0 .LUT_INIT=16'b0100010001010101;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_0_2_LC_15_17_0  (
            .in0(N__7292),
            .in1(N__8242),
            .in2(_gnd_net_),
            .in3(N__8152),
            .lcout(\DUT.uart_inst0.rx_countdown_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNI8P9F_2_LC_15_17_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNI8P9F_2_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNI8P9F_2_LC_15_17_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNI8P9F_2_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(N__11925),
            .in2(_gnd_net_),
            .in3(N__7291),
            .lcout(\DUT.uart_inst0.rx_m2_e_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_1_LC_15_17_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_1_LC_15_17_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_bits_remaining_1_LC_15_17_2 .LUT_INIT=16'b0010000111110000;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_1_LC_15_17_2  (
            .in0(N__7137),
            .in1(N__8154),
            .in2(N__7176),
            .in3(N__7206),
            .lcout(\DUT.uart_inst0.rx_bits_remainingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12112),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIUJI11_3_LC_15_17_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIUJI11_3_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_bits_remaining_RNIUJI11_3_LC_15_17_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \DUT.uart_inst0.rx_bits_remaining_RNIUJI11_3_LC_15_17_3  (
            .in0(N__7193),
            .in1(N__7169),
            .in2(N__7156),
            .in3(N__7136),
            .lcout(\DUT.uart_inst0.N_98_4 ),
            .ltout(\DUT.uart_inst0.N_98_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_2_LC_15_17_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_2_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_2_LC_15_17_4 .LUT_INIT=16'b1100010011110101;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_2_LC_15_17_4  (
            .in0(N__7294),
            .in1(N__8241),
            .in2(N__7315),
            .in3(N__8153),
            .lcout(),
            .ltout(\DUT.uart_inst0.r_N_5_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_2_LC_15_17_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_2_LC_15_17_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_2_LC_15_17_5 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \DUT.uart_inst0.recv_state_2_LC_15_17_5  (
            .in0(N__11525),
            .in1(N__7311),
            .in2(N__7297),
            .in3(N__7263),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12112),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_3_LC_15_17_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_3_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_3_LC_15_17_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_3_LC_15_17_6  (
            .in0(N__7293),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7273),
            .lcout(),
            .ltout(\DUT.uart_inst0.r_N_3_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_3_LC_15_17_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_3_LC_15_17_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_3_LC_15_17_7 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \DUT.uart_inst0.recv_state_3_LC_15_17_7  (
            .in0(N__11526),
            .in1(N__8262),
            .in2(N__7267),
            .in3(N__7264),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12112),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_4_LC_15_18_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_4_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_4_LC_15_18_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_0_4_LC_15_18_0  (
            .in0(N__9405),
            .in1(N__9513),
            .in2(N__7252),
            .in3(N__11396),
            .lcout(),
            .ltout(\DUT.uart_inst0.g3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_4_LC_15_18_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_4_LC_15_18_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_4_LC_15_18_1 .LUT_INIT=16'b0100100001011010;
    LogicCell40 \DUT.uart_inst0.tx_countdown_4_LC_15_18_1  (
            .in0(N__9335),
            .in1(N__12323),
            .in2(N__7255),
            .in3(N__9986),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12105),
            .ce(N__11844),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_4_2_LC_15_18_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_4_2_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_4_2_LC_15_18_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNO_4_2_LC_15_18_2  (
            .in0(N__9402),
            .in1(N__9333),
            .in2(_gnd_net_),
            .in3(N__9832),
            .lcout(\DUT.uart_inst0.un1_tx_bits_remaining_axbxc2_N_4L5_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_4_LC_15_18_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_4_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_4_LC_15_18_3 .LUT_INIT=16'b0000010100000101;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_1_4_LC_15_18_3  (
            .in0(N__9754),
            .in1(_gnd_net_),
            .in2(N__9850),
            .in3(_gnd_net_),
            .lcout(\DUT.uart_inst0.g3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_RNO_4_LC_15_18_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_RNO_4_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_out_RNO_4_LC_15_18_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_out_RNO_4_LC_15_18_4  (
            .in0(N__9403),
            .in1(N__9334),
            .in2(N__9463),
            .in3(N__9509),
            .lcout(\DUT.uart_inst0.g0_i_a4_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_3_3_LC_15_18_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_3_3_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_3_3_LC_15_18_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_3_3_LC_15_18_5  (
            .in0(N__9837),
            .in1(N__12322),
            .in2(N__9521),
            .in3(N__9461),
            .lcout(\DUT.uart_inst0.un1_m7_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_2_3_LC_15_18_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_2_3_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_2_3_LC_15_18_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_2_3_LC_15_18_6  (
            .in0(N__9404),
            .in1(N__9833),
            .in2(_gnd_net_),
            .in3(N__9753),
            .lcout(\DUT.uart_inst0.tx_countdown_0_c3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNIUUGK1_3_LC_15_19_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNIUUGK1_3_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNIUUGK1_3_LC_15_19_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNIUUGK1_3_LC_15_19_0  (
            .in0(N__9385),
            .in1(N__9831),
            .in2(N__9517),
            .in3(N__9740),
            .lcout(\DUT.uart_inst0.tx_countdown_0_c4_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_15_19_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_15_19_1 .LUT_INIT=16'b0010001011011101;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_0_3_LC_15_19_1  (
            .in0(N__11392),
            .in1(N__7342),
            .in2(_gnd_net_),
            .in3(N__9503),
            .lcout(\DUT.uart_inst0.tx_countdown_7_1_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_4_3_LC_15_19_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_4_3_LC_15_19_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_4_3_LC_15_19_2 .LUT_INIT=16'b0100000000010000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_4_3_LC_15_19_2  (
            .in0(N__9386),
            .in1(N__9741),
            .in2(N__12673),
            .in3(N__11393),
            .lcout(),
            .ltout(\DUT.uart_inst0.un1_tx_state_0_a4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_15_19_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_15_19_3 .LUT_INIT=16'b0100110011101100;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_1_3_LC_15_19_3  (
            .in0(N__7336),
            .in1(N__10288),
            .in2(N__7330),
            .in3(N__9343),
            .lcout(),
            .ltout(\DUT.uart_inst0.un1_tx_clk_divider_s1_sn_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_3_LC_15_19_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_3_LC_15_19_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_3_LC_15_19_4 .LUT_INIT=16'b1101000011011101;
    LogicCell40 \DUT.uart_inst0.tx_countdown_3_LC_15_19_4  (
            .in0(N__9966),
            .in1(N__12339),
            .in2(N__7327),
            .in3(N__7324),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12100),
            .ce(N__11848),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_1_LC_15_19_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_1_LC_15_19_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_1_LC_15_19_5 .LUT_INIT=16'b0000101011110101;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_0_1_LC_15_19_5  (
            .in0(N__11394),
            .in1(_gnd_net_),
            .in2(N__9764),
            .in3(N__9849),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_countdown_RNO_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_1_LC_15_19_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_1_LC_15_19_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_1_LC_15_19_6 .LUT_INIT=16'b0000111100000101;
    LogicCell40 \DUT.uart_inst0.tx_countdown_1_LC_15_19_6  (
            .in0(N__9965),
            .in1(_gnd_net_),
            .in2(N__7318),
            .in3(N__12338),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12100),
            .ce(N__11848),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_0_LC_15_19_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_0_LC_15_19_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_0_LC_15_19_7 .LUT_INIT=16'b0100100001011010;
    LogicCell40 \DUT.uart_inst0.tx_countdown_0_LC_15_19_7  (
            .in0(N__11395),
            .in1(N__12340),
            .in2(N__9765),
            .in3(N__9964),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12100),
            .ce(N__11848),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_4_LC_15_20_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_4_LC_15_20_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_4_LC_15_20_0 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \DUT.uart_inst0.tx_data_4_LC_15_20_0  (
            .in0(N__10896),
            .in1(N__7423),
            .in2(N__10075),
            .in3(N__9989),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12093),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_RNO_6_LC_15_20_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_RNO_6_LC_15_20_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_out_RNO_6_LC_15_20_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \DUT.uart_inst0.tx_out_RNO_6_LC_15_20_1  (
            .in0(N__9347),
            .in1(N__9505),
            .in2(N__9457),
            .in3(N__9399),
            .lcout(),
            .ltout(\DUT.uart_inst0.g0_i_o4_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_RNO_3_LC_15_20_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_RNO_3_LC_15_20_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_out_RNO_3_LC_15_20_2 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \DUT.uart_inst0.tx_out_RNO_3_LC_15_20_2  (
            .in0(N__12317),
            .in1(N__12662),
            .in2(N__7624),
            .in3(N__9842),
            .lcout(\DUT.uart_inst0.g0_i_o4_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIN79A_2_LC_15_20_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIN79A_2_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIN79A_2_LC_15_20_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNIN79A_2_LC_15_20_4  (
            .in0(N__7612),
            .in1(N__8683),
            .in2(N__7549),
            .in3(N__7473),
            .lcout(\DUT.fifo_tx_inst.rFifoData_awe3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_RNO_0_0_LC_15_20_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_RNO_0_0_LC_15_20_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_data_RNO_0_0_LC_15_20_7 .LUT_INIT=16'b1100010111000000;
    LogicCell40 \DUT.uart_inst0.tx_data_RNO_0_0_LC_15_20_7  (
            .in0(N__10026),
            .in1(N__8718),
            .in2(N__12675),
            .in3(N__7450),
            .lcout(\DUT.uart_inst0.tx_data_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_15_21_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_15_21_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_15_21_0 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNI33EC1_4_LC_15_21_0  (
            .in0(N__7444),
            .in1(N__9660),
            .in2(N__7675),
            .in3(N__7432),
            .lcout(),
            .ltout(\DUT.rFifoDatarx_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_RNO_0_4_LC_15_21_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_RNO_0_4_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_data_RNO_0_4_LC_15_21_1 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \DUT.uart_inst0.tx_data_RNO_0_4_LC_15_21_1  (
            .in0(N__12666),
            .in1(N__9007),
            .in2(N__7426),
            .in3(N__10030),
            .lcout(\DUT.uart_inst0.tx_data_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_15_21_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_15_21_3 .LUT_INIT=16'b0001000110101111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram0__RNI4U0H_6_LC_15_21_3  (
            .in0(N__9658),
            .in1(N__7417),
            .in2(N__7405),
            .in3(N__7391),
            .lcout(),
            .ltout(\DUT.fifo_tx_inst.rFifoData_ramout_3_ns_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_15_21_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_15_21_4 .LUT_INIT=16'b1100101000001111;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIBBEC1_6_LC_15_21_4  (
            .in0(N__7954),
            .in1(N__8836),
            .in2(N__7789),
            .in3(N__9659),
            .lcout(\DUT.rFifoDatarx_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_2_LC_15_21_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_2_LC_15_21_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_2_LC_15_21_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \DUT.uart_inst0.tx_data_2_LC_15_21_5  (
            .in0(N__7786),
            .in1(N__10904),
            .in2(N__8746),
            .in3(N__9993),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12088),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_2_LC_15_21_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_2_LC_15_21_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_2_LC_15_21_7 .LUT_INIT=16'b1110111011111111;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_0_2_LC_15_21_7  (
            .in0(N__9855),
            .in1(N__9771),
            .in2(_gnd_net_),
            .in3(N__11398),
            .lcout(\DUT.uart_inst0.N_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_15_22_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_15_22_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_15_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__0_LC_15_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8933),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12083),
            .ce(N__7903),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_15_22_1 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_15_22_1 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_15_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__1_LC_15_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8991),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12083),
            .ce(N__7903),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_15_22_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_15_22_2 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_15_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__2_LC_15_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7767),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12083),
            .ce(N__7903),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_15_22_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_15_22_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_15_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__3_LC_15_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10275),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12083),
            .ce(N__7903),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_15_22_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_15_22_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_15_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__4_LC_15_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7717),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12083),
            .ce(N__7903),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_15_22_5 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_15_22_5 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_15_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__5_LC_15_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7666),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12083),
            .ce(N__7903),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_15_22_6 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_15_22_6 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_15_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__6_LC_15_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8876),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12083),
            .ce(N__7903),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_15_22_7 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_15_22_7 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_15_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram3__7_LC_15_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7944),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12083),
            .ce(N__7903),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_RNO_0_7_LC_15_23_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_RNO_0_7_LC_15_23_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_data_RNO_0_7_LC_15_23_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \DUT.uart_inst0.tx_data_RNO_0_7_LC_15_23_3  (
            .in0(_gnd_net_),
            .in1(N__12672),
            .in2(_gnd_net_),
            .in3(N__7885),
            .lcout(\DUT.uart_inst0.tx_data_8_321_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.SUM_0_2_LC_16_10_3 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.SUM_0_2_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.SUM_0_2_LC_16_10_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \fifo_inst.ftdi_input_inst.SUM_0_2_LC_16_10_3  (
            .in0(N__7847),
            .in1(N__7868),
            .in2(_gnd_net_),
            .in3(N__7810),
            .lcout(),
            .ltout(G_152_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_2_LC_16_10_4 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_2_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_2_LC_16_10_4 .LUT_INIT=16'b0000000011100010;
    LogicCell40 \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_2_LC_16_10_4  (
            .in0(N__7869),
            .in1(N__7834),
            .in2(N__7879),
            .in3(N__12539),
            .lcout(G_151),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_1_LC_16_10_5 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_1_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_1_LC_16_10_5 .LUT_INIT=16'b0000011000001010;
    LogicCell40 \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_1_LC_16_10_5  (
            .in0(N__7848),
            .in1(N__7812),
            .in2(N__12541),
            .in3(N__7833),
            .lcout(G_150),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_0_LC_16_10_7 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_0_LC_16_10_7 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_0_LC_16_10_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.ftdi_input_inst.rRamWrAddr_latch_0_LC_16_10_7  (
            .in0(N__12535),
            .in1(N__7811),
            .in2(_gnd_net_),
            .in3(N__7832),
            .lcout(G_149),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_input_inst.oPacketAvail_latch_LC_16_11_0 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_input_inst.oPacketAvail_latch_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_input_inst.oPacketAvail_latch_LC_16_11_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_inst.ftdi_input_inst.oPacketAvail_latch_LC_16_11_0  (
            .in0(N__11920),
            .in1(N__9264),
            .in2(_gnd_net_),
            .in3(N__7795),
            .lcout(G_148),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNI237O_0_LC_16_13_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNI237O_0_LC_16_13_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNI237O_0_LC_16_13_6 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \DUT.uart_inst0.recv_state_RNI237O_0_LC_16_13_6  (
            .in0(N__8183),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8038),
            .lcout(\DUT.uart_inst0.N_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNI6B671_5_LC_16_14_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI6B671_5_LC_16_14_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI6B671_5_LC_16_14_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNI6B671_5_LC_16_14_1  (
            .in0(N__10397),
            .in1(N__10424),
            .in2(N__10372),
            .in3(N__10451),
            .lcout(\DUT.uart_inst0.un2_rx_clk_divider_a_10 ),
            .ltout(\DUT.uart_inst0.un2_rx_clk_divider_a_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIKU472_10_LC_16_14_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIKU472_10_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIKU472_10_LC_16_14_2 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIKU472_10_LC_16_14_2  (
            .in0(N__9030),
            .in1(_gnd_net_),
            .in2(N__8062),
            .in3(N__9045),
            .lcout(\DUT.uart_inst0.rx_clk_divider_RNIKU472Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_1_0_LC_16_14_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_1_0_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_1_0_LC_16_14_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_1_0_LC_16_14_6  (
            .in0(N__7965),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8013),
            .lcout(),
            .ltout(\DUT.uart_inst0.recv_state_RNO_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_0_LC_16_14_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_0_LC_16_14_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_0_LC_16_14_7 .LUT_INIT=16'b0101010101110101;
    LogicCell40 \DUT.uart_inst0.recv_state_0_LC_16_14_7  (
            .in0(N__8050),
            .in1(N__8426),
            .in2(N__8044),
            .in3(N__8370),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12133),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_1_LC_16_15_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_1_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_1_LC_16_15_0 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_0_1_LC_16_15_0  (
            .in0(N__8107),
            .in1(N__9128),
            .in2(N__8293),
            .in3(N__8545),
            .lcout(\DUT.uart_inst0.N_105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNI7H9R3_10_LC_16_15_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI7H9R3_10_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI7H9R3_10_LC_16_15_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNI7H9R3_10_LC_16_15_1  (
            .in0(N__8023),
            .in1(N__9046),
            .in2(N__9034),
            .in3(N__9192),
            .lcout(\DUT.uart_inst0.un2_rx_clk_divider_0 ),
            .ltout(\DUT.uart_inst0.un2_rx_clk_divider_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNI8UI86_3_LC_16_15_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNI8UI86_3_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNI8UI86_3_LC_16_15_2 .LUT_INIT=16'b1111010111000101;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNI8UI86_3_LC_16_15_2  (
            .in0(N__8485),
            .in1(N__8079),
            .in2(N__8017),
            .in3(N__8475),
            .lcout(\DUT.uart_inst0.rx_countdown_8_i_o2_1_2 ),
            .ltout(\DUT.uart_inst0.rx_countdown_8_i_o2_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_4_LC_16_15_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_4_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_4_LC_16_15_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_4_LC_16_15_3  (
            .in0(N__8291),
            .in1(N__8012),
            .in2(N__7975),
            .in3(N__8359),
            .lcout(),
            .ltout(\DUT.uart_inst0.recv_state_RNO_0Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_4_LC_16_15_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_4_LC_16_15_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.recv_state_4_LC_16_15_4 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \DUT.uart_inst0.recv_state_4_LC_16_15_4  (
            .in0(N__11531),
            .in1(N__7969),
            .in2(N__7972),
            .in3(N__8292),
            .lcout(\DUT.uart_inst0.recv_stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12129),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_3_LC_16_15_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_3_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNO_0_3_LC_16_15_6 .LUT_INIT=16'b0000000101000101;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNO_0_3_LC_16_15_6  (
            .in0(N__8288),
            .in1(N__9129),
            .in2(N__8512),
            .in3(N__8080),
            .lcout(\DUT.uart_inst0.N_102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.recv_state_RNO_0_5_LC_16_15_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.recv_state_RNO_0_5_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.recv_state_RNO_0_5_LC_16_15_7 .LUT_INIT=16'b0011011111110111;
    LogicCell40 \DUT.uart_inst0.recv_state_RNO_0_5_LC_16_15_7  (
            .in0(N__8263),
            .in1(N__11923),
            .in2(N__8240),
            .in3(N__8155),
            .lcout(\DUT.uart_inst0.recv_state_srsts_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_s1_c_LC_16_16_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_s1_c_LC_16_16_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_s1_c_LC_16_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_0_s1_c_LC_16_16_0  (
            .in0(_gnd_net_),
            .in1(N__9062),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_16_0_),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_0_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_s1_c_RNIKPDT_LC_16_16_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_s1_c_RNIKPDT_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_0_s1_c_RNIKPDT_LC_16_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_0_s1_c_RNIKPDT_LC_16_16_1  (
            .in0(_gnd_net_),
            .in1(N__12997),
            .in2(N__8544),
            .in3(N__8092),
            .lcout(\DUT.uart_inst0.rx_countdown_3_s1_1 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_countdown_3_cry_0_s1 ),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_s1_THRU_LUT4_0_LC_16_16_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_s1_THRU_LUT4_0_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_1_s1_THRU_LUT4_0_LC_16_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_1_s1_THRU_LUT4_0_LC_16_16_2  (
            .in0(_gnd_net_),
            .in1(N__13000),
            .in2(N__8313),
            .in3(N__8083),
            .lcout(\DUT.uart_inst0.rx_countdown_3_cry_1_s1_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_countdown_3_cry_1_s1 ),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_2_s1_c_RNIO52I_LC_16_16_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_2_s1_c_RNIO52I_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_2_s1_c_RNIO52I_LC_16_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_2_s1_c_RNIO52I_LC_16_16_3  (
            .in0(_gnd_net_),
            .in1(N__12998),
            .in2(N__8508),
            .in3(N__8071),
            .lcout(\DUT.uart_inst0.rx_countdown_3_s1_3 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_countdown_3_cry_2_s1 ),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_s1_c_RNIQBCS_LC_16_16_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_s1_c_RNIQBCS_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_3_s1_c_RNIQBCS_LC_16_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_3_s1_c_RNIQBCS_LC_16_16_4  (
            .in0(_gnd_net_),
            .in1(N__13001),
            .in2(N__8463),
            .in3(N__8068),
            .lcout(\DUT.uart_inst0.rx_countdown_3_s1_4 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_countdown_3_cry_3_s1 ),
            .carryout(\DUT.uart_inst0.rx_countdown_3_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_cry_4_s1_c_RNISHMM_LC_16_16_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_4_s1_c_RNISHMM_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_3_cry_4_s1_c_RNISHMM_LC_16_16_5 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_cry_4_s1_c_RNISHMM_LC_16_16_5  (
            .in0(N__9161),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8065),
            .lcout(\DUT.uart_inst0.rx_countdown_3_s1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_0_LC_16_16_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_0_LC_16_16_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_0_LC_16_16_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_0_LC_16_16_6  (
            .in0(N__12999),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11276),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12124),
            .ce(),
            .sr(N__12730));
    defparam \DUT.uart_inst0.rx_clk_divider_3_LC_16_17_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_3_LC_16_17_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_3_LC_16_17_0 .LUT_INIT=16'b1111111110110111;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_3_LC_16_17_0  (
            .in0(N__10501),
            .in1(N__11177),
            .in2(N__10530),
            .in3(N__9142),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12118),
            .ce(N__11845),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_1_LC_16_17_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_1_LC_16_17_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_1_LC_16_17_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \DUT.uart_inst0.rx_countdown_1_LC_16_17_2  (
            .in0(_gnd_net_),
            .in1(N__11175),
            .in2(_gnd_net_),
            .in3(N__8554),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12118),
            .ce(N__11845),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_3_LC_16_17_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_3_LC_16_17_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_3_LC_16_17_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \DUT.uart_inst0.rx_countdown_3_LC_16_17_3  (
            .in0(N__11176),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8521),
            .lcout(\DUT.uart_inst0.rx_countdownZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12118),
            .ce(N__11845),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_RNIFRQU_3_LC_16_17_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_RNIFRQU_3_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_countdown_RNIFRQU_3_LC_16_17_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \DUT.uart_inst0.rx_countdown_RNIFRQU_3_LC_16_17_4  (
            .in0(_gnd_net_),
            .in1(N__8459),
            .in2(_gnd_net_),
            .in3(N__8504),
            .lcout(\DUT.uart_inst0.rx_countdown_8_i_o2_1_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_4_LC_16_17_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_4_LC_16_17_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_4_LC_16_17_5 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \DUT.uart_inst0.rx_countdown_4_LC_16_17_5  (
            .in0(N__9143),
            .in1(N__9092),
            .in2(N__8464),
            .in3(N__8476),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12118),
            .ce(N__11845),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_2_LC_16_18_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_2_LC_16_18_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_2_LC_16_18_0 .LUT_INIT=16'b1111000011110001;
    LogicCell40 \DUT.uart_inst0.rx_countdown_2_LC_16_18_0  (
            .in0(N__8443),
            .in1(N__8430),
            .in2(N__8383),
            .in3(N__8371),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12113),
            .ce(N__11849),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_3_LC_16_18_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_3_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_3_LC_16_18_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_3_LC_16_18_1  (
            .in0(N__12435),
            .in1(N__12217),
            .in2(N__10333),
            .in3(N__12387),
            .lcout(\DUT.uart_inst0.N_159 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_1_2_LC_16_18_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_1_2_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_1_2_LC_16_18_2 .LUT_INIT=16'b0111110111111101;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNO_1_2_LC_16_18_2  (
            .in0(N__12388),
            .in1(N__8773),
            .in2(N__12676),
            .in3(N__8689),
            .lcout(\DUT.uart_inst0.tx_bits_remaining_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_RNIBPK2_0_LC_16_18_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNIBPK2_0_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNIBPK2_0_LC_16_18_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNIBPK2_0_LC_16_18_3  (
            .in0(_gnd_net_),
            .in1(N__11277),
            .in2(_gnd_net_),
            .in3(N__11257),
            .lcout(),
            .ltout(\DUT.uart_inst0.un1_tx_clk_divider_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_RNITC2S1_0_LC_16_18_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNITC2S1_0_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNITC2S1_0_LC_16_18_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNITC2S1_0_LC_16_18_4  (
            .in0(N__9529),
            .in1(N__9535),
            .in2(N__8701),
            .in3(N__9541),
            .lcout(\DUT.uart_inst0.un1_tx_clk_divider_0 ),
            .ltout(\DUT.uart_inst0.un1_tx_clk_divider_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_2_2_LC_16_18_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_2_2_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_2_2_LC_16_18_5 .LUT_INIT=16'b0010000000000010;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNO_2_2_LC_16_18_5  (
            .in0(N__8698),
            .in1(N__9885),
            .in2(N__8692),
            .in3(N__9755),
            .lcout(\DUT.uart_inst0.un1_tx_bits_remaining_axbxc2_N_4L5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIBPFM_1_LC_16_19_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIBPFM_1_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoCount_RNIBPFM_1_LC_16_19_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \DUT.fifo_tx_inst.rFifoCount_RNIBPFM_1_LC_16_19_0  (
            .in0(N__11602),
            .in1(N__8682),
            .in2(N__8629),
            .in3(N__8577),
            .lcout(\DUT.fifo_tx_inst.rFifoCount_RNIBPFMZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNI18BH1_5_LC_16_19_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNI18BH1_5_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNI18BH1_5_LC_16_19_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNI18BH1_5_LC_16_19_1  (
            .in0(N__9504),
            .in1(N__12654),
            .in2(N__9456),
            .in3(N__9838),
            .lcout(),
            .ltout(\DUT.uart_inst0.g0_0_0_a3_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNIP6303_4_LC_16_19_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNIP6303_4_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNIP6303_4_LC_16_19_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNIP6303_4_LC_16_19_2  (
            .in0(N__9339),
            .in1(N__8584),
            .in2(N__8590),
            .in3(N__9400),
            .lcout(),
            .ltout(\DUT.uart_inst0.g0_0_0_a3_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNI1BIT5_0_LC_16_19_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNI1BIT5_0_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNI1BIT5_0_LC_16_19_3 .LUT_INIT=16'b1110101010111010;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNI1BIT5_0_LC_16_19_3  (
            .in0(N__9682),
            .in1(N__9759),
            .in2(N__8587),
            .in3(N__11388),
            .lcout(\DUT.uart_inst0.N_152_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_0_3_LC_16_19_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_0_3_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_0_3_LC_16_19_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNI6CFK_0_3_LC_16_19_5  (
            .in0(N__12443),
            .in1(N__12216),
            .in2(N__10331),
            .in3(N__12389),
            .lcout(\DUT.uart_inst0.N_159_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.rTransmit_LC_16_19_6 .C_ON=1'b0;
    defparam \DUT.rTransmit_LC_16_19_6 .SEQ_MODE=4'b1000;
    defparam \DUT.rTransmit_LC_16_19_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DUT.rTransmit_LC_16_19_6  (
            .in0(N__12655),
            .in1(N__12324),
            .in2(_gnd_net_),
            .in3(N__8578),
            .lcout(\DUT.rTransmitZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12106),
            .ce(),
            .sr(N__12493));
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_5_LC_16_20_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_5_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_0_5_LC_16_20_0 .LUT_INIT=16'b1101001011110000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_0_5_LC_16_20_0  (
            .in0(N__11399),
            .in1(N__9348),
            .in2(N__9462),
            .in3(N__9291),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_countdown_0_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_5_LC_16_20_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_5_LC_16_20_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_5_LC_16_20_1 .LUT_INIT=16'b1010000011110000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_5_LC_16_20_1  (
            .in0(N__12328),
            .in1(_gnd_net_),
            .in2(N__8821),
            .in3(N__9968),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12101),
            .ce(N__11862),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_RNO_1_LC_16_20_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_RNO_1_LC_16_20_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_out_RNO_1_LC_16_20_5 .LUT_INIT=16'b0000101100001110;
    LogicCell40 \DUT.uart_inst0.tx_out_RNO_1_LC_16_20_5  (
            .in0(N__8818),
            .in1(N__11400),
            .in2(N__8796),
            .in3(N__9763),
            .lcout(),
            .ltout(\DUT.uart_inst0.N_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_LC_16_20_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_LC_16_20_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_out_LC_16_20_6 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \DUT.uart_inst0.tx_out_LC_16_20_6  (
            .in0(N__10294),
            .in1(N__12670),
            .in2(N__8812),
            .in3(N__9688),
            .lcout(P1A7_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12101),
            .ce(N__11862),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_2_LC_16_20_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_2_LC_16_20_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_countdown_2_LC_16_20_7 .LUT_INIT=16'b1010111001011101;
    LogicCell40 \DUT.uart_inst0.tx_countdown_2_LC_16_20_7  (
            .in0(N__8779),
            .in1(N__9967),
            .in2(N__12337),
            .in3(N__9401),
            .lcout(\DUT.uart_inst0.tx_countdownZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12101),
            .ce(N__11862),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_3_2_LC_16_21_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_3_2_LC_16_21_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_3_2_LC_16_21_1 .LUT_INIT=16'b0000001101000111;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNO_3_2_LC_16_21_1  (
            .in0(N__9451),
            .in1(N__12645),
            .in2(N__11623),
            .in3(N__9522),
            .lcout(\DUT.uart_inst0.un1_tx_bits_remaining_axbxc2_N_4L5_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_16_21_2 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_16_21_2 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_16_21_2 .LUT_INIT=16'b1011100000110011;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNINMDC1_1_LC_16_21_2  (
            .in0(N__8947),
            .in1(N__8764),
            .in2(N__8755),
            .in3(N__9676),
            .lcout(),
            .ltout(\DUT.rFifoDatarx_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_RNO_0_1_LC_16_21_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_RNO_0_1_LC_16_21_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_data_RNO_0_1_LC_16_21_3 .LUT_INIT=16'b1000100010111000;
    LogicCell40 \DUT.uart_inst0.tx_data_RNO_0_1_LC_16_21_3  (
            .in0(N__8739),
            .in1(N__12646),
            .in2(N__8728),
            .in3(N__10052),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_data_RNO_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_1_LC_16_21_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_1_LC_16_21_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_1_LC_16_21_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \DUT.uart_inst0.tx_data_1_LC_16_21_4  (
            .in0(N__9991),
            .in1(N__10900),
            .in2(N__8725),
            .in3(N__8722),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12094),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_0_LC_16_21_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_0_LC_16_21_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_0_LC_16_21_5 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \DUT.uart_inst0.tx_data_0_LC_16_21_5  (
            .in0(N__9870),
            .in1(N__8707),
            .in2(N__10906),
            .in3(N__9990),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12094),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_RNO_0_5_LC_16_21_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_RNO_0_5_LC_16_21_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_data_RNO_0_5_LC_16_21_6 .LUT_INIT=16'b1100010111000000;
    LogicCell40 \DUT.uart_inst0.tx_data_RNO_0_5_LC_16_21_6  (
            .in0(N__10053),
            .in1(N__10093),
            .in2(N__12671),
            .in3(N__9019),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_data_RNO_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_5_LC_16_21_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_5_LC_16_21_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_5_LC_16_21_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \DUT.uart_inst0.tx_data_5_LC_16_21_7  (
            .in0(N__10899),
            .in1(N__9006),
            .in2(N__9010),
            .in3(N__9992),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12094),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_16_22_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_16_22_0 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_16_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__1_LC_16_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8992),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12089),
            .ce(N__10237),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_16_22_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_16_22_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_16_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__0_LC_16_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8938),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12089),
            .ce(N__10237),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_16_22_4 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_16_22_4 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_16_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__6_LC_16_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8877),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12089),
            .ce(N__10237),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_7_LC_16_23_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_7_LC_16_23_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_7_LC_16_23_0 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \DUT.uart_inst0.tx_data_7_LC_16_23_0  (
            .in0(N__10905),
            .in1(N__8827),
            .in2(N__10116),
            .in3(N__10054),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12084),
            .ce(N__9997),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_0_LC_17_13_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_0_LC_17_13_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_0_LC_17_13_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_0_LC_17_13_0  (
            .in0(_gnd_net_),
            .in1(N__11145),
            .in2(_gnd_net_),
            .in3(N__10152),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12138),
            .ce(N__11832),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_6_LC_17_13_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_6_LC_17_13_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_6_LC_17_13_1 .LUT_INIT=16'b1111111110011111;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_6_LC_17_13_1  (
            .in0(N__10408),
            .in1(N__10426),
            .in2(N__11179),
            .in3(N__9145),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12138),
            .ce(N__11832),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_7_LC_17_13_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_7_LC_17_13_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_7_LC_17_13_4 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_7_LC_17_13_4  (
            .in0(N__10399),
            .in1(N__10381),
            .in2(_gnd_net_),
            .in3(N__11146),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12138),
            .ce(N__11832),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_5_LC_17_13_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_5_LC_17_13_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_5_LC_17_13_5 .LUT_INIT=16'b1111111110011111;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_5_LC_17_13_5  (
            .in0(N__10435),
            .in1(N__10453),
            .in2(N__11178),
            .in3(N__9144),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12138),
            .ce(N__11832),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIB99J_10_LC_17_14_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIB99J_10_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIB99J_10_LC_17_14_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIB99J_10_LC_17_14_0  (
            .in0(N__10796),
            .in1(N__10769),
            .in2(N__10723),
            .in3(N__10745),
            .lcout(\DUT.uart_inst0.un2_rx_clk_divider_a_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_9_LC_17_14_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_9_LC_17_14_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_9_LC_17_14_1 .LUT_INIT=16'b1000100001000100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_9_LC_17_14_1  (
            .in0(N__10798),
            .in1(N__11163),
            .in2(_gnd_net_),
            .in3(N__10780),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12136),
            .ce(N__11836),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_10_LC_17_14_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_10_LC_17_14_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_10_LC_17_14_2 .LUT_INIT=16'b1010000001010000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_10_LC_17_14_2  (
            .in0(N__10756),
            .in1(_gnd_net_),
            .in2(N__11180),
            .in3(N__10770),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12136),
            .ce(N__11836),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_11_LC_17_14_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_11_LC_17_14_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_11_LC_17_14_3 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_11_LC_17_14_3  (
            .in0(N__10746),
            .in1(N__10732),
            .in2(_gnd_net_),
            .in3(N__11156),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12136),
            .ce(N__11836),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_12_LC_17_14_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_12_LC_17_14_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_12_LC_17_14_4 .LUT_INIT=16'b1010000001010000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_12_LC_17_14_4  (
            .in0(N__10721),
            .in1(_gnd_net_),
            .in2(N__11181),
            .in3(N__10705),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12136),
            .ce(N__11836),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_LC_17_14_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_1_LC_17_14_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_LC_17_14_5 .LUT_INIT=16'b1000100001000100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_LC_17_14_5  (
            .in0(N__10570),
            .in1(N__11161),
            .in2(_gnd_net_),
            .in3(N__10588),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12136),
            .ce(N__11836),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_16_LC_17_14_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_16_LC_17_14_6 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_16_LC_17_14_6 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_16_LC_17_14_6  (
            .in0(N__11160),
            .in1(N__10597),
            .in2(_gnd_net_),
            .in3(N__10615),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12136),
            .ce(N__11836),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_4_LC_17_14_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_4_LC_17_14_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_4_LC_17_14_7 .LUT_INIT=16'b1000100001000100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_4_LC_17_14_7  (
            .in0(N__10462),
            .in1(N__11162),
            .in2(_gnd_net_),
            .in3(N__10484),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12136),
            .ce(N__11836),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNI3ALC_17_LC_17_15_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI3ALC_17_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNI3ALC_17_LC_17_15_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNI3ALC_17_LC_17_15_0  (
            .in0(N__10667),
            .in1(N__10694),
            .in2(N__11083),
            .in3(N__10640),
            .lcout(\DUT.uart_inst0.un2_rx_clk_divider_a_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_13_LC_17_15_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_13_LC_17_15_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_13_LC_17_15_1 .LUT_INIT=16'b1010010100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_13_LC_17_15_1  (
            .in0(N__10695),
            .in1(_gnd_net_),
            .in2(N__10681),
            .in3(N__11196),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12134),
            .ce(N__11843),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_14_LC_17_15_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_14_LC_17_15_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_14_LC_17_15_2 .LUT_INIT=16'b1010000001010000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_14_LC_17_15_2  (
            .in0(N__10651),
            .in1(_gnd_net_),
            .in2(N__11203),
            .in3(N__10669),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12134),
            .ce(N__11843),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_15_LC_17_15_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_15_LC_17_15_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_15_LC_17_15_3 .LUT_INIT=16'b1010010100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_15_LC_17_15_3  (
            .in0(N__10641),
            .in1(_gnd_net_),
            .in2(N__10627),
            .in3(N__11200),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12134),
            .ce(N__11843),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIIDCT_2_LC_17_15_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIIDCT_2_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIIDCT_2_LC_17_15_4 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIIDCT_2_LC_17_15_4  (
            .in0(_gnd_net_),
            .in1(N__10556),
            .in2(N__10485),
            .in3(N__10526),
            .lcout(),
            .ltout(\DUT.uart_inst0.un2_rx_clk_divider_a_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_RNIJI4K1_16_LC_17_15_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIJI4K1_16_LC_17_15_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_RNIJI4K1_16_LC_17_15_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_RNIJI4K1_16_LC_17_15_5  (
            .in0(N__10613),
            .in1(N__10153),
            .in2(N__9199),
            .in3(N__10586),
            .lcout(\DUT.uart_inst0.un2_rx_clk_divider_a_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_2_LC_17_15_7 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_2_LC_17_15_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_2_LC_17_15_7 .LUT_INIT=16'b1001100100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_2_LC_17_15_7  (
            .in0(N__10557),
            .in1(N__10543),
            .in2(_gnd_net_),
            .in3(N__11201),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12134),
            .ce(N__11843),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_5_LC_17_16_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_5_LC_17_16_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_5_LC_17_16_0 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \DUT.uart_inst0.rx_countdown_5_LC_17_16_0  (
            .in0(N__9165),
            .in1(N__9131),
            .in2(N__9097),
            .in3(N__9181),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12130),
            .ce(N__11846),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_countdown_0_LC_17_16_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_countdown_0_LC_17_16_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_countdown_0_LC_17_16_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \DUT.uart_inst0.rx_countdown_0_LC_17_16_1  (
            .in0(N__9130),
            .in1(N__9093),
            .in2(_gnd_net_),
            .in3(N__9068),
            .lcout(\DUT.uart_inst0.rx_countdownZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12130),
            .ce(N__11846),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_8_LC_17_16_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_8_LC_17_16_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_8_LC_17_16_3 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_8_LC_17_16_3  (
            .in0(N__11174),
            .in1(N__10345),
            .in2(_gnd_net_),
            .in3(N__10367),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12130),
            .ce(N__11846),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rRxF_n_1_LC_17_16_6 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rRxF_n_1_LC_17_16_6 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rRxF_n_1_LC_17_16_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \fifo_inst.ftdi_output_inst.rRxF_n_1_LC_17_16_6  (
            .in0(N__12165),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\fifo_inst.ftdi_output_inst.rRxF_nZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12130),
            .ce(N__11846),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rTxE_n_RNIJBK2_1_LC_17_17_0 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rTxE_n_RNIJBK2_1_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_output_inst.rTxE_n_RNIJBK2_1_LC_17_17_0 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \fifo_inst.ftdi_output_inst.rTxE_n_RNIJBK2_1_LC_17_17_0  (
            .in0(N__9271),
            .in1(N__10195),
            .in2(_gnd_net_),
            .in3(N__10171),
            .lcout(\fifo_inst.ftdi_output_inst.N_86_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_2_LC_17_17_2 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_2_LC_17_17_2 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_2_LC_17_17_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_2_LC_17_17_2  (
            .in0(N__11930),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11292),
            .lcout(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12125),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rRxF_n_RNIHPJ8_1_LC_17_17_3 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rRxF_n_RNIHPJ8_1_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_output_inst.rRxF_n_RNIHPJ8_1_LC_17_17_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rRxF_n_RNIHPJ8_1_LC_17_17_3  (
            .in0(N__12164),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11307),
            .lcout(\fifo_inst.ftdi_output_inst.N_95 ),
            .ltout(\fifo_inst.ftdi_output_inst.N_95_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_3_LC_17_17_4 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_3_LC_17_17_4 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_3_LC_17_17_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_3_LC_17_17_4  (
            .in0(N__9208),
            .in1(N__11935),
            .in2(N__9253),
            .in3(N__11329),
            .lcout(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12125),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_4_LC_17_17_5 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_4_LC_17_17_5 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_4_LC_17_17_5 .LUT_INIT=16'b1100110001000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_4_LC_17_17_5  (
            .in0(N__11012),
            .in1(N__11931),
            .in2(N__11043),
            .in3(N__9249),
            .lcout(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12125),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNO_0_0_LC_17_17_6 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNO_0_0_LC_17_17_6 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNO_0_0_LC_17_17_6 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_RNO_0_0_LC_17_17_6  (
            .in0(N__9228),
            .in1(N__11036),
            .in2(N__11941),
            .in3(N__11011),
            .lcout(),
            .ltout(\fifo_inst.ftdi_output_inst.m14_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_0_LC_17_17_7 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_0_LC_17_17_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_0_LC_17_17_7 .LUT_INIT=16'b0000111110001111;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_0_LC_17_17_7  (
            .in0(N__11328),
            .in1(N__9217),
            .in2(N__9211),
            .in3(N__9207),
            .lcout(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12125),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_1_LC_17_18_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_1_LC_17_18_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_bits_remaining_1_LC_17_18_0 .LUT_INIT=16'b1111011100001000;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_1_LC_17_18_0  (
            .in0(N__9983),
            .in1(N__10871),
            .in2(N__12405),
            .in3(N__12224),
            .lcout(\DUT.uart_inst0.tx_bits_remainingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12119),
            .ce(),
            .sr(N__11632));
    defparam \DUT.uart_inst0.tx_bits_remaining_0_LC_17_18_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_0_LC_17_18_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_bits_remaining_0_LC_17_18_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_0_LC_17_18_1  (
            .in0(N__10869),
            .in1(N__12396),
            .in2(_gnd_net_),
            .in3(N__9982),
            .lcout(\DUT.uart_inst0.tx_bits_remainingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12119),
            .ce(),
            .sr(N__11632));
    defparam \DUT.uart_inst0.tx_bits_remaining_3_LC_17_18_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_3_LC_17_18_2 .SEQ_MODE=4'b1001;
    defparam \DUT.uart_inst0.tx_bits_remaining_3_LC_17_18_2 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_3_LC_17_18_2  (
            .in0(N__9985),
            .in1(N__10870),
            .in2(N__12352),
            .in3(N__10327),
            .lcout(\DUT.uart_inst0.tx_bits_remainingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12119),
            .ce(),
            .sr(N__11632));
    defparam \DUT.uart_inst0.tx_bits_remaining_2_LC_17_18_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_2_LC_17_18_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_bits_remaining_2_LC_17_18_3 .LUT_INIT=16'b0110101010011010;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_2_LC_17_18_3  (
            .in0(N__12442),
            .in1(N__9984),
            .in2(N__12190),
            .in3(N__9547),
            .lcout(\DUT.uart_inst0.tx_bits_remainingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12119),
            .ce(),
            .sr(N__11632));
    defparam \DUT.uart_inst0.tx_clk_divider_RNI2V95_2_LC_17_19_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI2V95_2_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI2V95_2_LC_17_19_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNI2V95_2_LC_17_19_0  (
            .in0(N__11739),
            .in1(N__11758),
            .in2(N__11236),
            .in3(N__11217),
            .lcout(\DUT.uart_inst0.un1_tx_clk_divider_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_13_LC_17_19_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_13_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_13_LC_17_19_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_13_LC_17_19_1  (
            .in0(N__12762),
            .in1(N__11724),
            .in2(N__12745),
            .in3(N__11709),
            .lcout(\DUT.uart_inst0.un1_tx_clk_divider_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_8_LC_17_19_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_8_LC_17_19_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_8_LC_17_19_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_RNI8Q1Q_8_LC_17_19_2  (
            .in0(N__11694),
            .in1(N__11679),
            .in2(N__11650),
            .in3(N__11664),
            .lcout(\DUT.uart_inst0.un1_tx_clk_divider_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNIJ3F33_3_LC_17_19_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNIJ3F33_3_LC_17_19_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNIJ3F33_3_LC_17_19_3 .LUT_INIT=16'b0000011000000011;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNIJ3F33_3_LC_17_19_3  (
            .in0(N__9767),
            .in1(N__9851),
            .in2(N__9523),
            .in3(N__11376),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_data_i_m_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNIHJJ88_5_LC_17_19_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNIHJJ88_5_LC_17_19_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNIHJJ88_5_LC_17_19_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNIHJJ88_5_LC_17_19_4  (
            .in0(N__9452),
            .in1(N__9409),
            .in2(N__9352),
            .in3(N__9277),
            .lcout(\DUT.uart_inst0.N_345_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNIBSRA4_4_LC_17_19_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNIBSRA4_4_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNIBSRA4_4_LC_17_19_5 .LUT_INIT=16'b0111110111101110;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNIBSRA4_4_LC_17_19_5  (
            .in0(N__9766),
            .in1(N__9349),
            .in2(N__9295),
            .in3(N__11375),
            .lcout(\DUT.uart_inst0.tx_state_ns_0_o3_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_RNO_0_6_LC_17_20_0 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_RNO_0_6_LC_17_20_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_data_RNO_0_6_LC_17_20_0 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \DUT.uart_inst0.tx_data_RNO_0_6_LC_17_20_0  (
            .in0(N__12619),
            .in1(N__10132),
            .in2(N__10120),
            .in3(N__10043),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_data_RNO_0Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_6_LC_17_20_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_6_LC_17_20_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_6_LC_17_20_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \DUT.uart_inst0.tx_data_6_LC_17_20_1  (
            .in0(N__10898),
            .in1(N__10089),
            .in2(N__10096),
            .in3(N__9988),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12107),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_RNO_0_3_LC_17_20_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_RNO_0_3_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_data_RNO_0_3_LC_17_20_2 .LUT_INIT=16'b1010000011100100;
    LogicCell40 \DUT.uart_inst0.tx_data_RNO_0_3_LC_17_20_2  (
            .in0(N__12618),
            .in1(N__9553),
            .in2(N__10074),
            .in3(N__10042),
            .lcout(),
            .ltout(\DUT.uart_inst0.tx_data_RNO_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_data_3_LC_17_20_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_data_3_LC_17_20_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_data_3_LC_17_20_3 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \DUT.uart_inst0.tx_data_3_LC_17_20_3  (
            .in0(N__10897),
            .in1(N__9903),
            .in2(N__10000),
            .in3(N__9987),
            .lcout(\DUT.uart_inst0.tx_dataZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12107),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_RNO_5_LC_17_20_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_RNO_5_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_out_RNO_5_LC_17_20_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \DUT.uart_inst0.tx_out_RNO_5_LC_17_20_4  (
            .in0(N__12617),
            .in1(N__9889),
            .in2(N__9874),
            .in3(N__9856),
            .lcout(),
            .ltout(\DUT.uart_inst0.g0_i_a4_0_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_RNO_2_LC_17_20_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_RNO_2_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_out_RNO_2_LC_17_20_5 .LUT_INIT=16'b1000000000100000;
    LogicCell40 \DUT.uart_inst0.tx_out_RNO_2_LC_17_20_5  (
            .in0(N__9784),
            .in1(N__9772),
            .in2(N__9691),
            .in3(N__11401),
            .lcout(\DUT.uart_inst0.N_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNI5H8K_0_LC_17_20_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNI5H8K_0_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNI5H8K_0_LC_17_20_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \DUT.uart_inst0.tx_state_RNI5H8K_0_LC_17_20_6  (
            .in0(_gnd_net_),
            .in1(N__11586),
            .in2(_gnd_net_),
            .in3(N__12591),
            .lcout(\DUT.uart_inst0.N_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_17_21_0 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_17_21_0 .SEQ_MODE=4'b0000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_17_21_0 .LUT_INIT=16'b1000100011110011;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__RNIVUDC1_3_LC_17_21_0  (
            .in0(N__10246),
            .in1(N__9675),
            .in2(N__9577),
            .in3(N__9562),
            .lcout(\DUT.rFifoDatarx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNIB46K_3_LC_17_21_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNIB46K_3_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNIB46K_3_LC_17_21_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNIB46K_3_LC_17_21_1  (
            .in0(N__12614),
            .in1(N__10332),
            .in2(_gnd_net_),
            .in3(N__12444),
            .lcout(\DUT.uart_inst0.tx_state_ns_i_i_a2_0_0_0 ),
            .ltout(\DUT.uart_inst0.tx_state_ns_i_i_a2_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNICODU_1_LC_17_21_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNICODU_1_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNICODU_1_LC_17_21_2 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNICODU_1_LC_17_21_2  (
            .in0(_gnd_net_),
            .in1(N__12235),
            .in2(N__10297),
            .in3(N__12404),
            .lcout(\DUT.uart_inst0.tx_state_ns_i_i_a2_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_RNO_0_0_LC_17_21_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_RNO_0_0_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_RNO_0_0_LC_17_21_4 .LUT_INIT=16'b1010101010111011;
    LogicCell40 \DUT.uart_inst0.tx_state_RNO_0_0_LC_17_21_4  (
            .in0(N__12320),
            .in1(N__11610),
            .in2(_gnd_net_),
            .in3(N__12616),
            .lcout(\DUT.uart_inst0.tx_state_ns_i_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_out_RNO_0_LC_17_21_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_out_RNO_0_LC_17_21_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_out_RNO_0_LC_17_21_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \DUT.uart_inst0.tx_out_RNO_0_LC_17_21_5  (
            .in0(N__11609),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12319),
            .lcout(\DUT.uart_inst0.g0_i_a4_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_countdown_RNO_5_3_LC_17_21_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_countdown_RNO_5_3_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_countdown_RNO_5_3_LC_17_21_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \DUT.uart_inst0.tx_countdown_RNO_5_3_LC_17_21_6  (
            .in0(N__12318),
            .in1(N__11608),
            .in2(_gnd_net_),
            .in3(N__12615),
            .lcout(\DUT.uart_inst0.d_N_5_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_17_22_3 .C_ON=1'b0;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_17_22_3 .SEQ_MODE=4'b1000;
    defparam \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_17_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.fifo_tx_inst.rFifoData_rFifoData_ram2__3_LC_17_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10276),
            .lcout(\DUT.fifo_tx_inst.rFifoData_ram2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12095),
            .ce(N__10233),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rTxE_n_1_LC_17_23_6 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rTxE_n_1_LC_17_23_6 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rTxE_n_1_LC_17_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rTxE_n_1_LC_17_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10167),
            .lcout(\fifo_inst.ftdi_output_inst.rTxE_nZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12090),
            .ce(N__11866),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rTxE_n_0_LC_17_24_3 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rTxE_n_0_LC_17_24_3 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rTxE_n_0_LC_17_24_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \fifo_inst.ftdi_output_inst.rTxE_n_0_LC_17_24_3  (
            .in0(N__10183),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\fifo_inst.ftdi_output_inst.rTxE_nZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12085),
            .ce(N__11867),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_18_13_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_18_13_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_18_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_0_c_LC_18_13_0  (
            .in0(_gnd_net_),
            .in1(N__10151),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_13_0_),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_18_13_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_18_13_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_18_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_LUT4_0_LC_18_13_1  (
            .in0(_gnd_net_),
            .in1(N__10587),
            .in2(N__12991),
            .in3(N__10564),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_0 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_18_13_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_18_13_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_18_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_LUT4_0_LC_18_13_2  (
            .in0(_gnd_net_),
            .in1(N__10561),
            .in2(N__12995),
            .in3(N__10534),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_1 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_2_THRU_LUT4_0_LC_18_13_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_2_THRU_LUT4_0_LC_18_13_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_2_THRU_LUT4_0_LC_18_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_2_THRU_LUT4_0_LC_18_13_3  (
            .in0(_gnd_net_),
            .in1(N__10531),
            .in2(N__12992),
            .in3(N__10489),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_2 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_18_13_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_18_13_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_18_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_LUT4_0_LC_18_13_4  (
            .in0(_gnd_net_),
            .in1(N__12947),
            .in2(N__10486),
            .in3(N__10456),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_3 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_4_THRU_LUT4_0_LC_18_13_5 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_4_THRU_LUT4_0_LC_18_13_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_4_THRU_LUT4_0_LC_18_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_4_THRU_LUT4_0_LC_18_13_5  (
            .in0(_gnd_net_),
            .in1(N__10452),
            .in2(N__12993),
            .in3(N__10429),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_4 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_5_THRU_LUT4_0_LC_18_13_6 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_5_THRU_LUT4_0_LC_18_13_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_5_THRU_LUT4_0_LC_18_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_5_THRU_LUT4_0_LC_18_13_6  (
            .in0(_gnd_net_),
            .in1(N__10425),
            .in2(N__12996),
            .in3(N__10402),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_5 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_18_13_7 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_18_13_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_18_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_LUT4_0_LC_18_13_7  (
            .in0(_gnd_net_),
            .in1(N__10398),
            .in2(N__12994),
            .in3(N__10375),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_6 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_18_14_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_18_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_LUT4_0_LC_18_14_0  (
            .in0(_gnd_net_),
            .in1(N__10371),
            .in2(N__12989),
            .in3(N__10336),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_18_14_0_),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_18_14_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_18_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_LUT4_0_LC_18_14_1  (
            .in0(_gnd_net_),
            .in1(N__10797),
            .in2(N__12986),
            .in3(N__10774),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_8 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_LUT4_0_LC_18_14_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_LUT4_0_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_LUT4_0_LC_18_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_LUT4_0_LC_18_14_2  (
            .in0(_gnd_net_),
            .in1(N__10771),
            .in2(N__12990),
            .in3(N__10750),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_9 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_LUT4_0_LC_18_14_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_LUT4_0_LC_18_14_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_LUT4_0_LC_18_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_LUT4_0_LC_18_14_3  (
            .in0(_gnd_net_),
            .in1(N__10747),
            .in2(N__12983),
            .in3(N__10726),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_10 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_LUT4_0_LC_18_14_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_LUT4_0_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_LUT4_0_LC_18_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_LUT4_0_LC_18_14_4  (
            .in0(_gnd_net_),
            .in1(N__10722),
            .in2(N__12987),
            .in3(N__10699),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_11_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_11 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_LUT4_0_LC_18_14_5 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_LUT4_0_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_LUT4_0_LC_18_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_LUT4_0_LC_18_14_5  (
            .in0(_gnd_net_),
            .in1(N__10696),
            .in2(N__12984),
            .in3(N__10672),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_12 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_LUT4_0_LC_18_14_6 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_LUT4_0_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_LUT4_0_LC_18_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_LUT4_0_LC_18_14_6  (
            .in0(_gnd_net_),
            .in1(N__10668),
            .in2(N__12988),
            .in3(N__10645),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_13_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_13 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_LUT4_0_LC_18_14_7 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_LUT4_0_LC_18_14_7 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_LUT4_0_LC_18_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_LUT4_0_LC_18_14_7  (
            .in0(_gnd_net_),
            .in1(N__10642),
            .in2(N__12985),
            .in3(N__10618),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_14_THRU_CO ),
            .ltout(),
            .carryin(\DUT.uart_inst0.rx_clk_divider_1_cry_14 ),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_LUT4_0_LC_18_15_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_LUT4_0_LC_18_15_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_LUT4_0_LC_18_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_LUT4_0_LC_18_15_0  (
            .in0(_gnd_net_),
            .in1(N__10614),
            .in2(N__12982),
            .in3(N__10591),
            .lcout(\DUT.uart_inst0.rx_clk_divider_1_cry_15_THRU_CO ),
            .ltout(),
            .carryin(bfn_18_15_0_),
            .carryout(\DUT.uart_inst0.rx_clk_divider_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.rx_clk_divider_17_LC_18_15_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.rx_clk_divider_17_LC_18_15_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.rx_clk_divider_17_LC_18_15_1 .LUT_INIT=16'b1000100001000100;
    LogicCell40 \DUT.uart_inst0.rx_clk_divider_17_LC_18_15_1  (
            .in0(N__11082),
            .in1(N__11202),
            .in2(_gnd_net_),
            .in3(N__11086),
            .lcout(\DUT.uart_inst0.rx_clk_dividerZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12137),
            .ce(N__11847),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.oRamRdAddr_0_LC_18_16_0 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.oRamRdAddr_0_LC_18_16_0 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.oRamRdAddr_0_LC_18_16_0 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \fifo_inst.ftdi_output_inst.oRamRdAddr_0_LC_18_16_0  (
            .in0(N__10963),
            .in1(N__11035),
            .in2(N__11940),
            .in3(N__11014),
            .lcout(\fifo_inst.wRamRdAddr_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12135),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.oRamRdAddr_2_LC_18_16_1 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.oRamRdAddr_2_LC_18_16_1 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.oRamRdAddr_2_LC_18_16_1 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \fifo_inst.ftdi_output_inst.oRamRdAddr_2_LC_18_16_1  (
            .in0(N__10931),
            .in1(N__10965),
            .in2(N__11061),
            .in3(N__10981),
            .lcout(\fifo_inst.wRamRdAddr_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12135),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIBT9K_4_LC_18_16_6 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIBT9K_4_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_RNIBT9K_4_LC_18_16_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_RNIBT9K_4_LC_18_16_6  (
            .in0(N__11929),
            .in1(N__11034),
            .in2(_gnd_net_),
            .in3(N__11013),
            .lcout(\fifo_inst.ftdi_output_inst.N_3_0 ),
            .ltout(\fifo_inst.ftdi_output_inst.N_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.oRamRdAddr_1_LC_18_16_7 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.oRamRdAddr_1_LC_18_16_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.oRamRdAddr_1_LC_18_16_7 .LUT_INIT=16'b0110101001101010;
    LogicCell40 \fifo_inst.ftdi_output_inst.oRamRdAddr_1_LC_18_16_7  (
            .in0(N__10932),
            .in1(N__10964),
            .in2(N__10948),
            .in3(_gnd_net_),
            .lcout(\fifo_inst.wRamRdAddr_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12135),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_esr_1_LC_18_17_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_esr_1_LC_18_17_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_state_esr_1_LC_18_17_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \DUT.uart_inst0.tx_state_esr_1_LC_18_17_2  (
            .in0(N__10918),
            .in1(N__12223),
            .in2(_gnd_net_),
            .in3(N__12400),
            .lcout(\DUT.tx_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12131),
            .ce(N__10804),
            .sr(N__12495));
    defparam CONSTANT_ONE_LUT4_LC_18_18_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_18_18_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_18_18_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_18_18_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_esr_RNICLU7_1_LC_18_18_1 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_esr_RNICLU7_1_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_esr_RNICLU7_1_LC_18_18_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \DUT.uart_inst0.tx_state_esr_RNICLU7_1_LC_18_18_1  (
            .in0(_gnd_net_),
            .in1(N__11936),
            .in2(_gnd_net_),
            .in3(N__12266),
            .lcout(\DUT.uart_inst0.tx_state_0_sqmuxa_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_esr_RNO_1_LC_18_18_2 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_esr_RNO_1_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_esr_RNO_1_LC_18_18_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DUT.uart_inst0.tx_state_esr_RNO_1_LC_18_18_2  (
            .in0(_gnd_net_),
            .in1(N__10831),
            .in2(_gnd_net_),
            .in3(N__12693),
            .lcout(\DUT.uart_inst0.N_345_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_esr_RNIH67S_1_LC_18_18_3 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_esr_RNIH67S_1_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_esr_RNIH67S_1_LC_18_18_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \DUT.uart_inst0.tx_state_esr_RNIH67S_1_LC_18_18_3  (
            .in0(_gnd_net_),
            .in1(N__11937),
            .in2(_gnd_net_),
            .in3(N__11542),
            .lcout(\DUT.uart_inst0.tx_bits_remaining_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_esr_RNILOSP_1_LC_18_18_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_esr_RNILOSP_1_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_esr_RNILOSP_1_LC_18_18_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \DUT.uart_inst0.tx_state_esr_RNILOSP_1_LC_18_18_4  (
            .in0(N__12265),
            .in1(N__11622),
            .in2(_gnd_net_),
            .in3(N__12653),
            .lcout(\DUT.uart_inst0.tx_clk_divider_0_sqmuxa ),
            .ltout(\DUT.uart_inst0.tx_clk_divider_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_state_esr_RNIEJ9O2_1_LC_18_18_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_esr_RNIEJ9O2_1_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_state_esr_RNIEJ9O2_1_LC_18_18_5 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \DUT.uart_inst0.tx_state_esr_RNIEJ9O2_1_LC_18_18_5  (
            .in0(N__11494),
            .in1(_gnd_net_),
            .in2(N__11404),
            .in3(N__11397),
            .lcout(\DUT.uart_inst0.tx_clk_divider_1_sqmuxa_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rFifoState_1_LC_18_18_7 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_1_LC_18_18_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rFifoState_1_LC_18_18_7 .LUT_INIT=16'b0010101000000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rFifoState_1_LC_18_18_7  (
            .in0(N__11322),
            .in1(N__11311),
            .in2(N__12166),
            .in3(N__11938),
            .lcout(\fifo_inst.ftdi_output_inst.rFifoStateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12126),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_18_19_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_18_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_cry_c_0_LC_18_19_0  (
            .in0(_gnd_net_),
            .in1(N__11281),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_19_0_),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_clk_divider_1_LC_18_19_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_1_LC_18_19_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_1_LC_18_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_1_LC_18_19_1  (
            .in0(_gnd_net_),
            .in1(N__11253),
            .in2(N__12892),
            .in3(N__11239),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_1 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_0 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_1 ),
            .clk(N__12120),
            .ce(),
            .sr(N__12716));
    defparam \DUT.uart_inst0.tx_clk_divider_2_LC_18_19_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_2_LC_18_19_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_2_LC_18_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_2_LC_18_19_2  (
            .in0(_gnd_net_),
            .in1(N__11235),
            .in2(N__12896),
            .in3(N__11221),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_2 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_1 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_2 ),
            .clk(N__12120),
            .ce(),
            .sr(N__12716));
    defparam \DUT.uart_inst0.tx_clk_divider_3_LC_18_19_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_3_LC_18_19_3 .SEQ_MODE=4'b1001;
    defparam \DUT.uart_inst0.tx_clk_divider_3_LC_18_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_3_LC_18_19_3  (
            .in0(_gnd_net_),
            .in1(N__11218),
            .in2(N__12893),
            .in3(N__11206),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_3 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_2 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_3 ),
            .clk(N__12120),
            .ce(),
            .sr(N__12716));
    defparam \DUT.uart_inst0.tx_clk_divider_4_LC_18_19_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_4_LC_18_19_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_4_LC_18_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_4_LC_18_19_4  (
            .in0(_gnd_net_),
            .in1(N__11757),
            .in2(N__12897),
            .in3(N__11743),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_4 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_3 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_4 ),
            .clk(N__12120),
            .ce(),
            .sr(N__12716));
    defparam \DUT.uart_inst0.tx_clk_divider_5_LC_18_19_5 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_5_LC_18_19_5 .SEQ_MODE=4'b1001;
    defparam \DUT.uart_inst0.tx_clk_divider_5_LC_18_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_5_LC_18_19_5  (
            .in0(_gnd_net_),
            .in1(N__11740),
            .in2(N__12894),
            .in3(N__11728),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_5 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_4 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_5 ),
            .clk(N__12120),
            .ce(),
            .sr(N__12716));
    defparam \DUT.uart_inst0.tx_clk_divider_6_LC_18_19_6 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_6_LC_18_19_6 .SEQ_MODE=4'b1001;
    defparam \DUT.uart_inst0.tx_clk_divider_6_LC_18_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_6_LC_18_19_6  (
            .in0(_gnd_net_),
            .in1(N__11725),
            .in2(N__12898),
            .in3(N__11713),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_6 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_5 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_6 ),
            .clk(N__12120),
            .ce(),
            .sr(N__12716));
    defparam \DUT.uart_inst0.tx_clk_divider_7_LC_18_19_7 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_7_LC_18_19_7 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_7_LC_18_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_7_LC_18_19_7  (
            .in0(_gnd_net_),
            .in1(N__11710),
            .in2(N__12895),
            .in3(N__11698),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_7 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_6 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_7 ),
            .clk(N__12120),
            .ce(),
            .sr(N__12716));
    defparam \DUT.uart_inst0.tx_clk_divider_8_LC_18_20_0 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_8_LC_18_20_0 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_8_LC_18_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_8_LC_18_20_0  (
            .in0(_gnd_net_),
            .in1(N__11695),
            .in2(N__12979),
            .in3(N__11683),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_8 ),
            .ltout(),
            .carryin(bfn_18_20_0_),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_8 ),
            .clk(N__12114),
            .ce(),
            .sr(N__12729));
    defparam \DUT.uart_inst0.tx_clk_divider_9_LC_18_20_1 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_9_LC_18_20_1 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_9_LC_18_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_9_LC_18_20_1  (
            .in0(_gnd_net_),
            .in1(N__11680),
            .in2(N__12981),
            .in3(N__11668),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_9 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_8 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_9 ),
            .clk(N__12114),
            .ce(),
            .sr(N__12729));
    defparam \DUT.uart_inst0.tx_clk_divider_10_LC_18_20_2 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_10_LC_18_20_2 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_10_LC_18_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_10_LC_18_20_2  (
            .in0(_gnd_net_),
            .in1(N__11665),
            .in2(N__12977),
            .in3(N__11653),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_10 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_9 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_10 ),
            .clk(N__12114),
            .ce(),
            .sr(N__12729));
    defparam \DUT.uart_inst0.tx_clk_divider_11_LC_18_20_3 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_11_LC_18_20_3 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_11_LC_18_20_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_11_LC_18_20_3  (
            .in0(_gnd_net_),
            .in1(N__11649),
            .in2(N__12980),
            .in3(N__11635),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_11 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_10 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_11 ),
            .clk(N__12114),
            .ce(),
            .sr(N__12729));
    defparam \DUT.uart_inst0.tx_clk_divider_12_LC_18_20_4 .C_ON=1'b1;
    defparam \DUT.uart_inst0.tx_clk_divider_12_LC_18_20_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_12_LC_18_20_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_12_LC_18_20_4  (
            .in0(_gnd_net_),
            .in1(N__12763),
            .in2(N__12978),
            .in3(N__12751),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_12 ),
            .ltout(),
            .carryin(\DUT.uart_inst0.tx_clk_divider_cry_11 ),
            .carryout(\DUT.uart_inst0.tx_clk_divider_cry_12 ),
            .clk(N__12114),
            .ce(),
            .sr(N__12729));
    defparam \DUT.uart_inst0.tx_clk_divider_13_LC_18_20_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_clk_divider_13_LC_18_20_5 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_clk_divider_13_LC_18_20_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \DUT.uart_inst0.tx_clk_divider_13_LC_18_20_5  (
            .in0(_gnd_net_),
            .in1(N__12744),
            .in2(_gnd_net_),
            .in3(N__12748),
            .lcout(\DUT.uart_inst0.tx_clk_dividerZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12114),
            .ce(),
            .sr(N__12729));
    defparam \DUT.uart_inst0.tx_state_0_LC_18_21_4 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_state_0_LC_18_21_4 .SEQ_MODE=4'b1000;
    defparam \DUT.uart_inst0.tx_state_0_LC_18_21_4 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \DUT.uart_inst0.tx_state_0_LC_18_21_4  (
            .in0(N__12703),
            .in1(N__12697),
            .in2(_gnd_net_),
            .in3(N__12682),
            .lcout(\DUT.tx_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12108),
            .ce(),
            .sr(N__12494));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_18_21_5 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_18_21_5 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_18_21_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNO_0_3_LC_18_21_5  (
            .in0(N__12234),
            .in1(N__12445),
            .in2(_gnd_net_),
            .in3(N__12406),
            .lcout(\DUT.uart_inst0.tx_bits_remaining_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_0_2_LC_18_21_6 .C_ON=1'b0;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_0_2_LC_18_21_6 .SEQ_MODE=4'b0000;
    defparam \DUT.uart_inst0.tx_bits_remaining_RNO_0_2_LC_18_21_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \DUT.uart_inst0.tx_bits_remaining_RNO_0_2_LC_18_21_6  (
            .in0(N__11939),
            .in1(N__12321),
            .in2(_gnd_net_),
            .in3(N__12233),
            .lcout(\DUT.uart_inst0.tx_bits_remaining_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ftdi_output_inst.rRxF_n_0_LC_18_23_4 .C_ON=1'b0;
    defparam \fifo_inst.ftdi_output_inst.rRxF_n_0_LC_18_23_4 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ftdi_output_inst.rRxF_n_0_LC_18_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.ftdi_output_inst.rRxF_n_0_LC_18_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12175),
            .lcout(\fifo_inst.ftdi_output_inst.rRxF_nZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__12096),
            .ce(N__11868),
            .sr(_gnd_net_));
endmodule // top
