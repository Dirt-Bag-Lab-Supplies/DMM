// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Apr 5 2020 01:05:16

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top" view "INTERFACE"

module top (
    ioFifoData,
    P1A9,
    P1A1,
    P1A8,
    oRx_n,
    P1A7,
    P1A3,
    iTxE_n,
    iRxF_n,
    iClk,
    P1A2,
    BTN_N,
    BTN1,
    oTx_n,
    P1A4);

    inout [7:0] ioFifoData;
    output P1A9;
    input P1A1;
    output P1A8;
    output oRx_n;
    output P1A7;
    output P1A3;
    input iTxE_n;
    input iRxF_n;
    input iClk;
    output P1A2;
    input BTN_N;
    input BTN1;
    output oTx_n;
    output P1A4;

    wire N__17429;
    wire N__17415;
    wire N__17414;
    wire N__17413;
    wire N__17406;
    wire N__17405;
    wire N__17404;
    wire N__17397;
    wire N__17396;
    wire N__17395;
    wire N__17388;
    wire N__17387;
    wire N__17386;
    wire N__17379;
    wire N__17378;
    wire N__17377;
    wire N__17370;
    wire N__17369;
    wire N__17368;
    wire N__17361;
    wire N__17360;
    wire N__17359;
    wire N__17352;
    wire N__17351;
    wire N__17350;
    wire N__17343;
    wire N__17342;
    wire N__17341;
    wire N__17334;
    wire N__17333;
    wire N__17332;
    wire N__17325;
    wire N__17324;
    wire N__17323;
    wire N__17316;
    wire N__17315;
    wire N__17314;
    wire N__17307;
    wire N__17306;
    wire N__17305;
    wire N__17298;
    wire N__17297;
    wire N__17296;
    wire N__17289;
    wire N__17288;
    wire N__17287;
    wire N__17280;
    wire N__17279;
    wire N__17278;
    wire N__17271;
    wire N__17270;
    wire N__17269;
    wire N__17262;
    wire N__17261;
    wire N__17260;
    wire N__17253;
    wire N__17252;
    wire N__17251;
    wire N__17244;
    wire N__17243;
    wire N__17242;
    wire N__17225;
    wire N__17222;
    wire N__17219;
    wire N__17216;
    wire N__17213;
    wire N__17210;
    wire N__17209;
    wire N__17206;
    wire N__17203;
    wire N__17200;
    wire N__17195;
    wire N__17192;
    wire N__17189;
    wire N__17186;
    wire N__17183;
    wire N__17182;
    wire N__17179;
    wire N__17176;
    wire N__17173;
    wire N__17168;
    wire N__17165;
    wire N__17162;
    wire N__17159;
    wire N__17156;
    wire N__17155;
    wire N__17152;
    wire N__17149;
    wire N__17144;
    wire N__17141;
    wire N__17138;
    wire N__17135;
    wire N__17132;
    wire N__17129;
    wire N__17128;
    wire N__17125;
    wire N__17122;
    wire N__17117;
    wire N__17114;
    wire N__17111;
    wire N__17108;
    wire N__17105;
    wire N__17102;
    wire N__17099;
    wire N__17096;
    wire N__17095;
    wire N__17092;
    wire N__17089;
    wire N__17084;
    wire N__17081;
    wire N__17078;
    wire N__17075;
    wire N__17072;
    wire N__17069;
    wire N__17066;
    wire N__17063;
    wire N__17062;
    wire N__17061;
    wire N__17060;
    wire N__17059;
    wire N__17058;
    wire N__17057;
    wire N__17044;
    wire N__17041;
    wire N__17040;
    wire N__17035;
    wire N__17032;
    wire N__17029;
    wire N__17028;
    wire N__17027;
    wire N__17022;
    wire N__17019;
    wire N__17016;
    wire N__17011;
    wire N__17006;
    wire N__17005;
    wire N__17002;
    wire N__16999;
    wire N__16996;
    wire N__16991;
    wire N__16990;
    wire N__16989;
    wire N__16988;
    wire N__16987;
    wire N__16986;
    wire N__16985;
    wire N__16984;
    wire N__16983;
    wire N__16982;
    wire N__16981;
    wire N__16980;
    wire N__16979;
    wire N__16978;
    wire N__16977;
    wire N__16976;
    wire N__16975;
    wire N__16974;
    wire N__16973;
    wire N__16972;
    wire N__16971;
    wire N__16970;
    wire N__16969;
    wire N__16968;
    wire N__16967;
    wire N__16966;
    wire N__16965;
    wire N__16964;
    wire N__16963;
    wire N__16962;
    wire N__16961;
    wire N__16960;
    wire N__16959;
    wire N__16958;
    wire N__16957;
    wire N__16956;
    wire N__16955;
    wire N__16954;
    wire N__16953;
    wire N__16952;
    wire N__16951;
    wire N__16950;
    wire N__16949;
    wire N__16948;
    wire N__16947;
    wire N__16946;
    wire N__16945;
    wire N__16944;
    wire N__16943;
    wire N__16942;
    wire N__16941;
    wire N__16940;
    wire N__16939;
    wire N__16938;
    wire N__16937;
    wire N__16936;
    wire N__16935;
    wire N__16934;
    wire N__16933;
    wire N__16932;
    wire N__16931;
    wire N__16930;
    wire N__16929;
    wire N__16928;
    wire N__16927;
    wire N__16926;
    wire N__16925;
    wire N__16924;
    wire N__16923;
    wire N__16922;
    wire N__16921;
    wire N__16920;
    wire N__16919;
    wire N__16918;
    wire N__16917;
    wire N__16916;
    wire N__16915;
    wire N__16914;
    wire N__16913;
    wire N__16912;
    wire N__16911;
    wire N__16910;
    wire N__16909;
    wire N__16908;
    wire N__16907;
    wire N__16906;
    wire N__16905;
    wire N__16904;
    wire N__16903;
    wire N__16902;
    wire N__16901;
    wire N__16900;
    wire N__16899;
    wire N__16898;
    wire N__16897;
    wire N__16706;
    wire N__16703;
    wire N__16702;
    wire N__16701;
    wire N__16700;
    wire N__16699;
    wire N__16698;
    wire N__16697;
    wire N__16696;
    wire N__16695;
    wire N__16694;
    wire N__16693;
    wire N__16690;
    wire N__16689;
    wire N__16688;
    wire N__16687;
    wire N__16686;
    wire N__16685;
    wire N__16684;
    wire N__16683;
    wire N__16682;
    wire N__16681;
    wire N__16680;
    wire N__16679;
    wire N__16678;
    wire N__16677;
    wire N__16676;
    wire N__16675;
    wire N__16674;
    wire N__16671;
    wire N__16670;
    wire N__16667;
    wire N__16666;
    wire N__16665;
    wire N__16664;
    wire N__16663;
    wire N__16662;
    wire N__16661;
    wire N__16660;
    wire N__16659;
    wire N__16658;
    wire N__16657;
    wire N__16654;
    wire N__16653;
    wire N__16650;
    wire N__16649;
    wire N__16646;
    wire N__16645;
    wire N__16644;
    wire N__16641;
    wire N__16640;
    wire N__16639;
    wire N__16638;
    wire N__16637;
    wire N__16636;
    wire N__16635;
    wire N__16634;
    wire N__16633;
    wire N__16632;
    wire N__16631;
    wire N__16630;
    wire N__16629;
    wire N__16628;
    wire N__16627;
    wire N__16626;
    wire N__16625;
    wire N__16624;
    wire N__16623;
    wire N__16622;
    wire N__16621;
    wire N__16620;
    wire N__16619;
    wire N__16618;
    wire N__16615;
    wire N__16610;
    wire N__16607;
    wire N__16594;
    wire N__16589;
    wire N__16580;
    wire N__16577;
    wire N__16572;
    wire N__16569;
    wire N__16566;
    wire N__16563;
    wire N__16560;
    wire N__16555;
    wire N__16548;
    wire N__16541;
    wire N__16538;
    wire N__16531;
    wire N__16526;
    wire N__16523;
    wire N__16518;
    wire N__16511;
    wire N__16504;
    wire N__16497;
    wire N__16490;
    wire N__16483;
    wire N__16480;
    wire N__16473;
    wire N__16466;
    wire N__16459;
    wire N__16456;
    wire N__16455;
    wire N__16454;
    wire N__16453;
    wire N__16450;
    wire N__16449;
    wire N__16448;
    wire N__16445;
    wire N__16442;
    wire N__16439;
    wire N__16438;
    wire N__16437;
    wire N__16436;
    wire N__16433;
    wire N__16430;
    wire N__16429;
    wire N__16426;
    wire N__16425;
    wire N__16422;
    wire N__16421;
    wire N__16420;
    wire N__16419;
    wire N__16418;
    wire N__16417;
    wire N__16416;
    wire N__16415;
    wire N__16414;
    wire N__16413;
    wire N__16410;
    wire N__16407;
    wire N__16404;
    wire N__16401;
    wire N__16398;
    wire N__16395;
    wire N__16392;
    wire N__16389;
    wire N__16386;
    wire N__16385;
    wire N__16384;
    wire N__16381;
    wire N__16378;
    wire N__16375;
    wire N__16372;
    wire N__16369;
    wire N__16368;
    wire N__16367;
    wire N__16366;
    wire N__16363;
    wire N__16360;
    wire N__16359;
    wire N__16358;
    wire N__16357;
    wire N__16356;
    wire N__16355;
    wire N__16352;
    wire N__16351;
    wire N__16350;
    wire N__16347;
    wire N__16344;
    wire N__16341;
    wire N__16340;
    wire N__16217;
    wire N__16214;
    wire N__16211;
    wire N__16210;
    wire N__16207;
    wire N__16204;
    wire N__16201;
    wire N__16196;
    wire N__16193;
    wire N__16192;
    wire N__16189;
    wire N__16186;
    wire N__16183;
    wire N__16178;
    wire N__16175;
    wire N__16172;
    wire N__16169;
    wire N__16166;
    wire N__16163;
    wire N__16162;
    wire N__16159;
    wire N__16156;
    wire N__16153;
    wire N__16148;
    wire N__16147;
    wire N__16144;
    wire N__16141;
    wire N__16138;
    wire N__16137;
    wire N__16134;
    wire N__16131;
    wire N__16128;
    wire N__16125;
    wire N__16118;
    wire N__16115;
    wire N__16114;
    wire N__16111;
    wire N__16108;
    wire N__16105;
    wire N__16100;
    wire N__16097;
    wire N__16096;
    wire N__16093;
    wire N__16090;
    wire N__16087;
    wire N__16082;
    wire N__16081;
    wire N__16078;
    wire N__16075;
    wire N__16072;
    wire N__16067;
    wire N__16066;
    wire N__16063;
    wire N__16060;
    wire N__16057;
    wire N__16054;
    wire N__16049;
    wire N__16048;
    wire N__16045;
    wire N__16044;
    wire N__16041;
    wire N__16038;
    wire N__16037;
    wire N__16036;
    wire N__16035;
    wire N__16034;
    wire N__16033;
    wire N__16032;
    wire N__16029;
    wire N__16026;
    wire N__16023;
    wire N__16022;
    wire N__16019;
    wire N__16014;
    wire N__16009;
    wire N__16004;
    wire N__16001;
    wire N__15998;
    wire N__15995;
    wire N__15990;
    wire N__15985;
    wire N__15974;
    wire N__15973;
    wire N__15970;
    wire N__15969;
    wire N__15966;
    wire N__15965;
    wire N__15964;
    wire N__15961;
    wire N__15958;
    wire N__15953;
    wire N__15950;
    wire N__15943;
    wire N__15938;
    wire N__15937;
    wire N__15934;
    wire N__15933;
    wire N__15930;
    wire N__15927;
    wire N__15924;
    wire N__15923;
    wire N__15922;
    wire N__15921;
    wire N__15920;
    wire N__15913;
    wire N__15910;
    wire N__15903;
    wire N__15896;
    wire N__15895;
    wire N__15892;
    wire N__15891;
    wire N__15888;
    wire N__15885;
    wire N__15882;
    wire N__15875;
    wire N__15874;
    wire N__15871;
    wire N__15868;
    wire N__15865;
    wire N__15864;
    wire N__15861;
    wire N__15858;
    wire N__15855;
    wire N__15848;
    wire N__15845;
    wire N__15842;
    wire N__15839;
    wire N__15836;
    wire N__15835;
    wire N__15832;
    wire N__15829;
    wire N__15824;
    wire N__15823;
    wire N__15822;
    wire N__15821;
    wire N__15818;
    wire N__15815;
    wire N__15812;
    wire N__15809;
    wire N__15800;
    wire N__15799;
    wire N__15798;
    wire N__15795;
    wire N__15794;
    wire N__15791;
    wire N__15790;
    wire N__15789;
    wire N__15786;
    wire N__15783;
    wire N__15780;
    wire N__15777;
    wire N__15774;
    wire N__15771;
    wire N__15768;
    wire N__15755;
    wire N__15752;
    wire N__15751;
    wire N__15748;
    wire N__15745;
    wire N__15740;
    wire N__15737;
    wire N__15734;
    wire N__15731;
    wire N__15730;
    wire N__15727;
    wire N__15724;
    wire N__15719;
    wire N__15716;
    wire N__15713;
    wire N__15710;
    wire N__15709;
    wire N__15706;
    wire N__15703;
    wire N__15698;
    wire N__15695;
    wire N__15692;
    wire N__15689;
    wire N__15688;
    wire N__15685;
    wire N__15682;
    wire N__15677;
    wire N__15674;
    wire N__15671;
    wire N__15668;
    wire N__15665;
    wire N__15662;
    wire N__15659;
    wire N__15656;
    wire N__15655;
    wire N__15654;
    wire N__15651;
    wire N__15646;
    wire N__15641;
    wire N__15638;
    wire N__15637;
    wire N__15634;
    wire N__15631;
    wire N__15626;
    wire N__15623;
    wire N__15622;
    wire N__15619;
    wire N__15616;
    wire N__15613;
    wire N__15610;
    wire N__15605;
    wire N__15602;
    wire N__15599;
    wire N__15596;
    wire N__15595;
    wire N__15592;
    wire N__15589;
    wire N__15586;
    wire N__15581;
    wire N__15578;
    wire N__15575;
    wire N__15572;
    wire N__15569;
    wire N__15566;
    wire N__15563;
    wire N__15560;
    wire N__15557;
    wire N__15554;
    wire N__15551;
    wire N__15548;
    wire N__15545;
    wire N__15542;
    wire N__15539;
    wire N__15536;
    wire N__15533;
    wire N__15530;
    wire N__15527;
    wire N__15524;
    wire N__15521;
    wire N__15518;
    wire N__15515;
    wire N__15512;
    wire N__15511;
    wire N__15508;
    wire N__15505;
    wire N__15500;
    wire N__15497;
    wire N__15494;
    wire N__15491;
    wire N__15490;
    wire N__15487;
    wire N__15484;
    wire N__15479;
    wire N__15476;
    wire N__15473;
    wire N__15470;
    wire N__15467;
    wire N__15466;
    wire N__15463;
    wire N__15460;
    wire N__15455;
    wire N__15452;
    wire N__15449;
    wire N__15446;
    wire N__15445;
    wire N__15442;
    wire N__15439;
    wire N__15434;
    wire N__15431;
    wire N__15428;
    wire N__15425;
    wire N__15422;
    wire N__15419;
    wire N__15416;
    wire N__15413;
    wire N__15412;
    wire N__15411;
    wire N__15408;
    wire N__15403;
    wire N__15402;
    wire N__15401;
    wire N__15400;
    wire N__15399;
    wire N__15398;
    wire N__15397;
    wire N__15394;
    wire N__15391;
    wire N__15378;
    wire N__15377;
    wire N__15376;
    wire N__15369;
    wire N__15368;
    wire N__15367;
    wire N__15366;
    wire N__15365;
    wire N__15364;
    wire N__15363;
    wire N__15362;
    wire N__15361;
    wire N__15358;
    wire N__15355;
    wire N__15352;
    wire N__15349;
    wire N__15338;
    wire N__15331;
    wire N__15320;
    wire N__15319;
    wire N__15316;
    wire N__15313;
    wire N__15308;
    wire N__15305;
    wire N__15304;
    wire N__15301;
    wire N__15298;
    wire N__15293;
    wire N__15290;
    wire N__15287;
    wire N__15286;
    wire N__15283;
    wire N__15280;
    wire N__15277;
    wire N__15276;
    wire N__15271;
    wire N__15268;
    wire N__15263;
    wire N__15260;
    wire N__15257;
    wire N__15254;
    wire N__15253;
    wire N__15252;
    wire N__15249;
    wire N__15246;
    wire N__15243;
    wire N__15236;
    wire N__15233;
    wire N__15230;
    wire N__15229;
    wire N__15226;
    wire N__15225;
    wire N__15222;
    wire N__15219;
    wire N__15216;
    wire N__15209;
    wire N__15206;
    wire N__15203;
    wire N__15202;
    wire N__15199;
    wire N__15198;
    wire N__15195;
    wire N__15192;
    wire N__15189;
    wire N__15182;
    wire N__15179;
    wire N__15176;
    wire N__15173;
    wire N__15172;
    wire N__15169;
    wire N__15168;
    wire N__15165;
    wire N__15162;
    wire N__15159;
    wire N__15152;
    wire N__15149;
    wire N__15148;
    wire N__15145;
    wire N__15142;
    wire N__15137;
    wire N__15134;
    wire N__15131;
    wire N__15128;
    wire N__15127;
    wire N__15126;
    wire N__15123;
    wire N__15120;
    wire N__15117;
    wire N__15110;
    wire N__15107;
    wire N__15104;
    wire N__15101;
    wire N__15100;
    wire N__15099;
    wire N__15096;
    wire N__15093;
    wire N__15090;
    wire N__15083;
    wire N__15080;
    wire N__15079;
    wire N__15076;
    wire N__15073;
    wire N__15072;
    wire N__15069;
    wire N__15066;
    wire N__15063;
    wire N__15060;
    wire N__15053;
    wire N__15050;
    wire N__15047;
    wire N__15044;
    wire N__15043;
    wire N__15042;
    wire N__15039;
    wire N__15036;
    wire N__15033;
    wire N__15026;
    wire N__15025;
    wire N__15022;
    wire N__15017;
    wire N__15014;
    wire N__15011;
    wire N__15008;
    wire N__15007;
    wire N__15004;
    wire N__15001;
    wire N__14998;
    wire N__14993;
    wire N__14990;
    wire N__14987;
    wire N__14984;
    wire N__14983;
    wire N__14980;
    wire N__14977;
    wire N__14974;
    wire N__14969;
    wire N__14966;
    wire N__14963;
    wire N__14962;
    wire N__14961;
    wire N__14960;
    wire N__14957;
    wire N__14954;
    wire N__14951;
    wire N__14950;
    wire N__14949;
    wire N__14948;
    wire N__14947;
    wire N__14946;
    wire N__14945;
    wire N__14944;
    wire N__14943;
    wire N__14940;
    wire N__14937;
    wire N__14934;
    wire N__14931;
    wire N__14928;
    wire N__14925;
    wire N__14918;
    wire N__14911;
    wire N__14894;
    wire N__14893;
    wire N__14890;
    wire N__14887;
    wire N__14884;
    wire N__14879;
    wire N__14876;
    wire N__14873;
    wire N__14870;
    wire N__14867;
    wire N__14864;
    wire N__14861;
    wire N__14858;
    wire N__14855;
    wire N__14852;
    wire N__14849;
    wire N__14846;
    wire N__14843;
    wire N__14842;
    wire N__14841;
    wire N__14840;
    wire N__14837;
    wire N__14836;
    wire N__14831;
    wire N__14828;
    wire N__14825;
    wire N__14822;
    wire N__14815;
    wire N__14812;
    wire N__14807;
    wire N__14804;
    wire N__14801;
    wire N__14798;
    wire N__14797;
    wire N__14796;
    wire N__14793;
    wire N__14790;
    wire N__14787;
    wire N__14780;
    wire N__14777;
    wire N__14774;
    wire N__14771;
    wire N__14770;
    wire N__14767;
    wire N__14764;
    wire N__14761;
    wire N__14756;
    wire N__14753;
    wire N__14750;
    wire N__14749;
    wire N__14746;
    wire N__14743;
    wire N__14740;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14728;
    wire N__14725;
    wire N__14722;
    wire N__14717;
    wire N__14714;
    wire N__14711;
    wire N__14710;
    wire N__14707;
    wire N__14704;
    wire N__14699;
    wire N__14696;
    wire N__14693;
    wire N__14690;
    wire N__14689;
    wire N__14686;
    wire N__14683;
    wire N__14678;
    wire N__14675;
    wire N__14672;
    wire N__14671;
    wire N__14668;
    wire N__14665;
    wire N__14660;
    wire N__14657;
    wire N__14654;
    wire N__14653;
    wire N__14650;
    wire N__14647;
    wire N__14642;
    wire N__14639;
    wire N__14638;
    wire N__14637;
    wire N__14636;
    wire N__14635;
    wire N__14632;
    wire N__14629;
    wire N__14626;
    wire N__14623;
    wire N__14620;
    wire N__14617;
    wire N__14614;
    wire N__14607;
    wire N__14600;
    wire N__14599;
    wire N__14594;
    wire N__14593;
    wire N__14592;
    wire N__14591;
    wire N__14590;
    wire N__14587;
    wire N__14584;
    wire N__14581;
    wire N__14578;
    wire N__14575;
    wire N__14572;
    wire N__14569;
    wire N__14566;
    wire N__14555;
    wire N__14552;
    wire N__14551;
    wire N__14550;
    wire N__14549;
    wire N__14548;
    wire N__14547;
    wire N__14544;
    wire N__14543;
    wire N__14540;
    wire N__14537;
    wire N__14532;
    wire N__14529;
    wire N__14526;
    wire N__14523;
    wire N__14520;
    wire N__14517;
    wire N__14504;
    wire N__14501;
    wire N__14500;
    wire N__14497;
    wire N__14494;
    wire N__14489;
    wire N__14486;
    wire N__14483;
    wire N__14480;
    wire N__14477;
    wire N__14474;
    wire N__14471;
    wire N__14470;
    wire N__14467;
    wire N__14464;
    wire N__14459;
    wire N__14456;
    wire N__14453;
    wire N__14450;
    wire N__14449;
    wire N__14448;
    wire N__14445;
    wire N__14442;
    wire N__14439;
    wire N__14432;
    wire N__14431;
    wire N__14428;
    wire N__14425;
    wire N__14420;
    wire N__14419;
    wire N__14418;
    wire N__14415;
    wire N__14412;
    wire N__14409;
    wire N__14406;
    wire N__14399;
    wire N__14398;
    wire N__14397;
    wire N__14394;
    wire N__14391;
    wire N__14388;
    wire N__14381;
    wire N__14380;
    wire N__14377;
    wire N__14374;
    wire N__14371;
    wire N__14366;
    wire N__14363;
    wire N__14360;
    wire N__14357;
    wire N__14356;
    wire N__14353;
    wire N__14350;
    wire N__14347;
    wire N__14342;
    wire N__14339;
    wire N__14336;
    wire N__14333;
    wire N__14332;
    wire N__14331;
    wire N__14328;
    wire N__14325;
    wire N__14322;
    wire N__14315;
    wire N__14312;
    wire N__14309;
    wire N__14308;
    wire N__14307;
    wire N__14304;
    wire N__14301;
    wire N__14298;
    wire N__14295;
    wire N__14288;
    wire N__14287;
    wire N__14284;
    wire N__14281;
    wire N__14278;
    wire N__14275;
    wire N__14274;
    wire N__14271;
    wire N__14268;
    wire N__14265;
    wire N__14262;
    wire N__14255;
    wire N__14252;
    wire N__14249;
    wire N__14248;
    wire N__14245;
    wire N__14244;
    wire N__14241;
    wire N__14238;
    wire N__14235;
    wire N__14228;
    wire N__14225;
    wire N__14222;
    wire N__14219;
    wire N__14218;
    wire N__14217;
    wire N__14214;
    wire N__14211;
    wire N__14208;
    wire N__14201;
    wire N__14198;
    wire N__14195;
    wire N__14192;
    wire N__14189;
    wire N__14186;
    wire N__14183;
    wire N__14182;
    wire N__14181;
    wire N__14178;
    wire N__14175;
    wire N__14172;
    wire N__14165;
    wire N__14162;
    wire N__14159;
    wire N__14156;
    wire N__14155;
    wire N__14154;
    wire N__14151;
    wire N__14148;
    wire N__14145;
    wire N__14138;
    wire N__14135;
    wire N__14132;
    wire N__14131;
    wire N__14130;
    wire N__14127;
    wire N__14124;
    wire N__14121;
    wire N__14118;
    wire N__14115;
    wire N__14108;
    wire N__14105;
    wire N__14102;
    wire N__14101;
    wire N__14100;
    wire N__14097;
    wire N__14094;
    wire N__14091;
    wire N__14088;
    wire N__14085;
    wire N__14082;
    wire N__14081;
    wire N__14078;
    wire N__14075;
    wire N__14072;
    wire N__14069;
    wire N__14068;
    wire N__14063;
    wire N__14058;
    wire N__14055;
    wire N__14052;
    wire N__14049;
    wire N__14046;
    wire N__14039;
    wire N__14036;
    wire N__14035;
    wire N__14032;
    wire N__14029;
    wire N__14024;
    wire N__14023;
    wire N__14022;
    wire N__14021;
    wire N__14020;
    wire N__14017;
    wire N__14016;
    wire N__14015;
    wire N__14014;
    wire N__14013;
    wire N__14012;
    wire N__14011;
    wire N__14006;
    wire N__14005;
    wire N__14004;
    wire N__14003;
    wire N__14000;
    wire N__13999;
    wire N__13998;
    wire N__13995;
    wire N__13992;
    wire N__13987;
    wire N__13986;
    wire N__13983;
    wire N__13980;
    wire N__13977;
    wire N__13974;
    wire N__13971;
    wire N__13968;
    wire N__13963;
    wire N__13956;
    wire N__13953;
    wire N__13950;
    wire N__13947;
    wire N__13946;
    wire N__13943;
    wire N__13940;
    wire N__13937;
    wire N__13932;
    wire N__13929;
    wire N__13922;
    wire N__13921;
    wire N__13918;
    wire N__13913;
    wire N__13910;
    wire N__13907;
    wire N__13904;
    wire N__13895;
    wire N__13894;
    wire N__13891;
    wire N__13888;
    wire N__13885;
    wire N__13880;
    wire N__13875;
    wire N__13872;
    wire N__13869;
    wire N__13866;
    wire N__13857;
    wire N__13854;
    wire N__13851;
    wire N__13848;
    wire N__13845;
    wire N__13842;
    wire N__13839;
    wire N__13836;
    wire N__13829;
    wire N__13826;
    wire N__13825;
    wire N__13824;
    wire N__13823;
    wire N__13822;
    wire N__13819;
    wire N__13818;
    wire N__13817;
    wire N__13814;
    wire N__13807;
    wire N__13804;
    wire N__13799;
    wire N__13790;
    wire N__13787;
    wire N__13784;
    wire N__13781;
    wire N__13780;
    wire N__13779;
    wire N__13778;
    wire N__13775;
    wire N__13772;
    wire N__13771;
    wire N__13768;
    wire N__13765;
    wire N__13762;
    wire N__13759;
    wire N__13756;
    wire N__13749;
    wire N__13746;
    wire N__13739;
    wire N__13738;
    wire N__13735;
    wire N__13732;
    wire N__13729;
    wire N__13724;
    wire N__13721;
    wire N__13720;
    wire N__13719;
    wire N__13716;
    wire N__13713;
    wire N__13710;
    wire N__13707;
    wire N__13700;
    wire N__13697;
    wire N__13696;
    wire N__13693;
    wire N__13690;
    wire N__13685;
    wire N__13684;
    wire N__13681;
    wire N__13680;
    wire N__13679;
    wire N__13676;
    wire N__13673;
    wire N__13670;
    wire N__13667;
    wire N__13664;
    wire N__13661;
    wire N__13658;
    wire N__13655;
    wire N__13652;
    wire N__13643;
    wire N__13640;
    wire N__13637;
    wire N__13634;
    wire N__13631;
    wire N__13630;
    wire N__13629;
    wire N__13628;
    wire N__13625;
    wire N__13622;
    wire N__13619;
    wire N__13616;
    wire N__13611;
    wire N__13604;
    wire N__13603;
    wire N__13602;
    wire N__13601;
    wire N__13600;
    wire N__13599;
    wire N__13598;
    wire N__13597;
    wire N__13596;
    wire N__13595;
    wire N__13594;
    wire N__13593;
    wire N__13592;
    wire N__13591;
    wire N__13562;
    wire N__13559;
    wire N__13556;
    wire N__13555;
    wire N__13554;
    wire N__13551;
    wire N__13550;
    wire N__13549;
    wire N__13548;
    wire N__13547;
    wire N__13546;
    wire N__13545;
    wire N__13544;
    wire N__13543;
    wire N__13542;
    wire N__13541;
    wire N__13538;
    wire N__13529;
    wire N__13526;
    wire N__13511;
    wire N__13510;
    wire N__13505;
    wire N__13500;
    wire N__13497;
    wire N__13490;
    wire N__13487;
    wire N__13484;
    wire N__13483;
    wire N__13480;
    wire N__13477;
    wire N__13472;
    wire N__13469;
    wire N__13466;
    wire N__13463;
    wire N__13460;
    wire N__13457;
    wire N__13456;
    wire N__13453;
    wire N__13450;
    wire N__13447;
    wire N__13442;
    wire N__13441;
    wire N__13438;
    wire N__13435;
    wire N__13430;
    wire N__13427;
    wire N__13426;
    wire N__13423;
    wire N__13420;
    wire N__13415;
    wire N__13414;
    wire N__13411;
    wire N__13408;
    wire N__13403;
    wire N__13400;
    wire N__13397;
    wire N__13394;
    wire N__13393;
    wire N__13388;
    wire N__13385;
    wire N__13382;
    wire N__13379;
    wire N__13376;
    wire N__13373;
    wire N__13372;
    wire N__13371;
    wire N__13370;
    wire N__13367;
    wire N__13364;
    wire N__13359;
    wire N__13352;
    wire N__13351;
    wire N__13348;
    wire N__13345;
    wire N__13342;
    wire N__13337;
    wire N__13334;
    wire N__13333;
    wire N__13330;
    wire N__13327;
    wire N__13324;
    wire N__13319;
    wire N__13318;
    wire N__13317;
    wire N__13316;
    wire N__13315;
    wire N__13312;
    wire N__13309;
    wire N__13304;
    wire N__13299;
    wire N__13298;
    wire N__13291;
    wire N__13290;
    wire N__13287;
    wire N__13284;
    wire N__13281;
    wire N__13274;
    wire N__13271;
    wire N__13268;
    wire N__13265;
    wire N__13264;
    wire N__13263;
    wire N__13260;
    wire N__13259;
    wire N__13258;
    wire N__13255;
    wire N__13254;
    wire N__13251;
    wire N__13250;
    wire N__13247;
    wire N__13242;
    wire N__13239;
    wire N__13236;
    wire N__13231;
    wire N__13226;
    wire N__13217;
    wire N__13216;
    wire N__13213;
    wire N__13210;
    wire N__13205;
    wire N__13202;
    wire N__13199;
    wire N__13196;
    wire N__13193;
    wire N__13190;
    wire N__13187;
    wire N__13184;
    wire N__13181;
    wire N__13180;
    wire N__13177;
    wire N__13174;
    wire N__13169;
    wire N__13168;
    wire N__13165;
    wire N__13162;
    wire N__13157;
    wire N__13156;
    wire N__13155;
    wire N__13154;
    wire N__13151;
    wire N__13148;
    wire N__13147;
    wire N__13146;
    wire N__13143;
    wire N__13142;
    wire N__13141;
    wire N__13140;
    wire N__13137;
    wire N__13134;
    wire N__13131;
    wire N__13126;
    wire N__13123;
    wire N__13118;
    wire N__13115;
    wire N__13110;
    wire N__13103;
    wire N__13094;
    wire N__13093;
    wire N__13092;
    wire N__13091;
    wire N__13090;
    wire N__13089;
    wire N__13088;
    wire N__13085;
    wire N__13082;
    wire N__13075;
    wire N__13070;
    wire N__13061;
    wire N__13058;
    wire N__13055;
    wire N__13052;
    wire N__13049;
    wire N__13046;
    wire N__13043;
    wire N__13042;
    wire N__13041;
    wire N__13040;
    wire N__13037;
    wire N__13034;
    wire N__13031;
    wire N__13028;
    wire N__13019;
    wire N__13016;
    wire N__13013;
    wire N__13012;
    wire N__13007;
    wire N__13004;
    wire N__13003;
    wire N__13002;
    wire N__13001;
    wire N__13000;
    wire N__12997;
    wire N__12994;
    wire N__12991;
    wire N__12986;
    wire N__12981;
    wire N__12974;
    wire N__12971;
    wire N__12968;
    wire N__12967;
    wire N__12966;
    wire N__12963;
    wire N__12962;
    wire N__12959;
    wire N__12958;
    wire N__12957;
    wire N__12954;
    wire N__12949;
    wire N__12942;
    wire N__12935;
    wire N__12934;
    wire N__12931;
    wire N__12930;
    wire N__12929;
    wire N__12928;
    wire N__12927;
    wire N__12922;
    wire N__12917;
    wire N__12912;
    wire N__12905;
    wire N__12902;
    wire N__12899;
    wire N__12896;
    wire N__12893;
    wire N__12890;
    wire N__12887;
    wire N__12884;
    wire N__12881;
    wire N__12878;
    wire N__12875;
    wire N__12872;
    wire N__12869;
    wire N__12866;
    wire N__12863;
    wire N__12860;
    wire N__12857;
    wire N__12854;
    wire N__12851;
    wire N__12850;
    wire N__12847;
    wire N__12844;
    wire N__12841;
    wire N__12838;
    wire N__12835;
    wire N__12832;
    wire N__12827;
    wire N__12824;
    wire N__12821;
    wire N__12818;
    wire N__12815;
    wire N__12812;
    wire N__12809;
    wire N__12806;
    wire N__12803;
    wire N__12800;
    wire N__12797;
    wire N__12796;
    wire N__12793;
    wire N__12790;
    wire N__12787;
    wire N__12784;
    wire N__12779;
    wire N__12776;
    wire N__12775;
    wire N__12772;
    wire N__12769;
    wire N__12764;
    wire N__12763;
    wire N__12762;
    wire N__12759;
    wire N__12758;
    wire N__12757;
    wire N__12756;
    wire N__12755;
    wire N__12754;
    wire N__12751;
    wire N__12750;
    wire N__12749;
    wire N__12746;
    wire N__12743;
    wire N__12732;
    wire N__12729;
    wire N__12726;
    wire N__12725;
    wire N__12722;
    wire N__12719;
    wire N__12712;
    wire N__12709;
    wire N__12706;
    wire N__12695;
    wire N__12692;
    wire N__12691;
    wire N__12690;
    wire N__12689;
    wire N__12688;
    wire N__12687;
    wire N__12686;
    wire N__12683;
    wire N__12680;
    wire N__12675;
    wire N__12668;
    wire N__12665;
    wire N__12656;
    wire N__12653;
    wire N__12652;
    wire N__12651;
    wire N__12650;
    wire N__12647;
    wire N__12646;
    wire N__12645;
    wire N__12642;
    wire N__12641;
    wire N__12638;
    wire N__12637;
    wire N__12634;
    wire N__12631;
    wire N__12628;
    wire N__12625;
    wire N__12618;
    wire N__12613;
    wire N__12610;
    wire N__12599;
    wire N__12598;
    wire N__12595;
    wire N__12594;
    wire N__12593;
    wire N__12592;
    wire N__12589;
    wire N__12588;
    wire N__12587;
    wire N__12586;
    wire N__12583;
    wire N__12580;
    wire N__12577;
    wire N__12574;
    wire N__12567;
    wire N__12564;
    wire N__12561;
    wire N__12548;
    wire N__12545;
    wire N__12542;
    wire N__12539;
    wire N__12536;
    wire N__12533;
    wire N__12530;
    wire N__12527;
    wire N__12524;
    wire N__12521;
    wire N__12518;
    wire N__12515;
    wire N__12512;
    wire N__12509;
    wire N__12506;
    wire N__12503;
    wire N__12502;
    wire N__12501;
    wire N__12498;
    wire N__12495;
    wire N__12492;
    wire N__12487;
    wire N__12482;
    wire N__12479;
    wire N__12476;
    wire N__12473;
    wire N__12470;
    wire N__12467;
    wire N__12464;
    wire N__12461;
    wire N__12460;
    wire N__12459;
    wire N__12458;
    wire N__12457;
    wire N__12456;
    wire N__12455;
    wire N__12454;
    wire N__12453;
    wire N__12452;
    wire N__12451;
    wire N__12450;
    wire N__12449;
    wire N__12446;
    wire N__12443;
    wire N__12440;
    wire N__12439;
    wire N__12436;
    wire N__12433;
    wire N__12430;
    wire N__12427;
    wire N__12424;
    wire N__12421;
    wire N__12418;
    wire N__12415;
    wire N__12412;
    wire N__12409;
    wire N__12408;
    wire N__12407;
    wire N__12406;
    wire N__12405;
    wire N__12404;
    wire N__12403;
    wire N__12402;
    wire N__12399;
    wire N__12390;
    wire N__12385;
    wire N__12378;
    wire N__12369;
    wire N__12366;
    wire N__12363;
    wire N__12360;
    wire N__12357;
    wire N__12356;
    wire N__12353;
    wire N__12352;
    wire N__12349;
    wire N__12348;
    wire N__12345;
    wire N__12344;
    wire N__12343;
    wire N__12342;
    wire N__12341;
    wire N__12340;
    wire N__12339;
    wire N__12338;
    wire N__12327;
    wire N__12322;
    wire N__12317;
    wire N__12316;
    wire N__12315;
    wire N__12314;
    wire N__12313;
    wire N__12300;
    wire N__12297;
    wire N__12294;
    wire N__12291;
    wire N__12288;
    wire N__12285;
    wire N__12282;
    wire N__12279;
    wire N__12278;
    wire N__12271;
    wire N__12268;
    wire N__12267;
    wire N__12264;
    wire N__12261;
    wire N__12258;
    wire N__12257;
    wire N__12256;
    wire N__12253;
    wire N__12246;
    wire N__12237;
    wire N__12234;
    wire N__12229;
    wire N__12226;
    wire N__12223;
    wire N__12218;
    wire N__12215;
    wire N__12212;
    wire N__12205;
    wire N__12202;
    wire N__12197;
    wire N__12192;
    wire N__12189;
    wire N__12186;
    wire N__12183;
    wire N__12180;
    wire N__12177;
    wire N__12172;
    wire N__12169;
    wire N__12166;
    wire N__12163;
    wire N__12158;
    wire N__12149;
    wire N__12148;
    wire N__12145;
    wire N__12144;
    wire N__12141;
    wire N__12138;
    wire N__12133;
    wire N__12128;
    wire N__12125;
    wire N__12122;
    wire N__12119;
    wire N__12116;
    wire N__12115;
    wire N__12112;
    wire N__12109;
    wire N__12104;
    wire N__12101;
    wire N__12098;
    wire N__12095;
    wire N__12092;
    wire N__12089;
    wire N__12086;
    wire N__12083;
    wire N__12080;
    wire N__12077;
    wire N__12076;
    wire N__12075;
    wire N__12072;
    wire N__12069;
    wire N__12066;
    wire N__12063;
    wire N__12056;
    wire N__12053;
    wire N__12050;
    wire N__12047;
    wire N__12046;
    wire N__12045;
    wire N__12042;
    wire N__12039;
    wire N__12036;
    wire N__12029;
    wire N__12026;
    wire N__12023;
    wire N__12020;
    wire N__12019;
    wire N__12018;
    wire N__12015;
    wire N__12012;
    wire N__12009;
    wire N__12002;
    wire N__11999;
    wire N__11996;
    wire N__11993;
    wire N__11992;
    wire N__11989;
    wire N__11988;
    wire N__11985;
    wire N__11982;
    wire N__11979;
    wire N__11972;
    wire N__11969;
    wire N__11966;
    wire N__11963;
    wire N__11960;
    wire N__11959;
    wire N__11956;
    wire N__11955;
    wire N__11952;
    wire N__11949;
    wire N__11946;
    wire N__11939;
    wire N__11936;
    wire N__11933;
    wire N__11930;
    wire N__11927;
    wire N__11926;
    wire N__11925;
    wire N__11922;
    wire N__11917;
    wire N__11912;
    wire N__11909;
    wire N__11906;
    wire N__11903;
    wire N__11902;
    wire N__11901;
    wire N__11898;
    wire N__11893;
    wire N__11888;
    wire N__11885;
    wire N__11882;
    wire N__11879;
    wire N__11876;
    wire N__11875;
    wire N__11874;
    wire N__11873;
    wire N__11868;
    wire N__11865;
    wire N__11862;
    wire N__11861;
    wire N__11860;
    wire N__11859;
    wire N__11858;
    wire N__11857;
    wire N__11856;
    wire N__11855;
    wire N__11854;
    wire N__11853;
    wire N__11850;
    wire N__11845;
    wire N__11840;
    wire N__11831;
    wire N__11824;
    wire N__11813;
    wire N__11810;
    wire N__11807;
    wire N__11804;
    wire N__11801;
    wire N__11798;
    wire N__11795;
    wire N__11792;
    wire N__11789;
    wire N__11788;
    wire N__11787;
    wire N__11784;
    wire N__11781;
    wire N__11778;
    wire N__11771;
    wire N__11768;
    wire N__11765;
    wire N__11762;
    wire N__11759;
    wire N__11756;
    wire N__11753;
    wire N__11752;
    wire N__11751;
    wire N__11750;
    wire N__11749;
    wire N__11748;
    wire N__11745;
    wire N__11734;
    wire N__11729;
    wire N__11726;
    wire N__11725;
    wire N__11722;
    wire N__11719;
    wire N__11716;
    wire N__11711;
    wire N__11710;
    wire N__11707;
    wire N__11704;
    wire N__11701;
    wire N__11698;
    wire N__11693;
    wire N__11692;
    wire N__11691;
    wire N__11688;
    wire N__11685;
    wire N__11682;
    wire N__11675;
    wire N__11672;
    wire N__11669;
    wire N__11666;
    wire N__11665;
    wire N__11662;
    wire N__11661;
    wire N__11660;
    wire N__11659;
    wire N__11658;
    wire N__11655;
    wire N__11654;
    wire N__11653;
    wire N__11652;
    wire N__11651;
    wire N__11650;
    wire N__11649;
    wire N__11648;
    wire N__11645;
    wire N__11640;
    wire N__11637;
    wire N__11634;
    wire N__11631;
    wire N__11628;
    wire N__11625;
    wire N__11620;
    wire N__11613;
    wire N__11606;
    wire N__11591;
    wire N__11588;
    wire N__11587;
    wire N__11584;
    wire N__11583;
    wire N__11582;
    wire N__11581;
    wire N__11580;
    wire N__11579;
    wire N__11576;
    wire N__11575;
    wire N__11572;
    wire N__11569;
    wire N__11566;
    wire N__11565;
    wire N__11562;
    wire N__11561;
    wire N__11560;
    wire N__11557;
    wire N__11556;
    wire N__11553;
    wire N__11552;
    wire N__11549;
    wire N__11546;
    wire N__11543;
    wire N__11540;
    wire N__11535;
    wire N__11528;
    wire N__11521;
    wire N__11518;
    wire N__11501;
    wire N__11498;
    wire N__11495;
    wire N__11492;
    wire N__11489;
    wire N__11486;
    wire N__11483;
    wire N__11482;
    wire N__11479;
    wire N__11476;
    wire N__11473;
    wire N__11470;
    wire N__11465;
    wire N__11464;
    wire N__11459;
    wire N__11456;
    wire N__11455;
    wire N__11452;
    wire N__11449;
    wire N__11444;
    wire N__11441;
    wire N__11438;
    wire N__11435;
    wire N__11432;
    wire N__11431;
    wire N__11430;
    wire N__11429;
    wire N__11428;
    wire N__11425;
    wire N__11422;
    wire N__11419;
    wire N__11414;
    wire N__11405;
    wire N__11404;
    wire N__11403;
    wire N__11402;
    wire N__11399;
    wire N__11396;
    wire N__11391;
    wire N__11384;
    wire N__11381;
    wire N__11378;
    wire N__11375;
    wire N__11374;
    wire N__11371;
    wire N__11368;
    wire N__11363;
    wire N__11360;
    wire N__11357;
    wire N__11354;
    wire N__11353;
    wire N__11350;
    wire N__11347;
    wire N__11342;
    wire N__11339;
    wire N__11336;
    wire N__11333;
    wire N__11332;
    wire N__11331;
    wire N__11328;
    wire N__11325;
    wire N__11322;
    wire N__11315;
    wire N__11314;
    wire N__11311;
    wire N__11308;
    wire N__11305;
    wire N__11300;
    wire N__11297;
    wire N__11296;
    wire N__11293;
    wire N__11290;
    wire N__11287;
    wire N__11282;
    wire N__11279;
    wire N__11276;
    wire N__11275;
    wire N__11274;
    wire N__11273;
    wire N__11270;
    wire N__11267;
    wire N__11262;
    wire N__11255;
    wire N__11252;
    wire N__11249;
    wire N__11246;
    wire N__11245;
    wire N__11244;
    wire N__11243;
    wire N__11242;
    wire N__11231;
    wire N__11230;
    wire N__11229;
    wire N__11228;
    wire N__11225;
    wire N__11218;
    wire N__11217;
    wire N__11216;
    wire N__11211;
    wire N__11208;
    wire N__11205;
    wire N__11198;
    wire N__11195;
    wire N__11192;
    wire N__11189;
    wire N__11186;
    wire N__11183;
    wire N__11180;
    wire N__11179;
    wire N__11176;
    wire N__11173;
    wire N__11168;
    wire N__11167;
    wire N__11164;
    wire N__11161;
    wire N__11156;
    wire N__11155;
    wire N__11152;
    wire N__11151;
    wire N__11148;
    wire N__11145;
    wire N__11142;
    wire N__11139;
    wire N__11136;
    wire N__11131;
    wire N__11130;
    wire N__11129;
    wire N__11128;
    wire N__11123;
    wire N__11118;
    wire N__11115;
    wire N__11108;
    wire N__11105;
    wire N__11104;
    wire N__11103;
    wire N__11096;
    wire N__11093;
    wire N__11090;
    wire N__11087;
    wire N__11084;
    wire N__11081;
    wire N__11078;
    wire N__11077;
    wire N__11074;
    wire N__11071;
    wire N__11068;
    wire N__11063;
    wire N__11062;
    wire N__11059;
    wire N__11056;
    wire N__11051;
    wire N__11048;
    wire N__11045;
    wire N__11044;
    wire N__11041;
    wire N__11038;
    wire N__11033;
    wire N__11032;
    wire N__11029;
    wire N__11026;
    wire N__11023;
    wire N__11018;
    wire N__11017;
    wire N__11014;
    wire N__11011;
    wire N__11008;
    wire N__11003;
    wire N__11000;
    wire N__10997;
    wire N__10994;
    wire N__10993;
    wire N__10992;
    wire N__10989;
    wire N__10986;
    wire N__10983;
    wire N__10976;
    wire N__10975;
    wire N__10970;
    wire N__10967;
    wire N__10966;
    wire N__10963;
    wire N__10962;
    wire N__10961;
    wire N__10958;
    wire N__10955;
    wire N__10954;
    wire N__10951;
    wire N__10948;
    wire N__10943;
    wire N__10942;
    wire N__10939;
    wire N__10934;
    wire N__10931;
    wire N__10928;
    wire N__10925;
    wire N__10916;
    wire N__10913;
    wire N__10912;
    wire N__10909;
    wire N__10906;
    wire N__10901;
    wire N__10898;
    wire N__10895;
    wire N__10892;
    wire N__10889;
    wire N__10886;
    wire N__10883;
    wire N__10880;
    wire N__10877;
    wire N__10874;
    wire N__10871;
    wire N__10868;
    wire N__10865;
    wire N__10862;
    wire N__10859;
    wire N__10856;
    wire N__10853;
    wire N__10850;
    wire N__10847;
    wire N__10844;
    wire N__10841;
    wire N__10838;
    wire N__10835;
    wire N__10832;
    wire N__10829;
    wire N__10826;
    wire N__10823;
    wire N__10820;
    wire N__10817;
    wire N__10814;
    wire N__10811;
    wire N__10808;
    wire N__10805;
    wire N__10802;
    wire N__10799;
    wire N__10796;
    wire N__10793;
    wire N__10792;
    wire N__10789;
    wire N__10786;
    wire N__10781;
    wire N__10778;
    wire N__10775;
    wire N__10772;
    wire N__10769;
    wire N__10768;
    wire N__10765;
    wire N__10762;
    wire N__10757;
    wire N__10756;
    wire N__10751;
    wire N__10748;
    wire N__10745;
    wire N__10742;
    wire N__10739;
    wire N__10736;
    wire N__10733;
    wire N__10730;
    wire N__10727;
    wire N__10724;
    wire N__10723;
    wire N__10720;
    wire N__10717;
    wire N__10712;
    wire N__10711;
    wire N__10708;
    wire N__10705;
    wire N__10700;
    wire N__10699;
    wire N__10696;
    wire N__10693;
    wire N__10688;
    wire N__10687;
    wire N__10684;
    wire N__10681;
    wire N__10678;
    wire N__10673;
    wire N__10672;
    wire N__10669;
    wire N__10666;
    wire N__10663;
    wire N__10658;
    wire N__10657;
    wire N__10656;
    wire N__10653;
    wire N__10652;
    wire N__10649;
    wire N__10646;
    wire N__10643;
    wire N__10640;
    wire N__10637;
    wire N__10636;
    wire N__10633;
    wire N__10628;
    wire N__10625;
    wire N__10622;
    wire N__10613;
    wire N__10610;
    wire N__10609;
    wire N__10608;
    wire N__10607;
    wire N__10604;
    wire N__10601;
    wire N__10600;
    wire N__10597;
    wire N__10594;
    wire N__10593;
    wire N__10588;
    wire N__10585;
    wire N__10582;
    wire N__10579;
    wire N__10576;
    wire N__10571;
    wire N__10566;
    wire N__10563;
    wire N__10560;
    wire N__10555;
    wire N__10552;
    wire N__10549;
    wire N__10546;
    wire N__10543;
    wire N__10540;
    wire N__10537;
    wire N__10532;
    wire N__10531;
    wire N__10530;
    wire N__10527;
    wire N__10526;
    wire N__10525;
    wire N__10524;
    wire N__10523;
    wire N__10520;
    wire N__10517;
    wire N__10514;
    wire N__10511;
    wire N__10508;
    wire N__10503;
    wire N__10500;
    wire N__10499;
    wire N__10496;
    wire N__10491;
    wire N__10484;
    wire N__10481;
    wire N__10472;
    wire N__10469;
    wire N__10466;
    wire N__10463;
    wire N__10460;
    wire N__10457;
    wire N__10454;
    wire N__10451;
    wire N__10448;
    wire N__10445;
    wire N__10442;
    wire N__10441;
    wire N__10436;
    wire N__10433;
    wire N__10430;
    wire N__10427;
    wire N__10424;
    wire N__10421;
    wire N__10418;
    wire N__10417;
    wire N__10414;
    wire N__10411;
    wire N__10406;
    wire N__10405;
    wire N__10402;
    wire N__10399;
    wire N__10394;
    wire N__10393;
    wire N__10390;
    wire N__10387;
    wire N__10382;
    wire N__10379;
    wire N__10376;
    wire N__10373;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10361;
    wire N__10360;
    wire N__10357;
    wire N__10354;
    wire N__10349;
    wire N__10348;
    wire N__10345;
    wire N__10342;
    wire N__10337;
    wire N__10334;
    wire N__10333;
    wire N__10330;
    wire N__10327;
    wire N__10324;
    wire N__10319;
    wire N__10316;
    wire N__10313;
    wire N__10310;
    wire N__10307;
    wire N__10304;
    wire N__10303;
    wire N__10300;
    wire N__10297;
    wire N__10292;
    wire N__10291;
    wire N__10288;
    wire N__10285;
    wire N__10280;
    wire N__10279;
    wire N__10278;
    wire N__10277;
    wire N__10276;
    wire N__10275;
    wire N__10266;
    wire N__10265;
    wire N__10262;
    wire N__10259;
    wire N__10256;
    wire N__10253;
    wire N__10250;
    wire N__10247;
    wire N__10238;
    wire N__10235;
    wire N__10234;
    wire N__10229;
    wire N__10226;
    wire N__10225;
    wire N__10224;
    wire N__10217;
    wire N__10214;
    wire N__10213;
    wire N__10210;
    wire N__10207;
    wire N__10202;
    wire N__10199;
    wire N__10198;
    wire N__10197;
    wire N__10196;
    wire N__10191;
    wire N__10188;
    wire N__10185;
    wire N__10178;
    wire N__10175;
    wire N__10174;
    wire N__10173;
    wire N__10170;
    wire N__10167;
    wire N__10164;
    wire N__10163;
    wire N__10162;
    wire N__10161;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10151;
    wire N__10148;
    wire N__10147;
    wire N__10144;
    wire N__10143;
    wire N__10138;
    wire N__10135;
    wire N__10132;
    wire N__10127;
    wire N__10122;
    wire N__10119;
    wire N__10106;
    wire N__10103;
    wire N__10102;
    wire N__10099;
    wire N__10096;
    wire N__10093;
    wire N__10088;
    wire N__10087;
    wire N__10084;
    wire N__10081;
    wire N__10076;
    wire N__10075;
    wire N__10072;
    wire N__10069;
    wire N__10068;
    wire N__10065;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10057;
    wire N__10056;
    wire N__10055;
    wire N__10052;
    wire N__10049;
    wire N__10044;
    wire N__10041;
    wire N__10038;
    wire N__10035;
    wire N__10032;
    wire N__10029;
    wire N__10024;
    wire N__10021;
    wire N__10018;
    wire N__10015;
    wire N__10012;
    wire N__10009;
    wire N__10004;
    wire N__9995;
    wire N__9992;
    wire N__9989;
    wire N__9988;
    wire N__9985;
    wire N__9982;
    wire N__9977;
    wire N__9974;
    wire N__9971;
    wire N__9970;
    wire N__9967;
    wire N__9964;
    wire N__9959;
    wire N__9958;
    wire N__9957;
    wire N__9956;
    wire N__9955;
    wire N__9952;
    wire N__9947;
    wire N__9944;
    wire N__9941;
    wire N__9938;
    wire N__9929;
    wire N__9928;
    wire N__9927;
    wire N__9926;
    wire N__9925;
    wire N__9918;
    wire N__9915;
    wire N__9912;
    wire N__9905;
    wire N__9902;
    wire N__9899;
    wire N__9896;
    wire N__9893;
    wire N__9890;
    wire N__9887;
    wire N__9884;
    wire N__9881;
    wire N__9878;
    wire N__9875;
    wire N__9874;
    wire N__9873;
    wire N__9870;
    wire N__9865;
    wire N__9860;
    wire N__9857;
    wire N__9854;
    wire N__9851;
    wire N__9850;
    wire N__9849;
    wire N__9848;
    wire N__9845;
    wire N__9842;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9832;
    wire N__9829;
    wire N__9826;
    wire N__9823;
    wire N__9820;
    wire N__9817;
    wire N__9814;
    wire N__9803;
    wire N__9800;
    wire N__9797;
    wire N__9796;
    wire N__9793;
    wire N__9792;
    wire N__9789;
    wire N__9786;
    wire N__9783;
    wire N__9780;
    wire N__9773;
    wire N__9770;
    wire N__9767;
    wire N__9766;
    wire N__9763;
    wire N__9760;
    wire N__9757;
    wire N__9752;
    wire N__9749;
    wire N__9748;
    wire N__9743;
    wire N__9740;
    wire N__9737;
    wire N__9734;
    wire N__9731;
    wire N__9728;
    wire N__9725;
    wire N__9724;
    wire N__9721;
    wire N__9718;
    wire N__9713;
    wire N__9710;
    wire N__9709;
    wire N__9706;
    wire N__9703;
    wire N__9698;
    wire N__9695;
    wire N__9694;
    wire N__9691;
    wire N__9688;
    wire N__9683;
    wire N__9682;
    wire N__9679;
    wire N__9676;
    wire N__9671;
    wire N__9668;
    wire N__9667;
    wire N__9664;
    wire N__9661;
    wire N__9656;
    wire N__9655;
    wire N__9652;
    wire N__9649;
    wire N__9644;
    wire N__9641;
    wire N__9638;
    wire N__9635;
    wire N__9634;
    wire N__9631;
    wire N__9628;
    wire N__9623;
    wire N__9622;
    wire N__9619;
    wire N__9616;
    wire N__9611;
    wire N__9610;
    wire N__9607;
    wire N__9604;
    wire N__9599;
    wire N__9596;
    wire N__9593;
    wire N__9592;
    wire N__9591;
    wire N__9590;
    wire N__9589;
    wire N__9588;
    wire N__9587;
    wire N__9584;
    wire N__9581;
    wire N__9578;
    wire N__9571;
    wire N__9568;
    wire N__9565;
    wire N__9562;
    wire N__9551;
    wire N__9548;
    wire N__9545;
    wire N__9542;
    wire N__9539;
    wire N__9536;
    wire N__9535;
    wire N__9530;
    wire N__9527;
    wire N__9526;
    wire N__9523;
    wire N__9522;
    wire N__9519;
    wire N__9514;
    wire N__9509;
    wire N__9508;
    wire N__9507;
    wire N__9506;
    wire N__9501;
    wire N__9500;
    wire N__9499;
    wire N__9496;
    wire N__9493;
    wire N__9490;
    wire N__9489;
    wire N__9488;
    wire N__9487;
    wire N__9484;
    wire N__9481;
    wire N__9478;
    wire N__9475;
    wire N__9472;
    wire N__9465;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9443;
    wire N__9440;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9422;
    wire N__9419;
    wire N__9416;
    wire N__9415;
    wire N__9412;
    wire N__9409;
    wire N__9404;
    wire N__9403;
    wire N__9400;
    wire N__9397;
    wire N__9392;
    wire N__9389;
    wire N__9386;
    wire N__9383;
    wire N__9380;
    wire N__9377;
    wire N__9374;
    wire N__9371;
    wire N__9368;
    wire N__9365;
    wire N__9362;
    wire N__9359;
    wire N__9356;
    wire N__9353;
    wire N__9350;
    wire N__9349;
    wire N__9346;
    wire N__9341;
    wire N__9338;
    wire N__9335;
    wire N__9332;
    wire N__9329;
    wire N__9326;
    wire N__9323;
    wire N__9322;
    wire N__9319;
    wire N__9316;
    wire N__9311;
    wire N__9310;
    wire N__9307;
    wire N__9304;
    wire N__9303;
    wire N__9302;
    wire N__9299;
    wire N__9296;
    wire N__9295;
    wire N__9292;
    wire N__9289;
    wire N__9288;
    wire N__9283;
    wire N__9280;
    wire N__9275;
    wire N__9272;
    wire N__9263;
    wire N__9260;
    wire N__9259;
    wire N__9258;
    wire N__9257;
    wire N__9254;
    wire N__9253;
    wire N__9252;
    wire N__9251;
    wire N__9248;
    wire N__9243;
    wire N__9240;
    wire N__9239;
    wire N__9238;
    wire N__9237;
    wire N__9232;
    wire N__9227;
    wire N__9222;
    wire N__9219;
    wire N__9214;
    wire N__9203;
    wire N__9202;
    wire N__9197;
    wire N__9194;
    wire N__9191;
    wire N__9188;
    wire N__9187;
    wire N__9184;
    wire N__9183;
    wire N__9180;
    wire N__9179;
    wire N__9174;
    wire N__9171;
    wire N__9168;
    wire N__9161;
    wire N__9160;
    wire N__9159;
    wire N__9156;
    wire N__9155;
    wire N__9150;
    wire N__9147;
    wire N__9144;
    wire N__9137;
    wire N__9134;
    wire N__9131;
    wire N__9128;
    wire N__9127;
    wire N__9124;
    wire N__9121;
    wire N__9116;
    wire N__9113;
    wire N__9110;
    wire N__9107;
    wire N__9104;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9092;
    wire N__9089;
    wire N__9086;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9076;
    wire N__9075;
    wire N__9074;
    wire N__9073;
    wire N__9072;
    wire N__9071;
    wire N__9066;
    wire N__9061;
    wire N__9056;
    wire N__9053;
    wire N__9044;
    wire N__9041;
    wire N__9038;
    wire N__9035;
    wire N__9032;
    wire N__9031;
    wire N__9028;
    wire N__9025;
    wire N__9020;
    wire N__9017;
    wire N__9014;
    wire N__9011;
    wire N__9008;
    wire N__9005;
    wire N__9002;
    wire N__8999;
    wire N__8996;
    wire N__8995;
    wire N__8992;
    wire N__8989;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8975;
    wire N__8972;
    wire N__8969;
    wire N__8966;
    wire N__8965;
    wire N__8962;
    wire N__8959;
    wire N__8954;
    wire N__8951;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8941;
    wire N__8938;
    wire N__8935;
    wire N__8930;
    wire N__8927;
    wire N__8924;
    wire N__8921;
    wire N__8918;
    wire N__8917;
    wire N__8914;
    wire N__8911;
    wire N__8906;
    wire N__8903;
    wire N__8900;
    wire N__8897;
    wire N__8894;
    wire N__8891;
    wire N__8890;
    wire N__8887;
    wire N__8884;
    wire N__8879;
    wire N__8876;
    wire N__8873;
    wire N__8870;
    wire N__8869;
    wire N__8866;
    wire N__8863;
    wire N__8858;
    wire N__8855;
    wire N__8852;
    wire N__8849;
    wire N__8846;
    wire N__8843;
    wire N__8840;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8828;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8807;
    wire N__8806;
    wire N__8803;
    wire N__8800;
    wire N__8795;
    wire N__8792;
    wire N__8789;
    wire N__8786;
    wire N__8783;
    wire N__8780;
    wire N__8777;
    wire N__8776;
    wire N__8775;
    wire N__8772;
    wire N__8767;
    wire N__8762;
    wire N__8759;
    wire N__8756;
    wire N__8753;
    wire N__8750;
    wire N__8747;
    wire N__8744;
    wire N__8743;
    wire N__8742;
    wire N__8739;
    wire N__8736;
    wire N__8733;
    wire N__8730;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8713;
    wire N__8712;
    wire N__8709;
    wire N__8706;
    wire N__8703;
    wire N__8696;
    wire N__8693;
    wire N__8692;
    wire N__8689;
    wire N__8686;
    wire N__8685;
    wire N__8682;
    wire N__8679;
    wire N__8676;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8662;
    wire N__8661;
    wire N__8658;
    wire N__8655;
    wire N__8652;
    wire N__8645;
    wire N__8644;
    wire N__8641;
    wire N__8638;
    wire N__8635;
    wire N__8632;
    wire N__8629;
    wire N__8626;
    wire N__8623;
    wire N__8620;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8602;
    wire N__8599;
    wire N__8596;
    wire N__8593;
    wire N__8590;
    wire N__8585;
    wire N__8584;
    wire N__8583;
    wire N__8582;
    wire N__8581;
    wire N__8580;
    wire N__8579;
    wire N__8576;
    wire N__8575;
    wire N__8574;
    wire N__8563;
    wire N__8562;
    wire N__8559;
    wire N__8556;
    wire N__8551;
    wire N__8548;
    wire N__8545;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8525;
    wire N__8522;
    wire N__8519;
    wire N__8516;
    wire N__8515;
    wire N__8514;
    wire N__8511;
    wire N__8510;
    wire N__8509;
    wire N__8506;
    wire N__8505;
    wire N__8502;
    wire N__8499;
    wire N__8496;
    wire N__8493;
    wire N__8492;
    wire N__8491;
    wire N__8488;
    wire N__8485;
    wire N__8480;
    wire N__8477;
    wire N__8476;
    wire N__8475;
    wire N__8470;
    wire N__8467;
    wire N__8462;
    wire N__8457;
    wire N__8454;
    wire N__8451;
    wire N__8448;
    wire N__8445;
    wire N__8440;
    wire N__8429;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8419;
    wire N__8414;
    wire N__8411;
    wire N__8410;
    wire N__8409;
    wire N__8408;
    wire N__8407;
    wire N__8404;
    wire N__8401;
    wire N__8394;
    wire N__8387;
    wire N__8386;
    wire N__8383;
    wire N__8382;
    wire N__8381;
    wire N__8378;
    wire N__8375;
    wire N__8370;
    wire N__8367;
    wire N__8360;
    wire N__8357;
    wire N__8356;
    wire N__8355;
    wire N__8352;
    wire N__8351;
    wire N__8350;
    wire N__8349;
    wire N__8346;
    wire N__8343;
    wire N__8340;
    wire N__8337;
    wire N__8332;
    wire N__8321;
    wire N__8318;
    wire N__8317;
    wire N__8316;
    wire N__8315;
    wire N__8314;
    wire N__8311;
    wire N__8308;
    wire N__8305;
    wire N__8302;
    wire N__8301;
    wire N__8300;
    wire N__8297;
    wire N__8292;
    wire N__8289;
    wire N__8286;
    wire N__8283;
    wire N__8280;
    wire N__8267;
    wire N__8264;
    wire N__8261;
    wire N__8258;
    wire N__8257;
    wire N__8256;
    wire N__8253;
    wire N__8248;
    wire N__8245;
    wire N__8240;
    wire N__8237;
    wire N__8236;
    wire N__8235;
    wire N__8232;
    wire N__8227;
    wire N__8222;
    wire N__8221;
    wire N__8220;
    wire N__8217;
    wire N__8214;
    wire N__8211;
    wire N__8204;
    wire N__8201;
    wire N__8200;
    wire N__8199;
    wire N__8196;
    wire N__8193;
    wire N__8190;
    wire N__8183;
    wire N__8180;
    wire N__8179;
    wire N__8176;
    wire N__8175;
    wire N__8172;
    wire N__8167;
    wire N__8162;
    wire N__8159;
    wire N__8156;
    wire N__8153;
    wire N__8150;
    wire N__8147;
    wire N__8146;
    wire N__8143;
    wire N__8140;
    wire N__8137;
    wire N__8134;
    wire N__8133;
    wire N__8130;
    wire N__8127;
    wire N__8124;
    wire N__8117;
    wire N__8116;
    wire N__8113;
    wire N__8110;
    wire N__8107;
    wire N__8104;
    wire N__8103;
    wire N__8098;
    wire N__8095;
    wire N__8090;
    wire N__8087;
    wire N__8084;
    wire N__8081;
    wire N__8078;
    wire N__8077;
    wire N__8074;
    wire N__8071;
    wire N__8068;
    wire N__8067;
    wire N__8064;
    wire N__8061;
    wire N__8058;
    wire N__8051;
    wire N__8048;
    wire N__8045;
    wire N__8042;
    wire N__8039;
    wire N__8036;
    wire N__8035;
    wire N__8034;
    wire N__8031;
    wire N__8026;
    wire N__8021;
    wire N__8018;
    wire N__8015;
    wire N__8014;
    wire N__8011;
    wire N__8008;
    wire N__8005;
    wire N__8002;
    wire N__7999;
    wire N__7996;
    wire N__7993;
    wire N__7990;
    wire N__7989;
    wire N__7986;
    wire N__7983;
    wire N__7980;
    wire N__7973;
    wire N__7970;
    wire N__7967;
    wire N__7966;
    wire N__7963;
    wire N__7960;
    wire N__7955;
    wire N__7952;
    wire N__7951;
    wire N__7948;
    wire N__7945;
    wire N__7942;
    wire N__7939;
    wire N__7934;
    wire N__7931;
    wire N__7928;
    wire N__7927;
    wire N__7924;
    wire N__7923;
    wire N__7920;
    wire N__7919;
    wire N__7918;
    wire N__7915;
    wire N__7912;
    wire N__7909;
    wire N__7906;
    wire N__7903;
    wire N__7900;
    wire N__7897;
    wire N__7894;
    wire N__7891;
    wire N__7886;
    wire N__7877;
    wire N__7874;
    wire N__7873;
    wire N__7870;
    wire N__7867;
    wire N__7866;
    wire N__7863;
    wire N__7860;
    wire N__7857;
    wire N__7854;
    wire N__7847;
    wire N__7844;
    wire N__7841;
    wire N__7838;
    wire N__7837;
    wire N__7834;
    wire N__7831;
    wire N__7826;
    wire N__7825;
    wire N__7820;
    wire N__7819;
    wire N__7816;
    wire N__7815;
    wire N__7814;
    wire N__7813;
    wire N__7810;
    wire N__7807;
    wire N__7804;
    wire N__7799;
    wire N__7796;
    wire N__7787;
    wire N__7786;
    wire N__7785;
    wire N__7780;
    wire N__7777;
    wire N__7774;
    wire N__7773;
    wire N__7772;
    wire N__7771;
    wire N__7770;
    wire N__7769;
    wire N__7766;
    wire N__7763;
    wire N__7758;
    wire N__7753;
    wire N__7750;
    wire N__7739;
    wire N__7736;
    wire N__7735;
    wire N__7734;
    wire N__7731;
    wire N__7726;
    wire N__7721;
    wire N__7720;
    wire N__7719;
    wire N__7718;
    wire N__7717;
    wire N__7712;
    wire N__7711;
    wire N__7710;
    wire N__7709;
    wire N__7706;
    wire N__7701;
    wire N__7698;
    wire N__7695;
    wire N__7690;
    wire N__7679;
    wire N__7676;
    wire N__7673;
    wire N__7670;
    wire N__7667;
    wire N__7664;
    wire N__7661;
    wire N__7658;
    wire N__7655;
    wire N__7652;
    wire N__7649;
    wire N__7646;
    wire N__7643;
    wire N__7640;
    wire N__7637;
    wire N__7634;
    wire N__7631;
    wire N__7628;
    wire N__7625;
    wire N__7622;
    wire N__7619;
    wire N__7616;
    wire N__7613;
    wire N__7610;
    wire N__7607;
    wire N__7606;
    wire N__7603;
    wire N__7600;
    wire N__7595;
    wire N__7592;
    wire N__7589;
    wire N__7586;
    wire N__7583;
    wire N__7580;
    wire N__7577;
    wire N__7574;
    wire N__7571;
    wire N__7568;
    wire N__7567;
    wire N__7564;
    wire N__7563;
    wire N__7560;
    wire N__7557;
    wire N__7554;
    wire N__7547;
    wire N__7544;
    wire N__7541;
    wire N__7538;
    wire N__7535;
    wire N__7532;
    wire N__7529;
    wire N__7526;
    wire N__7523;
    wire N__7520;
    wire N__7517;
    wire N__7514;
    wire N__7511;
    wire N__7508;
    wire N__7505;
    wire N__7502;
    wire N__7499;
    wire N__7496;
    wire N__7493;
    wire N__7490;
    wire N__7487;
    wire N__7484;
    wire N__7481;
    wire N__7478;
    wire N__7475;
    wire N__7472;
    wire N__7469;
    wire N__7466;
    wire N__7463;
    wire N__7460;
    wire N__7457;
    wire N__7454;
    wire N__7451;
    wire N__7448;
    wire N__7445;
    wire N__7442;
    wire N__7439;
    wire N__7436;
    wire N__7435;
    wire N__7432;
    wire N__7431;
    wire N__7428;
    wire N__7425;
    wire N__7422;
    wire N__7415;
    wire N__7412;
    wire N__7409;
    wire N__7406;
    wire N__7405;
    wire N__7402;
    wire N__7401;
    wire N__7398;
    wire N__7395;
    wire N__7392;
    wire N__7385;
    wire N__7382;
    wire N__7379;
    wire N__7376;
    wire N__7375;
    wire N__7372;
    wire N__7371;
    wire N__7368;
    wire N__7365;
    wire N__7362;
    wire N__7355;
    wire N__7352;
    wire N__7349;
    wire N__7346;
    wire N__7343;
    wire N__7340;
    wire N__7339;
    wire N__7338;
    wire N__7335;
    wire N__7332;
    wire N__7329;
    wire N__7322;
    wire N__7319;
    wire N__7316;
    wire N__7313;
    wire N__7310;
    wire N__7309;
    wire N__7306;
    wire N__7303;
    wire N__7298;
    wire N__7295;
    wire N__7292;
    wire N__7289;
    wire N__7286;
    wire N__7283;
    wire N__7280;
    wire N__7277;
    wire N__7274;
    wire N__7271;
    wire N__7270;
    wire N__7267;
    wire N__7264;
    wire N__7263;
    wire N__7258;
    wire N__7255;
    wire N__7250;
    wire N__7247;
    wire N__7244;
    wire N__7241;
    wire N__7238;
    wire N__7235;
    wire N__7232;
    wire N__7229;
    wire N__7226;
    wire N__7223;
    wire N__7220;
    wire N__7217;
    wire N__7214;
    wire N__7211;
    wire N__7208;
    wire N__7205;
    wire N__7202;
    wire N__7199;
    wire N__7196;
    wire N__7193;
    wire N__7190;
    wire N__7187;
    wire N__7184;
    wire N__7183;
    wire N__7178;
    wire N__7175;
    wire N__7172;
    wire N__7169;
    wire N__7166;
    wire N__7163;
    wire N__7160;
    wire N__7157;
    wire N__7154;
    wire N__7151;
    wire N__7148;
    wire N__7145;
    wire N__7142;
    wire N__7139;
    wire N__7136;
    wire N__7135;
    wire N__7132;
    wire N__7131;
    wire N__7128;
    wire N__7125;
    wire N__7122;
    wire N__7119;
    wire N__7112;
    wire N__7109;
    wire N__7106;
    wire N__7103;
    wire N__7102;
    wire N__7101;
    wire N__7098;
    wire N__7095;
    wire N__7092;
    wire N__7085;
    wire N__7082;
    wire N__7079;
    wire N__7078;
    wire N__7075;
    wire N__7074;
    wire N__7071;
    wire N__7068;
    wire N__7065;
    wire N__7058;
    wire N__7055;
    wire N__7052;
    wire N__7049;
    wire N__7046;
    wire N__7045;
    wire N__7042;
    wire N__7039;
    wire N__7038;
    wire N__7035;
    wire N__7032;
    wire N__7029;
    wire N__7026;
    wire N__7023;
    wire N__7016;
    wire N__7013;
    wire N__7010;
    wire N__7007;
    wire N__7004;
    wire N__7001;
    wire N__6998;
    wire N__6995;
    wire N__6994;
    wire N__6991;
    wire N__6988;
    wire N__6983;
    wire N__6980;
    wire N__6977;
    wire N__6974;
    wire N__6971;
    wire N__6970;
    wire N__6969;
    wire N__6966;
    wire N__6963;
    wire N__6960;
    wire N__6953;
    wire N__6950;
    wire N__6947;
    wire N__6944;
    wire N__6941;
    wire N__6940;
    wire N__6939;
    wire N__6936;
    wire N__6933;
    wire N__6930;
    wire N__6923;
    wire N__6920;
    wire N__6917;
    wire N__6914;
    wire N__6911;
    wire N__6910;
    wire N__6909;
    wire N__6906;
    wire N__6903;
    wire N__6900;
    wire N__6893;
    wire N__6890;
    wire N__6887;
    wire N__6884;
    wire N__6881;
    wire N__6880;
    wire N__6879;
    wire N__6876;
    wire N__6873;
    wire N__6870;
    wire N__6863;
    wire N__6860;
    wire N__6857;
    wire N__6854;
    wire N__6851;
    wire N__6850;
    wire N__6847;
    wire N__6844;
    wire N__6843;
    wire N__6840;
    wire N__6837;
    wire N__6834;
    wire N__6829;
    wire N__6824;
    wire N__6821;
    wire N__6820;
    wire N__6817;
    wire N__6814;
    wire N__6811;
    wire N__6808;
    wire N__6805;
    wire N__6802;
    wire N__6801;
    wire N__6798;
    wire N__6795;
    wire N__6792;
    wire N__6785;
    wire N__6782;
    wire N__6779;
    wire N__6776;
    wire N__6775;
    wire N__6772;
    wire N__6769;
    wire N__6764;
    wire N__6761;
    wire N__6758;
    wire N__6755;
    wire N__6752;
    wire N__6749;
    wire N__6746;
    wire N__6743;
    wire N__6740;
    wire N__6737;
    wire N__6736;
    wire N__6733;
    wire N__6730;
    wire N__6725;
    wire N__6724;
    wire N__6721;
    wire N__6718;
    wire N__6713;
    wire N__6712;
    wire N__6709;
    wire N__6706;
    wire N__6703;
    wire N__6698;
    wire N__6697;
    wire N__6694;
    wire N__6691;
    wire N__6686;
    wire N__6683;
    wire N__6680;
    wire N__6679;
    wire N__6678;
    wire N__6675;
    wire N__6672;
    wire N__6669;
    wire N__6662;
    wire N__6661;
    wire N__6660;
    wire N__6657;
    wire N__6654;
    wire N__6651;
    wire N__6644;
    wire N__6641;
    wire N__6638;
    wire N__6635;
    wire N__6632;
    wire N__6629;
    wire N__6626;
    wire N__6625;
    wire N__6622;
    wire N__6619;
    wire N__6614;
    wire N__6613;
    wire N__6610;
    wire N__6607;
    wire N__6602;
    wire N__6601;
    wire N__6598;
    wire N__6595;
    wire N__6592;
    wire N__6587;
    wire N__6586;
    wire N__6583;
    wire N__6580;
    wire N__6575;
    wire N__6572;
    wire N__6571;
    wire N__6568;
    wire N__6565;
    wire N__6560;
    wire N__6559;
    wire N__6556;
    wire N__6553;
    wire N__6550;
    wire N__6545;
    wire N__6542;
    wire N__6541;
    wire N__6538;
    wire N__6535;
    wire N__6530;
    wire N__6527;
    wire N__6526;
    wire N__6523;
    wire N__6520;
    wire N__6515;
    wire N__6514;
    wire N__6511;
    wire N__6508;
    wire N__6503;
    wire N__6502;
    wire N__6499;
    wire N__6496;
    wire N__6491;
    wire N__6488;
    wire N__6485;
    wire N__6482;
    wire N__6479;
    wire N__6476;
    wire N__6473;
    wire N__6470;
    wire N__6467;
    wire N__6464;
    wire N__6461;
    wire N__6458;
    wire N__6455;
    wire N__6452;
    wire N__6449;
    wire \INVfifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net ;
    wire \INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net ;
    wire BTN_N_c;
    wire \INVfifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net ;
    wire \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net ;
    wire VCCG0;
    wire GNDG0;
    wire \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO ;
    wire bfn_9_14_0_;
    wire \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_0 ;
    wire \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_1 ;
    wire \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_2 ;
    wire \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_3 ;
    wire \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_4 ;
    wire \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_5 ;
    wire \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_6 ;
    wire \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_7 ;
    wire bfn_9_15_0_;
    wire \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_8 ;
    wire \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_9 ;
    wire \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_10 ;
    wire \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_11 ;
    wire \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_12 ;
    wire \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_13 ;
    wire \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_8 ;
    wire \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_7 ;
    wire \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_14 ;
    wire \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_10 ;
    wire \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_11 ;
    wire \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_12 ;
    wire \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_9 ;
    wire \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_13 ;
    wire \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_6 ;
    wire \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_5 ;
    wire \uart_inst0.uart_inst0.un1_rx_clk_divider_10 ;
    wire \uart_inst0.uart_inst0.un1_rx_clk_divider_9 ;
    wire \uart_inst0.uart_inst0.un1_rx_clk_divider_7_cascade_ ;
    wire \uart_inst0.uart_inst0.un1_rx_clk_divider_0_cascade_ ;
    wire \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_3 ;
    wire \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_1 ;
    wire \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_4 ;
    wire \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_2 ;
    wire \uart_inst0.uart_inst0.un1_rx_clk_divider_8 ;
    wire \uart_inst0.uart_inst0.rx_clk_dividerZ0Z_0 ;
    wire \uart_inst0.uart_inst0.rx_clk_divider_1_sqmuxa_i ;
    wire P1A3_c;
    wire N_86_mux;
    wire \uart_inst0.tx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_0_cascade_ ;
    wire \uart_inst0.tx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_6 ;
    wire GB_BUFFER_wPllLocked_i_g_THRU_CO;
    wire fifo_inst_tx_fifo_inst_wRamWrEn_cascade_;
    wire \uart_inst0.tx_uart_fifo_inst.m68_eZ0Z_5_cascade_ ;
    wire \uart_inst0.tx_uart_fifo_inst.m68_eZ0Z_6 ;
    wire \uart_inst0.tx_uart_fifo_inst.N_92 ;
    wire fifo_inst_tx_fifo_inst_rRamWrAddr_0;
    wire rRamWrAddr_RNI10581_0;
    wire bfn_13_2_0_;
    wire fifo_inst_tx_fifo_inst_rRamWrAddr_1;
    wire \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_0 ;
    wire fifo_inst_tx_fifo_inst_rRamWrAddr_2;
    wire \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_1 ;
    wire fifo_inst_tx_fifo_inst_rRamWrAddr_3;
    wire un1_rRamWrAddr_cry_2_c_RNISJKU;
    wire \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_2 ;
    wire fifo_inst_tx_fifo_inst_rRamWrAddr_4;
    wire \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_3 ;
    wire fifo_inst_tx_fifo_inst_rRamWrAddr_5;
    wire \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_4 ;
    wire fifo_inst_tx_fifo_inst_rRamWrAddr_6;
    wire \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_5 ;
    wire fifo_inst_tx_fifo_inst_rRamWrAddr_7;
    wire \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_6 ;
    wire \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_7 ;
    wire bfn_13_3_0_;
    wire fifo_inst_tx_fifo_inst_rRamWrAddr_8;
    wire fifo_inst_ft2232h_inst_un1_rFifoState_12_0_i_cascade_;
    wire \fifo_inst.tx_fifo_inst.un1_rDataCount_ac0_1_a1_1 ;
    wire \uart_inst0.tx_uart_fifo_inst.m78_bmZ0 ;
    wire \uart_inst0.tx_uart_fifo_inst.m78_nsZ0Z_1_cascade_ ;
    wire \fifo_inst.ft2232h_inst.un1_rFifoState_12_0_i_0 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c2_d_cascade_ ;
    wire N_84_mux_cascade_;
    wire \uart_inst0.tx_uart_fifo_inst.m65_bmZ0_cascade_ ;
    wire \fifo_inst.rx_fifo_inst.un1_rDataCount_c2_1_1_0_cascade_ ;
    wire \uart_inst0.tx_uart_fifo_inst.m65_nsZ0Z_1 ;
    wire \fifo_inst.rx_fifo_inst.un1_rDataCount_c2_1 ;
    wire fifo_inst_rx_fifo_inst_rDataCount_0_sqmuxa;
    wire \fifo_inst.rx_fifo_inst.un1_rDataCount_ac0_2 ;
    wire rUartTxEnZ0;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c3_0_0 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c2_d ;
    wire \uart_inst0.tx_uart_fifo_inst.rDataCount_0_sqmuxa ;
    wire \uart_inst0.wTxRdEmpty_cascade_ ;
    wire \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_0 ;
    wire \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_1 ;
    wire \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_2 ;
    wire \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_3 ;
    wire \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_4 ;
    wire \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_5 ;
    wire \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_6 ;
    wire \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_7 ;
    wire \INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net ;
    wire \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ1Z_0 ;
    wire \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNO_0Z0Z_0 ;
    wire bfn_13_12_0_;
    wire \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ1Z_1 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_0 ;
    wire \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ0Z_2 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_1 ;
    wire \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_3 ;
    wire \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNO_0Z0Z_3 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_2 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_3 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_4 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_5 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_6 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_7 ;
    wire bfn_13_13_0_;
    wire \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_8 ;
    wire \uart_inst0.wTxRdData_0 ;
    wire \uart_inst0.wTxRdData_1 ;
    wire \uart_inst0.uart_inst0.rTxDataZ0Z_1 ;
    wire \uart_inst0.wTxRdData_6 ;
    wire \uart_inst0.wTxRdData_3 ;
    wire \uart_inst0.wTxRdData_4 ;
    wire \uart_inst0.uart_inst0.rTxDataZ0Z_4 ;
    wire \uart_inst0.uart_inst0.rTxDataZ0Z_3 ;
    wire \uart_inst0.wTxRdData_2 ;
    wire \uart_inst0.uart_inst0.rTxDataZ0Z_2 ;
    wire \uart_inst0.uart_inst0.rTxDataZ0Z_6 ;
    wire \uart_inst0.wTxRdData_5 ;
    wire \uart_inst0.uart_inst0.rTxDataZ0Z_5 ;
    wire \uart_inst0.wTxRdData_7 ;
    wire \uart_inst0.uart_inst0.rTxDataZ0Z_7 ;
    wire N_97_cascade_;
    wire \uart_inst0.tx_uart_fifo_inst.m8_xZ0Z0_cascade_ ;
    wire \fifo_inst.tx_fifo_inst.un1_rDataCount_axbxc3_2_tz ;
    wire \fifo_inst.tx_fifo_inst.un1_rDataCount_axbxc3_a0_2 ;
    wire \fifo_inst.tx_fifo_inst.un1_rDataCount_c2_0 ;
    wire fifo_inst_tx_fifo_inst_wRamWrEn;
    wire \fifo_inst.tx_fifo_inst.un1_rDataCount_ac0_1_a0_0 ;
    wire \fifo_inst.tx_fifo_inst.un1_rDataCount_c2_1_cascade_ ;
    wire \fifo_inst.tx_fifo_inst.un1_rDataCount_ac0_2 ;
    wire fifo_inst_tx_fifo_inst_un1_rDataCount15_2_0_0;
    wire fifo_inst_tx_fifo_inst_rDataCount_2;
    wire fifo_inst_tx_fifo_inst_rDataCount_1;
    wire fifo_inst_tx_fifo_inst_rDataCount_fast_3;
    wire fifo_inst_tx_fifo_inst_rDataCount_0;
    wire \fifo_inst.rx_fifo_inst.un1_rDataCount_axbxc3_1_1_cascade_ ;
    wire \uart_inst0.tx_uart_fifo_inst.m15_xZ0Z0_cascade_ ;
    wire \fifo_inst.rx_fifo_inst.un1_rDataCount_axbxc3_1_1 ;
    wire fifo_inst_rx_fifo_inst_rDataCount_fast_3;
    wire P1A4_c;
    wire fifo_inst_ft2232h_inst_rFifoState_3;
    wire fifo_inst_rx_fifo_inst_un1_rDataCount15_2_0_0;
    wire fifo_inst_rx_fifo_inst_rDataCount_fast_0;
    wire N_84_mux;
    wire rUartTxEn_4_cascade_;
    wire rFtdiRxStateZ0Z_0;
    wire \fifo_inst.ft2232h_inst.rFifoStatesr_0 ;
    wire \fifo_inst.ft2232h_inst.rFifoStateZ0Z_2 ;
    wire iRxF_n_c;
    wire fifo_inst_ft2232h_inst_rFifoState_0;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c2 ;
    wire \uart_inst0.tx_uart_fifo_inst.wRamWrEn_1 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rDataCount_axbxc1_0 ;
    wire \uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_1 ;
    wire \uart_inst0.tx_uart_fifo_inst.rDataCountZ0Z_2 ;
    wire \uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_0 ;
    wire \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIJHQM1Z0Z_2_cascade_ ;
    wire \uart_inst0.tx_uart_fifo_inst.wUartTxFull ;
    wire bfn_14_11_0_;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_0 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_1 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_2 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_3 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_4 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_5 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_6 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_7 ;
    wire bfn_14_12_0_;
    wire \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_7 ;
    wire \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_5 ;
    wire \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_6 ;
    wire \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_4 ;
    wire \uart_inst0.tx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_5 ;
    wire P1A7_c;
    wire \uart_inst0.uart_inst0.tx_state_81_d ;
    wire \uart_inst0.uart_inst0.rTxDataZ0Z_0 ;
    wire \uart_inst0.uart_inst0.rTx_6_f1_0 ;
    wire \uart_inst0.uart_inst0.N_141_0 ;
    wire \uart_inst0.uart_inst0.N_143_0 ;
    wire \uart_inst0.uart_inst0.N_143_0_cascade_ ;
    wire \uart_inst0.uart_inst0.N_143_0_0 ;
    wire \uart_inst0.uart_inst0.un1_m3_0_a2_2_1 ;
    wire \uart_inst0.uart_inst0.N_136_0_cascade_ ;
    wire \uart_inst0.uart_inst0.un1_tx_bits_remaining_c1 ;
    wire \uart_inst0.uart_inst0.N_136_0 ;
    wire \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_0 ;
    wire wTxRdData_0;
    wire \INVfifo_inst.tx_fifo_inst.ram512x8_inst.RDATA_0C_net ;
    wire bfn_15_3_0_;
    wire \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_0 ;
    wire \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_1 ;
    wire \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_2 ;
    wire \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_3 ;
    wire \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIMJ1QZ0 ;
    wire \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_4 ;
    wire \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIOM2QZ0 ;
    wire \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_5 ;
    wire \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIQP3QZ0 ;
    wire \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_6 ;
    wire \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_7 ;
    wire bfn_15_4_0_;
    wire \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIE7TPZ0 ;
    wire \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNISS4QZ0 ;
    wire fifo_inst_wRxWrEn;
    wire bfn_15_5_0_;
    wire \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_0 ;
    wire \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNICK0CZ0 ;
    wire \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_1 ;
    wire \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_2 ;
    wire \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_3 ;
    wire \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_4 ;
    wire \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIK05CZ0 ;
    wire \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_5 ;
    wire \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_6 ;
    wire \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_7 ;
    wire bfn_15_6_0_;
    wire \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIIT3CZ0 ;
    wire rTxEnZ0;
    wire fifo_inst_wTxRdEn;
    wire fifo_inst_tx_fifo_inst_rDataCount_0_sqmuxa;
    wire fifo_inst_ft2232h_inst_rWrDelay;
    wire fifo_inst_ft2232h_inst_rFifoState_4;
    wire \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNIO67CZ0 ;
    wire rUartTxDataZ0Z_6;
    wire rUartTxDataZ0Z_5;
    wire rUartTxDataZ0Z_1;
    wire rUartRxDataZ0Z_5;
    wire rUartRxDataZ0Z_6;
    wire rUartRxDataZ0Z_1;
    wire \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_2 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNISGZ0Z74 ;
    wire \uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_5_cascade_ ;
    wire \uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7_cascade_ ;
    wire \uart_inst0.tx_uart_fifo_inst.wRamRdEn_1 ;
    wire \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0 ;
    wire \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIBDOK2Z0Z_0 ;
    wire \uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7 ;
    wire \uart_inst0.wTxRdEn_0 ;
    wire \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_5 ;
    wire \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_6 ;
    wire \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_7 ;
    wire \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_0 ;
    wire \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_3 ;
    wire \uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_4 ;
    wire \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_3 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIUJZ0Z84 ;
    wire \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_4 ;
    wire \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_5 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNI2QAZ0Z4 ;
    wire \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_6 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI4TBZ0Z4 ;
    wire \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_7 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI60DZ0Z4 ;
    wire \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_8 ;
    wire \uart_inst0.uart_inst0.rx_state_srsts_0_o2_3_3_cascade_ ;
    wire \uart_inst0.uart_inst0.N_257_0_cascade_ ;
    wire \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_2 ;
    wire \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_3 ;
    wire \uart_inst0.uart_inst0.N_157 ;
    wire \uart_inst0.uart_inst0.N_157_cascade_ ;
    wire \uart_inst0.uart_inst0.N_147_0_cascade_ ;
    wire \uart_inst0.uart_inst0.N_277_cascade_ ;
    wire \uart_inst0.uart_inst0.rx_state_srsts_0_a5_1_0 ;
    wire \uart_inst0.uart_inst0.N_280_cascade_ ;
    wire \uart_inst0.uart_inst0.rx_stateZ0Z_4 ;
    wire \uart_inst0.uart_inst0.N_261_0 ;
    wire \uart_inst0.wTxRdEmpty ;
    wire \uart_inst0.uart_inst0.tx_state_ns_0_0_0_cascade_ ;
    wire \uart_inst0.uart_inst0.tx_state_1_sqmuxa_1_0_a3_0 ;
    wire \uart_inst0.uart_inst0.tx_state_RNI1319Z0Z_0 ;
    wire \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_1 ;
    wire \uart_inst0.uart_inst0.tx_bits_remainingZ0Z_0 ;
    wire \uart_inst0.uart_inst0.un1_tx_bits_remaining_ac0_1_a0_0_cascade_ ;
    wire \uart_inst0.uart_inst0.un1_tx_bits_remaining_ac0_1 ;
    wire \uart_inst0.uart_inst0.un1_rx_state49_i_cascade_ ;
    wire \uart_inst0.uart_inst0.tx_countdown_RNO_0Z0Z_3_cascade_ ;
    wire \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_11_3_cascade_ ;
    wire \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13 ;
    wire wTxFull;
    wire rTxDataZ0Z_0;
    wire rTxBusReady;
    wire un1_rRamRdAddr_cry_2_c_RNIMVKN;
    wire m74;
    wire fifo_inst_tx_fifo_inst_rRamRdAddr_5;
    wire fifo_inst_tx_fifo_inst_rRamRdAddr_7;
    wire fifo_inst_tx_fifo_inst_rRamRdAddr_6;
    wire \uart_inst0.tx_uart_fifo_inst.m72_eZ0Z_5_cascade_ ;
    wire \uart_inst0.tx_uart_fifo_inst.N_100_cascade_ ;
    wire m73;
    wire fifo_inst_tx_fifo_inst_rRamRdAddr_3;
    wire fifo_inst_tx_fifo_inst_rRamRdAddr_1;
    wire fifo_inst_tx_fifo_inst_rRamRdAddr_8;
    wire \uart_inst0.tx_uart_fifo_inst.m72_eZ0Z_6 ;
    wire \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIKG0QZ0 ;
    wire fifo_inst_tx_fifo_inst_rRamRdAddr_4;
    wire fifo_inst_tx_fifo_inst_wRamRdEn;
    wire rRamRdAddr_RNI9KL42_0;
    wire \uart_inst0.tx_uart_fifo_inst.N_100 ;
    wire fifo_inst_tx_fifo_inst_rRamRdAddr_0;
    wire \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIM36CZ0 ;
    wire \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIAHVBZ0 ;
    wire un1_rRamRdAddr_cry_2_c_RNII9N9;
    wire m60;
    wire \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIGQ2CZ0 ;
    wire fifo_inst_rx_fifo_inst_rRamRdAddr_3;
    wire fifo_inst_rx_fifo_inst_rRamRdAddr_1;
    wire fifo_inst_rx_fifo_inst_rRamRdAddr_8;
    wire N_101;
    wire N_97;
    wire iTxE_n_c;
    wire N_8_0;
    wire fifo_inst_ft2232h_inst_un1_rFifoState_1_sqmuxa_0_i_cascade_;
    wire \fifo_inst.ft2232h_inst.un1_rFifoState_1_sqmuxa_0_i_0 ;
    wire m59;
    wire fifo_inst_rx_fifo_inst_rRamRdAddr_5;
    wire fifo_inst_rx_fifo_inst_rRamRdAddr_4;
    wire fifo_inst_rx_fifo_inst_rRamRdAddr_2;
    wire fifo_inst_rx_fifo_inst_rRamRdAddr_7;
    wire fifo_inst_rx_fifo_inst_rRamRdAddr_6;
    wire \uart_inst0.tx_uart_fifo_inst.m58_eZ0Z_5_cascade_ ;
    wire \uart_inst0.tx_uart_fifo_inst.m58_eZ0Z_6 ;
    wire \uart_inst0.tx_uart_fifo_inst.N_99 ;
    wire rRamRdAddr_RNI0S8U_0;
    wire fifo_inst_rx_fifo_inst_wRamRdEn;
    wire \uart_inst0.tx_uart_fifo_inst.N_99_cascade_ ;
    wire fifo_inst_rx_fifo_inst_rRamRdAddr_0;
    wire rUartRxDataZ0Z_3;
    wire rUartTxDataZ0Z_3;
    wire rUartRxDataZ0Z_4;
    wire rRxDataZ0Z_4;
    wire rUartTxDataZ0Z_4;
    wire rUartRxDataZ0Z_7;
    wire rUartTxDataZ0Z_7;
    wire rUartRxDataZ0Z_2;
    wire rUartTxDataZ0Z_2;
    wire rUartRxDataZ0Z_0;
    wire rUartRxFlagZ0;
    wire rUartTxDataZ0Z_0;
    wire rUartTxEn_4_0;
    wire rUartRxState_0_0;
    wire \uart_inst0.uart_inst0.rx_stateZ0Z_0 ;
    wire \uart_inst0.wRxWrEn_0 ;
    wire \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_0_0 ;
    wire \uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ1Z_1 ;
    wire \uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ0Z_2 ;
    wire \uart_inst0.uart_inst0.rx_stateZ0Z_5 ;
    wire \uart_inst0.uart_inst0.N_283_cascade_ ;
    wire \uart_inst0.uart_inst0.rx_stateZ0Z_6 ;
    wire \uart_inst0.uart_inst0.rx_state_srsts_0_o2_3_3 ;
    wire \uart_inst0.uart_inst0.rx_countdown_2_sqmuxa_i_1 ;
    wire \uart_inst0.uart_inst0.un1_rx_clk_divider_0 ;
    wire \uart_inst0.uart_inst0.N_258_0_cascade_ ;
    wire \uart_inst0.uart_inst0.rx_countdownZ0Z_0 ;
    wire bfn_16_15_0_;
    wire \uart_inst0.uart_inst0.rx_countdownZ0Z_1 ;
    wire \uart_inst0.uart_inst0.rx_countdown_s_1 ;
    wire \uart_inst0.uart_inst0.rx_countdown_cry_0 ;
    wire \uart_inst0.uart_inst0.rx_countdownZ0Z_2 ;
    wire \uart_inst0.uart_inst0.rx_countdown_s_2 ;
    wire \uart_inst0.uart_inst0.rx_countdown_cry_1 ;
    wire \uart_inst0.uart_inst0.rx_countdownZ0Z_3 ;
    wire \uart_inst0.uart_inst0.rx_countdown_s_3 ;
    wire \uart_inst0.uart_inst0.rx_countdown_cry_2 ;
    wire \uart_inst0.uart_inst0.rx_countdownZ0Z_4 ;
    wire \uart_inst0.uart_inst0.rx_countdown_cry_3_THRU_CO ;
    wire \uart_inst0.uart_inst0.rx_countdown_cry_3 ;
    wire \uart_inst0.uart_inst0.N_252_0_i ;
    wire \uart_inst0.uart_inst0.rx_countdown_cry_4 ;
    wire \uart_inst0.uart_inst0.rx_countdownZ0Z_5 ;
    wire \uart_inst0.uart_inst0.rx_countdowne_0_i ;
    wire \uart_inst0.uart_inst0.N_258_0 ;
    wire \uart_inst0.uart_inst0.N_276_cascade_ ;
    wire \uart_inst0.uart_inst0.tx_stateZ0Z_0 ;
    wire \uart_inst0.uart_inst0.tx_stateZ0Z_1 ;
    wire \uart_inst0.uart_inst0.un1_m3_0_a2_0 ;
    wire \uart_inst0.uart_inst0.N_275 ;
    wire \uart_inst0.uart_inst0.N_147_0 ;
    wire bfn_16_18_0_;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_0_s1_THRU_CO ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_0_s1 ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_1_s1_THRU_CO ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_1_s1 ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_2_s1 ;
    wire \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_4 ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_3_s1_THRU_CO ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_3_s1 ;
    wire \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_5 ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_4_s1_THRU_CO ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_4_s1 ;
    wire \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_6 ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_5_s1_THRU_CO ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_5_s1 ;
    wire \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_7 ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_6_s1_THRU_CO ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_6_s1 ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_7_s1 ;
    wire \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_8 ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_7_s1_THRU_CO ;
    wire bfn_16_19_0_;
    wire \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_9 ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_8_s1_THRU_CO ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_8_s1 ;
    wire \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_10 ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_9_s1_THRU_CO ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_9_s1 ;
    wire \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_11 ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_10_s1_THRU_CO ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_10_s1 ;
    wire \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_12 ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_11_s1_THRU_CO ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_11_s1 ;
    wire CONSTANT_ONE_NET;
    wire \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_13 ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_12_s1_THRU_CO ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_12_s1 ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_13_s1 ;
    wire \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_14 ;
    wire \uart_inst0.uart_inst0.N_147_0_i_0 ;
    wire bfn_17_2_0_;
    wire \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_0 ;
    wire \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_1 ;
    wire \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_2 ;
    wire \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_3 ;
    wire \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_4 ;
    wire \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_5 ;
    wire \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_6 ;
    wire \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_7 ;
    wire bfn_17_3_0_;
    wire \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIGAUPZ0 ;
    wire fifo_inst_tx_fifo_inst_rRamRdAddr_2;
    wire fifo_inst_wRxWrFull;
    wire fifo_inst_rx_fifo_inst_rDataCount_2;
    wire fifo_inst_rx_fifo_inst_rDataCount_0;
    wire fifo_inst_rx_fifo_inst_rDataCount_1;
    wire rRxDataZ0Z_6;
    wire rRxDataZ0Z_1;
    wire rRxDataZ0Z_2;
    wire rRxDataZ0Z_3;
    wire rRxDataZ0Z_0;
    wire rRxDataZ0Z_5;
    wire rRxDataZ0Z_7;
    wire N_27_0;
    wire bfn_17_6_0_;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_0 ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_1 ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_2 ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_3 ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_4 ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_5 ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_6 ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_7 ;
    wire bfn_17_7_0_;
    wire \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNO_0_0_3 ;
    wire \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNO_0_0_0 ;
    wire wUartRxEmpty_cascade_;
    wire \uart_inst0.rx_uart_fifo_inst.wRamWrEn ;
    wire \uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_0 ;
    wire \uart_inst0.rx_uart_fifo_inst.rDataCount_RNI3V391Z0Z_2_cascade_ ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rDataCount15_2_0_0_0 ;
    wire \uart_inst0.rx_uart_fifo_inst.wRamRdEn_cascade_ ;
    wire rUartRxStateZ0Z_0;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rDataCount_c2 ;
    wire \uart_inst0.rx_uart_fifo_inst.rDataCount_0_sqmuxa ;
    wire \uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_2 ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rDataCount_axbxc3_1_1 ;
    wire \uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_1 ;
    wire \uart_inst0.wRxWrFull_0 ;
    wire bfn_17_10_0_;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIK0HSZ0 ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_0 ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_1 ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_2 ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_3 ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_4 ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_5 ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_6 ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_7 ;
    wire bfn_17_11_0_;
    wire \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_1 ;
    wire \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_2 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIOAZ0Z54 ;
    wire \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_0 ;
    wire \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_6 ;
    wire \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_5 ;
    wire \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_7 ;
    wire \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_4 ;
    wire \uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_5 ;
    wire \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_8 ;
    wire \uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_4 ;
    wire wUartRxEmpty;
    wire \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_0 ;
    wire \uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_3 ;
    wire P1A1_c;
    wire \uart_inst0.uart_inst0.rx_stateZ0Z_1 ;
    wire wPllLocked_i;
    wire \uart_inst0.uart_inst0.rRxData_0_sqmuxa ;
    wire wPllLocked;
    wire \uart_inst0.uart_inst0.N_257_0 ;
    wire \uart_inst0.uart_inst0.N_273_cascade_ ;
    wire \uart_inst0.uart_inst0.rx_stateZ0Z_3 ;
    wire \uart_inst0.uart_inst0.rx_state_srsts_0_a5_0_0_3 ;
    wire \uart_inst0.uart_inst0.N_274_2 ;
    wire \uart_inst0.uart_inst0.un1_rx_bits_remaining_c3_cascade_ ;
    wire \uart_inst0.uart_inst0.rx_bits_remainingZ0Z_3 ;
    wire \uart_inst0.uart_inst0.tx_countdownZ0Z_3 ;
    wire \uart_inst0.uart_inst0.tx_N_2 ;
    wire \uart_inst0.uart_inst0.tx_countdownZ0Z_2 ;
    wire N_292_g;
    wire \uart_inst0.uart_inst0.N_147_0_i ;
    wire \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_2_s1_THRU_CO ;
    wire \uart_inst0.uart_inst0.un1_rx_state49_i ;
    wire \uart_inst0.uart_inst0.tx_countdownZ0Z_1 ;
    wire \uart_inst0.uart_inst0.tx_countdownZ0Z_0 ;
    wire \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_9 ;
    wire \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_11_3 ;
    wire \uart_inst0.uart_inst0.tx_m5_0_2_cascade_ ;
    wire \uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_11_4 ;
    wire \uart_inst0.uart_inst0.tx_N_11_mux ;
    wire \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_2 ;
    wire \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_0 ;
    wire \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_3 ;
    wire \uart_inst0.uart_inst0.tx_clk_dividerZ0Z_1 ;
    wire \uart_inst0.uart_inst0.tx_m5_0 ;
    wire ioFifoData_in_5;
    wire \fifo_inst.wRxWrData_5 ;
    wire fifo_inst_rx_fifo_inst_rRamWrAddr_5;
    wire fifo_inst_rx_fifo_inst_rRamWrAddr_4;
    wire fifo_inst_rx_fifo_inst_rRamWrAddr_2;
    wire fifo_inst_rx_fifo_inst_rRamWrAddr_7;
    wire fifo_inst_rx_fifo_inst_rRamWrAddr_6;
    wire \uart_inst0.tx_uart_fifo_inst.m54_eZ0Z_5_cascade_ ;
    wire \uart_inst0.tx_uart_fifo_inst.N_91_cascade_ ;
    wire un1_rRamWrAddr_cry_2_c_RNIOTMG;
    wire fifo_inst_rx_fifo_inst_rRamWrAddr_3;
    wire fifo_inst_rx_fifo_inst_rRamWrAddr_1;
    wire fifo_inst_rx_fifo_inst_rRamWrAddr_8;
    wire \uart_inst0.tx_uart_fifo_inst.m54_eZ0Z_6 ;
    wire rRamWrAddr_RNI9D19_0;
    wire \uart_inst0.tx_uart_fifo_inst.N_91 ;
    wire fifo_inst_rx_fifo_inst_wRamWrEn;
    wire fifo_inst_rx_fifo_inst_rRamWrAddr_0;
    wire \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_4 ;
    wire wRxData_4;
    wire \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_3 ;
    wire wRxData_3;
    wire \INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_4C_net ;
    wire \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_7 ;
    wire wRxData_7;
    wire \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_5 ;
    wire wRxData_5;
    wire \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_1 ;
    wire wRxData_1;
    wire \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_2 ;
    wire wRxData_2;
    wire \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_6 ;
    wire wRxData_6;
    wire \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_0 ;
    wire P1A2_c;
    wire wRxData_0;
    wire \INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7C_net ;
    wire N_84_mux_i;
    wire \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_8 ;
    wire \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_3 ;
    wire \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_2 ;
    wire \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_1 ;
    wire \uart_inst0.rx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_0_cascade_ ;
    wire \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_0 ;
    wire \uart_inst0.rx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_6 ;
    wire \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_6 ;
    wire \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_5 ;
    wire \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_7 ;
    wire \uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_4 ;
    wire \uart_inst0.rx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_5 ;
    wire \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_5 ;
    wire wUartRxData_5;
    wire \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_6 ;
    wire wUartRxData_6;
    wire \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_7 ;
    wire rUartRxEnZ0;
    wire wUartRxData_7;
    wire \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_5C_net ;
    wire \uart_inst0.rx_uart_fifo_inst.wUartRxEmpty_i ;
    wire \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_0 ;
    wire wUartRxData_0;
    wire \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_1 ;
    wire wUartRxData_1;
    wire \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_2 ;
    wire wUartRxData_2;
    wire \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_3 ;
    wire wUartRxData_3;
    wire \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_4 ;
    wire wUartRxData_4;
    wire \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIUFMSZ0 ;
    wire \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_5_0 ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIQ9KSZ0 ;
    wire \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_3_0 ;
    wire \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNID4JC2Z0Z_0 ;
    wire \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_8 ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNISCLSZ0 ;
    wire \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_4_0 ;
    wire \uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7 ;
    wire \uart_inst0.rx_uart_fifo_inst.wRamRdEn ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNIO6JSZ0 ;
    wire \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_2_0 ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI0JNSZ0 ;
    wire \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_6_0 ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIM3ISZ0 ;
    wire \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_1_0 ;
    wire \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI2MOSZ0 ;
    wire \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_7_0 ;
    wire \uart_inst0.uart_inst0.un1_rx_bits_remaining_c1 ;
    wire \uart_inst0.uart_inst0.rx_bits_remaining_2_sqmuxa ;
    wire \uart_inst0.uart_inst0.rx_bits_remainingZ0Z_2 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIQDZ0Z64 ;
    wire \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_1 ;
    wire \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNI0NZ0Z94 ;
    wire \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_4 ;
    wire \uart_inst0.wRxWrData_4 ;
    wire \uart_inst0.wRxWrData_1 ;
    wire \uart_inst0.wRxWrData_0 ;
    wire \uart_inst0.wRxWrData_5 ;
    wire \uart_inst0.wRxWrData_7 ;
    wire \uart_inst0.wRxWrData_6 ;
    wire \uart_inst0.wRxWrData_3 ;
    wire \uart_inst0.wRxWrData_2 ;
    wire \uart_inst0.uart_inst0.rRxData_0_sqmuxa_0 ;
    wire \uart_inst0.uart_inst0.rx_stateZ0Z_2 ;
    wire \uart_inst0.uart_inst0.rx_bits_remainingZ0Z_0 ;
    wire \uart_inst0.uart_inst0.N_283 ;
    wire \uart_inst0.uart_inst0.rx_bits_remainingZ0Z_1 ;
    wire \uart_inst0.uart_inst0.rx_state_2_sqmuxa ;
    wire ioFifoData_in_2;
    wire \fifo_inst.wRxWrData_2 ;
    wire ioFifoData_in_1;
    wire \fifo_inst.wRxWrData_1 ;
    wire ioFifoData_in_3;
    wire \fifo_inst.wRxWrData_3 ;
    wire ioFifoData_in_4;
    wire \fifo_inst.wRxWrData_4 ;
    wire ioFifoData_in_0;
    wire \fifo_inst.wRxWrData_0 ;
    wire ioFifoData_in_7;
    wire \fifo_inst.wRxWrData_7 ;
    wire ioFifoData_in_6;
    wire \fifo_inst.ft2232h_inst.rFifoStateZ0Z_1 ;
    wire \fifo_inst.wRxWrData_6 ;
    wire _gnd_net_;
    wire clk_48mhz;
    wire wPllLocked_i_g;

    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical .WRITE_MODE=1;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical .READ_MODE=1;
    SB_RAM40_4K \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_0,\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_7 ,dangling_wire_1,\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_6 ,dangling_wire_2,\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_5 ,dangling_wire_3,\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_4 ,dangling_wire_4,\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_3 ,dangling_wire_5,\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_2 ,dangling_wire_6,\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_1 ,dangling_wire_7,\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_0 }),
            .RADDR({dangling_wire_8,dangling_wire_9,N__15677,N__15719,N__15500,N__15434,N__15479,N__15740,N__15698,N__11093,N__15455}),
            .WADDR({dangling_wire_10,dangling_wire_11,N__15290,N__15083,N__15137,N__15110,N__15053,N__15263,N__15236,N__15209,N__15179}),
            .MASK({dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27}),
            .WDATA({dangling_wire_28,N__16147,dangling_wire_29,N__16118,dangling_wire_30,N__16166,dangling_wire_31,N__16211,dangling_wire_32,N__16100,dangling_wire_33,N__16082,dangling_wire_34,N__16196,dangling_wire_35,N__16178}),
            .RCLKE(),
            .RCLK(N__16965),
            .RE(N__12278),
            .WCLKE(N__13155),
            .WCLK(\INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net ),
            .WE(N__12257));
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical .WRITE_MODE=1;
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical .READ_MODE=1;
    SB_RAM40_4K \fifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_36,\fifo_inst.rx_fifo_inst.ram512x8_inst.mem_7 ,dangling_wire_37,\fifo_inst.rx_fifo_inst.ram512x8_inst.mem_6 ,dangling_wire_38,\fifo_inst.rx_fifo_inst.ram512x8_inst.mem_5 ,dangling_wire_39,\fifo_inst.rx_fifo_inst.ram512x8_inst.mem_4 ,dangling_wire_40,\fifo_inst.rx_fifo_inst.ram512x8_inst.mem_3 ,dangling_wire_41,\fifo_inst.rx_fifo_inst.ram512x8_inst.mem_2 ,dangling_wire_42,\fifo_inst.rx_fifo_inst.ram512x8_inst.mem_1 ,dangling_wire_43,\fifo_inst.rx_fifo_inst.ram512x8_inst.mem_0 }),
            .RADDR({dangling_wire_44,dangling_wire_45,N__9137,N__10802,N__9008,N__9332,N__10733,N__10748,N__9041,N__10781,N__10460}),
            .WADDR({dangling_wire_46,dangling_wire_47,N__14138,N__14255,N__14228,N__14342,N__14315,N__14189,N__14288,N__14165,N__14804}),
            .MASK({dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51,dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63}),
            .WDATA({dangling_wire_64,N__17095,dangling_wire_65,N__17006,dangling_wire_66,N__14360,dangling_wire_67,N__17155,dangling_wire_68,N__17186,dangling_wire_69,N__15835,dangling_wire_70,N__17210,dangling_wire_71,N__17128}),
            .RCLKE(),
            .RCLK(N__16985),
            .RE(N__12313),
            .WCLKE(N__14836),
            .WCLK(\INVfifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net ),
            .WE(N__12256));
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical .WRITE_MODE=1;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical .READ_MODE=1;
    SB_RAM40_4K \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_72,\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_7 ,dangling_wire_73,\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_6 ,dangling_wire_74,\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_5 ,dangling_wire_75,\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_4 ,dangling_wire_76,\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_3 ,dangling_wire_77,\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_2 ,dangling_wire_78,\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_1 ,dangling_wire_79,\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_0 }),
            .RADDR({dangling_wire_80,dangling_wire_81,N__9428,N__9440,N__9452,N__15581,N__9737,N__9365,N__15605,N__13469,N__9551}),
            .WADDR({dangling_wire_82,dangling_wire_83,N__7577,N__8747,N__8696,N__8723,N__8669,N__7352,N__7382,N__7409,N__7445}),
            .MASK({dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99}),
            .WDATA({dangling_wire_100,N__10838,dangling_wire_101,N__9116,dangling_wire_102,N__9104,dangling_wire_103,N__10859,dangling_wire_104,N__10892,dangling_wire_105,N__10817,dangling_wire_106,N__9092,dangling_wire_107,N__11198}),
            .RCLKE(),
            .RCLK(N__16950),
            .RE(N__12267),
            .WCLKE(N__8510),
            .WCLK(\INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net ),
            .WE(N__12316));
    defparam \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical .WRITE_MODE=1;
    defparam \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical .READ_MODE=1;
    SB_RAM40_4K \fifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0_physical  (
            .RDATA({dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,dangling_wire_122,\fifo_inst.tx_fifo_inst.ram512x8_inst.mem_0 }),
            .RADDR({dangling_wire_123,dangling_wire_124,N__8879,N__8927,N__8951,N__8975,N__10313,N__10433,N__12803,N__8900,N__10376}),
            .WADDR({dangling_wire_125,dangling_wire_126,N__7052,N__7082,N__7109,N__7142,N__6850,N__6890,N__6920,N__6947,N__6983}),
            .MASK({dangling_wire_127,dangling_wire_128,dangling_wire_129,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,dangling_wire_140,dangling_wire_141,dangling_wire_142}),
            .WDATA({dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,N__10106}),
            .RCLKE(),
            .RCLK(N__16990),
            .RE(N__12314),
            .WCLKE(N__7928),
            .WCLK(\INVfifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net ),
            .WE(N__12315));
    defparam \top_pll_inst.top_pll_inst_pll .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \top_pll_inst.top_pll_inst_pll .TEST_MODE=1'b0;
    defparam \top_pll_inst.top_pll_inst_pll .SHIFTREG_DIV_MODE=2'b00;
    defparam \top_pll_inst.top_pll_inst_pll .PLLOUT_SELECT="GENCLK";
    defparam \top_pll_inst.top_pll_inst_pll .FILTER_RANGE=3'b001;
    defparam \top_pll_inst.top_pll_inst_pll .FEEDBACK_PATH="SIMPLE";
    defparam \top_pll_inst.top_pll_inst_pll .FDA_RELATIVE=4'b0000;
    defparam \top_pll_inst.top_pll_inst_pll .FDA_FEEDBACK=4'b0000;
    defparam \top_pll_inst.top_pll_inst_pll .ENABLE_ICEGATE=1'b0;
    defparam \top_pll_inst.top_pll_inst_pll .DIVR=4'b0000;
    defparam \top_pll_inst.top_pll_inst_pll .DIVQ=3'b100;
    defparam \top_pll_inst.top_pll_inst_pll .DIVF=7'b0111111;
    defparam \top_pll_inst.top_pll_inst_pll .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    PLL40 \top_pll_inst.top_pll_inst_pll  (
            .PLLOUTGLOBAL(clk_48mhz),
            .SDI(GNDG0),
            .BYPASS(GNDG0),
            .RESETB(N__6461),
            .PLLOUTCORE(),
            .LOCK(\PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO ),
            .SDO(),
            .SCLK(GNDG0),
            .LATCHINPUTVALUE(GNDG0),
            .EXTFEEDBACK(GNDG0),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLIN(N__17429));
    IO_PAD \top_pll_inst.top_pll_inst_iopad  (
            .OE(VCCG0),
            .DIN(),
            .DOUT(N__17429),
            .PACKAGEPIN(iClk));
    IO_PAD P1A8_obuft_iopad (
            .OE(N__17415),
            .DIN(N__17414),
            .DOUT(N__17413),
            .PACKAGEPIN(P1A8));
    defparam P1A8_obuft_preio.NEG_TRIGGER=1'b0;
    defparam P1A8_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO P1A8_obuft_preio (
            .PADOEN(N__17415),
            .PADOUT(N__17414),
            .PADIN(N__17413),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A4_obuf_iopad (
            .OE(N__17406),
            .DIN(N__17405),
            .DOUT(N__17404),
            .PACKAGEPIN(P1A4));
    defparam P1A4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO P1A4_obuf_preio (
            .PADOEN(N__17406),
            .PADOUT(N__17405),
            .PADIN(N__17404),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8014),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD oRx_n_obuf_iopad (
            .OE(N__17397),
            .DIN(N__17396),
            .DOUT(N__17395),
            .PACKAGEPIN(oRx_n));
    defparam oRx_n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam oRx_n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO oRx_n_obuf_preio (
            .PADOEN(N__17397),
            .PADOUT(N__17396),
            .PADIN(N__17395),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6820),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD iRxF_n_ibuf_iopad (
            .OE(N__17388),
            .DIN(N__17387),
            .DOUT(N__17386),
            .PACKAGEPIN(iRxF_n));
    defparam iRxF_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam iRxF_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO iRxF_n_ibuf_preio (
            .PADOEN(N__17388),
            .PADOUT(N__17387),
            .PADIN(N__17386),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(iRxF_n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A7_obuf_iopad (
            .OE(N__17379),
            .DIN(N__17378),
            .DOUT(N__17377),
            .PACKAGEPIN(P1A7));
    defparam P1A7_obuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A7_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO P1A7_obuf_preio (
            .PADOEN(N__17379),
            .PADOUT(N__17378),
            .PADIN(N__17377),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8615),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_7_iopad (
            .OE(N__17370),
            .DIN(N__17369),
            .DOUT(N__17368),
            .PACKAGEPIN(ioFifoData[7]));
    defparam ioFifoData_iobuf_7_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_7_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_7_preio (
            .PADOEN(N__17370),
            .PADOUT(N__17369),
            .PADIN(N__17368),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10088),
            .DIN0(ioFifoData_in_7),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BTN_N_ibuf_iopad (
            .OE(N__17361),
            .DIN(N__17360),
            .DOUT(N__17359),
            .PACKAGEPIN(BTN_N));
    defparam BTN_N_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam BTN_N_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO BTN_N_ibuf_preio (
            .PADOEN(N__17361),
            .PADOUT(N__17360),
            .PADIN(N__17359),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(BTN_N_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_4_iopad (
            .OE(N__17352),
            .DIN(N__17351),
            .DOUT(N__17350),
            .PACKAGEPIN(ioFifoData[4]));
    defparam ioFifoData_iobuf_4_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_4_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_4_preio (
            .PADOEN(N__17352),
            .PADOUT(N__17351),
            .PADIN(N__17350),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10056),
            .DIN0(ioFifoData_in_4),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_1_iopad (
            .OE(N__17343),
            .DIN(N__17342),
            .DOUT(N__17341),
            .PACKAGEPIN(ioFifoData[1]));
    defparam ioFifoData_iobuf_1_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_1_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_1_preio (
            .PADOEN(N__17343),
            .PADOUT(N__17342),
            .PADIN(N__17341),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10055),
            .DIN0(ioFifoData_in_1),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_5_iopad (
            .OE(N__17334),
            .DIN(N__17333),
            .DOUT(N__17332),
            .PACKAGEPIN(ioFifoData[5]));
    defparam ioFifoData_iobuf_5_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_5_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_5_preio (
            .PADOEN(N__17334),
            .PADOUT(N__17333),
            .PADIN(N__17332),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10057),
            .DIN0(ioFifoData_in_5),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD oTx_n_obuf_iopad (
            .OE(N__17325),
            .DIN(N__17324),
            .DOUT(N__17323),
            .PACKAGEPIN(oTx_n));
    defparam oTx_n_obuf_preio.NEG_TRIGGER=1'b0;
    defparam oTx_n_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO oTx_n_obuf_preio (
            .PADOEN(N__17325),
            .PADOUT(N__17324),
            .PADIN(N__17323),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8021),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD iTxE_n_ibuf_iopad (
            .OE(N__17316),
            .DIN(N__17315),
            .DOUT(N__17314),
            .PACKAGEPIN(iTxE_n));
    defparam iTxE_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam iTxE_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO iTxE_n_ibuf_preio (
            .PADOEN(N__17316),
            .PADOUT(N__17315),
            .PADIN(N__17314),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(iTxE_n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A1_ibuf_iopad (
            .OE(N__17307),
            .DIN(N__17306),
            .DOUT(N__17305),
            .PACKAGEPIN(P1A1));
    defparam P1A1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO P1A1_ibuf_preio (
            .PADOEN(N__17307),
            .PADOUT(N__17306),
            .PADIN(N__17305),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(P1A1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_2_iopad (
            .OE(N__17298),
            .DIN(N__17297),
            .DOUT(N__17296),
            .PACKAGEPIN(ioFifoData[2]));
    defparam ioFifoData_iobuf_2_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_2_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_2_preio (
            .PADOEN(N__17298),
            .PADOUT(N__17297),
            .PADIN(N__17296),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10075),
            .DIN0(ioFifoData_in_2),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A9_obuft_iopad (
            .OE(N__17289),
            .DIN(N__17288),
            .DOUT(N__17287),
            .PACKAGEPIN(P1A9));
    defparam P1A9_obuft_preio.NEG_TRIGGER=1'b0;
    defparam P1A9_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO P1A9_obuft_preio (
            .PADOEN(N__17289),
            .PADOUT(N__17288),
            .PADIN(N__17287),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_6_iopad (
            .OE(N__17280),
            .DIN(N__17279),
            .DOUT(N__17278),
            .PACKAGEPIN(ioFifoData[6]));
    defparam ioFifoData_iobuf_6_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_6_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_6_preio (
            .PADOEN(N__17280),
            .PADOUT(N__17279),
            .PADIN(N__17278),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10087),
            .DIN0(ioFifoData_in_6),
            .DOUT0(N__12470),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_3_iopad (
            .OE(N__17271),
            .DIN(N__17270),
            .DOUT(N__17269),
            .PACKAGEPIN(ioFifoData[3]));
    defparam ioFifoData_iobuf_3_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_3_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_3_preio (
            .PADOEN(N__17271),
            .PADOUT(N__17270),
            .PADIN(N__17269),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10068),
            .DIN0(ioFifoData_in_3),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A2_obuf_iopad (
            .OE(N__17262),
            .DIN(N__17261),
            .DOUT(N__17260),
            .PACKAGEPIN(P1A2));
    defparam P1A2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO P1A2_obuf_preio (
            .PADOEN(N__17262),
            .PADOUT(N__17261),
            .PADIN(N__17260),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__15419),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ioFifoData_iobuf_0_iopad (
            .OE(N__17253),
            .DIN(N__17252),
            .DOUT(N__17251),
            .PACKAGEPIN(ioFifoData[0]));
    defparam ioFifoData_iobuf_0_preio.NEG_TRIGGER=1'b0;
    defparam ioFifoData_iobuf_0_preio.PIN_TYPE=6'b101001;
    PRE_IO ioFifoData_iobuf_0_preio (
            .PADOEN(N__17253),
            .PADOUT(N__17252),
            .PADIN(N__17251),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__10064),
            .DIN0(ioFifoData_in_0),
            .DOUT0(N__8846),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD P1A3_obuf_iopad (
            .OE(N__17244),
            .DIN(N__17243),
            .DOUT(N__17242),
            .PACKAGEPIN(P1A3));
    defparam P1A3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam P1A3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO P1A3_obuf_preio (
            .PADOEN(N__17244),
            .PADOUT(N__17243),
            .PADIN(N__17242),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6821),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__4123 (
            .O(N__17225),
            .I(N__17222));
    LocalMux I__4122 (
            .O(N__17222),
            .I(N__17219));
    Span4Mux_h I__4121 (
            .O(N__17219),
            .I(N__17216));
    IoSpan4Mux I__4120 (
            .O(N__17216),
            .I(N__17213));
    Odrv4 I__4119 (
            .O(N__17213),
            .I(ioFifoData_in_1));
    InMux I__4118 (
            .O(N__17210),
            .I(N__17206));
    InMux I__4117 (
            .O(N__17209),
            .I(N__17203));
    LocalMux I__4116 (
            .O(N__17206),
            .I(N__17200));
    LocalMux I__4115 (
            .O(N__17203),
            .I(\fifo_inst.wRxWrData_1 ));
    Odrv4 I__4114 (
            .O(N__17200),
            .I(\fifo_inst.wRxWrData_1 ));
    InMux I__4113 (
            .O(N__17195),
            .I(N__17192));
    LocalMux I__4112 (
            .O(N__17192),
            .I(N__17189));
    Odrv4 I__4111 (
            .O(N__17189),
            .I(ioFifoData_in_3));
    InMux I__4110 (
            .O(N__17186),
            .I(N__17183));
    LocalMux I__4109 (
            .O(N__17183),
            .I(N__17179));
    InMux I__4108 (
            .O(N__17182),
            .I(N__17176));
    Span4Mux_h I__4107 (
            .O(N__17179),
            .I(N__17173));
    LocalMux I__4106 (
            .O(N__17176),
            .I(\fifo_inst.wRxWrData_3 ));
    Odrv4 I__4105 (
            .O(N__17173),
            .I(\fifo_inst.wRxWrData_3 ));
    InMux I__4104 (
            .O(N__17168),
            .I(N__17165));
    LocalMux I__4103 (
            .O(N__17165),
            .I(N__17162));
    IoSpan4Mux I__4102 (
            .O(N__17162),
            .I(N__17159));
    Odrv4 I__4101 (
            .O(N__17159),
            .I(ioFifoData_in_4));
    InMux I__4100 (
            .O(N__17156),
            .I(N__17152));
    InMux I__4099 (
            .O(N__17155),
            .I(N__17149));
    LocalMux I__4098 (
            .O(N__17152),
            .I(\fifo_inst.wRxWrData_4 ));
    LocalMux I__4097 (
            .O(N__17149),
            .I(\fifo_inst.wRxWrData_4 ));
    InMux I__4096 (
            .O(N__17144),
            .I(N__17141));
    LocalMux I__4095 (
            .O(N__17141),
            .I(N__17138));
    Sp12to4 I__4094 (
            .O(N__17138),
            .I(N__17135));
    Span12Mux_h I__4093 (
            .O(N__17135),
            .I(N__17132));
    Odrv12 I__4092 (
            .O(N__17132),
            .I(ioFifoData_in_0));
    InMux I__4091 (
            .O(N__17129),
            .I(N__17125));
    InMux I__4090 (
            .O(N__17128),
            .I(N__17122));
    LocalMux I__4089 (
            .O(N__17125),
            .I(\fifo_inst.wRxWrData_0 ));
    LocalMux I__4088 (
            .O(N__17122),
            .I(\fifo_inst.wRxWrData_0 ));
    InMux I__4087 (
            .O(N__17117),
            .I(N__17114));
    LocalMux I__4086 (
            .O(N__17114),
            .I(N__17111));
    Span4Mux_h I__4085 (
            .O(N__17111),
            .I(N__17108));
    Sp12to4 I__4084 (
            .O(N__17108),
            .I(N__17105));
    Span12Mux_v I__4083 (
            .O(N__17105),
            .I(N__17102));
    Span12Mux_v I__4082 (
            .O(N__17102),
            .I(N__17099));
    Odrv12 I__4081 (
            .O(N__17099),
            .I(ioFifoData_in_7));
    InMux I__4080 (
            .O(N__17096),
            .I(N__17092));
    InMux I__4079 (
            .O(N__17095),
            .I(N__17089));
    LocalMux I__4078 (
            .O(N__17092),
            .I(\fifo_inst.wRxWrData_7 ));
    LocalMux I__4077 (
            .O(N__17089),
            .I(\fifo_inst.wRxWrData_7 ));
    InMux I__4076 (
            .O(N__17084),
            .I(N__17081));
    LocalMux I__4075 (
            .O(N__17081),
            .I(N__17078));
    Span4Mux_v I__4074 (
            .O(N__17078),
            .I(N__17075));
    Sp12to4 I__4073 (
            .O(N__17075),
            .I(N__17072));
    Span12Mux_s6_h I__4072 (
            .O(N__17072),
            .I(N__17069));
    Span12Mux_v I__4071 (
            .O(N__17069),
            .I(N__17066));
    Odrv12 I__4070 (
            .O(N__17066),
            .I(ioFifoData_in_6));
    InMux I__4069 (
            .O(N__17063),
            .I(N__17044));
    InMux I__4068 (
            .O(N__17062),
            .I(N__17044));
    InMux I__4067 (
            .O(N__17061),
            .I(N__17044));
    InMux I__4066 (
            .O(N__17060),
            .I(N__17044));
    InMux I__4065 (
            .O(N__17059),
            .I(N__17044));
    InMux I__4064 (
            .O(N__17058),
            .I(N__17044));
    InMux I__4063 (
            .O(N__17057),
            .I(N__17041));
    LocalMux I__4062 (
            .O(N__17044),
            .I(N__17035));
    LocalMux I__4061 (
            .O(N__17041),
            .I(N__17035));
    InMux I__4060 (
            .O(N__17040),
            .I(N__17032));
    Span4Mux_v I__4059 (
            .O(N__17035),
            .I(N__17029));
    LocalMux I__4058 (
            .O(N__17032),
            .I(N__17022));
    Sp12to4 I__4057 (
            .O(N__17029),
            .I(N__17022));
    InMux I__4056 (
            .O(N__17028),
            .I(N__17019));
    InMux I__4055 (
            .O(N__17027),
            .I(N__17016));
    Span12Mux_s11_h I__4054 (
            .O(N__17022),
            .I(N__17011));
    LocalMux I__4053 (
            .O(N__17019),
            .I(N__17011));
    LocalMux I__4052 (
            .O(N__17016),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_1 ));
    Odrv12 I__4051 (
            .O(N__17011),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_1 ));
    InMux I__4050 (
            .O(N__17006),
            .I(N__17002));
    InMux I__4049 (
            .O(N__17005),
            .I(N__16999));
    LocalMux I__4048 (
            .O(N__17002),
            .I(N__16996));
    LocalMux I__4047 (
            .O(N__16999),
            .I(\fifo_inst.wRxWrData_6 ));
    Odrv4 I__4046 (
            .O(N__16996),
            .I(\fifo_inst.wRxWrData_6 ));
    ClkMux I__4045 (
            .O(N__16991),
            .I(N__16706));
    ClkMux I__4044 (
            .O(N__16990),
            .I(N__16706));
    ClkMux I__4043 (
            .O(N__16989),
            .I(N__16706));
    ClkMux I__4042 (
            .O(N__16988),
            .I(N__16706));
    ClkMux I__4041 (
            .O(N__16987),
            .I(N__16706));
    ClkMux I__4040 (
            .O(N__16986),
            .I(N__16706));
    ClkMux I__4039 (
            .O(N__16985),
            .I(N__16706));
    ClkMux I__4038 (
            .O(N__16984),
            .I(N__16706));
    ClkMux I__4037 (
            .O(N__16983),
            .I(N__16706));
    ClkMux I__4036 (
            .O(N__16982),
            .I(N__16706));
    ClkMux I__4035 (
            .O(N__16981),
            .I(N__16706));
    ClkMux I__4034 (
            .O(N__16980),
            .I(N__16706));
    ClkMux I__4033 (
            .O(N__16979),
            .I(N__16706));
    ClkMux I__4032 (
            .O(N__16978),
            .I(N__16706));
    ClkMux I__4031 (
            .O(N__16977),
            .I(N__16706));
    ClkMux I__4030 (
            .O(N__16976),
            .I(N__16706));
    ClkMux I__4029 (
            .O(N__16975),
            .I(N__16706));
    ClkMux I__4028 (
            .O(N__16974),
            .I(N__16706));
    ClkMux I__4027 (
            .O(N__16973),
            .I(N__16706));
    ClkMux I__4026 (
            .O(N__16972),
            .I(N__16706));
    ClkMux I__4025 (
            .O(N__16971),
            .I(N__16706));
    ClkMux I__4024 (
            .O(N__16970),
            .I(N__16706));
    ClkMux I__4023 (
            .O(N__16969),
            .I(N__16706));
    ClkMux I__4022 (
            .O(N__16968),
            .I(N__16706));
    ClkMux I__4021 (
            .O(N__16967),
            .I(N__16706));
    ClkMux I__4020 (
            .O(N__16966),
            .I(N__16706));
    ClkMux I__4019 (
            .O(N__16965),
            .I(N__16706));
    ClkMux I__4018 (
            .O(N__16964),
            .I(N__16706));
    ClkMux I__4017 (
            .O(N__16963),
            .I(N__16706));
    ClkMux I__4016 (
            .O(N__16962),
            .I(N__16706));
    ClkMux I__4015 (
            .O(N__16961),
            .I(N__16706));
    ClkMux I__4014 (
            .O(N__16960),
            .I(N__16706));
    ClkMux I__4013 (
            .O(N__16959),
            .I(N__16706));
    ClkMux I__4012 (
            .O(N__16958),
            .I(N__16706));
    ClkMux I__4011 (
            .O(N__16957),
            .I(N__16706));
    ClkMux I__4010 (
            .O(N__16956),
            .I(N__16706));
    ClkMux I__4009 (
            .O(N__16955),
            .I(N__16706));
    ClkMux I__4008 (
            .O(N__16954),
            .I(N__16706));
    ClkMux I__4007 (
            .O(N__16953),
            .I(N__16706));
    ClkMux I__4006 (
            .O(N__16952),
            .I(N__16706));
    ClkMux I__4005 (
            .O(N__16951),
            .I(N__16706));
    ClkMux I__4004 (
            .O(N__16950),
            .I(N__16706));
    ClkMux I__4003 (
            .O(N__16949),
            .I(N__16706));
    ClkMux I__4002 (
            .O(N__16948),
            .I(N__16706));
    ClkMux I__4001 (
            .O(N__16947),
            .I(N__16706));
    ClkMux I__4000 (
            .O(N__16946),
            .I(N__16706));
    ClkMux I__3999 (
            .O(N__16945),
            .I(N__16706));
    ClkMux I__3998 (
            .O(N__16944),
            .I(N__16706));
    ClkMux I__3997 (
            .O(N__16943),
            .I(N__16706));
    ClkMux I__3996 (
            .O(N__16942),
            .I(N__16706));
    ClkMux I__3995 (
            .O(N__16941),
            .I(N__16706));
    ClkMux I__3994 (
            .O(N__16940),
            .I(N__16706));
    ClkMux I__3993 (
            .O(N__16939),
            .I(N__16706));
    ClkMux I__3992 (
            .O(N__16938),
            .I(N__16706));
    ClkMux I__3991 (
            .O(N__16937),
            .I(N__16706));
    ClkMux I__3990 (
            .O(N__16936),
            .I(N__16706));
    ClkMux I__3989 (
            .O(N__16935),
            .I(N__16706));
    ClkMux I__3988 (
            .O(N__16934),
            .I(N__16706));
    ClkMux I__3987 (
            .O(N__16933),
            .I(N__16706));
    ClkMux I__3986 (
            .O(N__16932),
            .I(N__16706));
    ClkMux I__3985 (
            .O(N__16931),
            .I(N__16706));
    ClkMux I__3984 (
            .O(N__16930),
            .I(N__16706));
    ClkMux I__3983 (
            .O(N__16929),
            .I(N__16706));
    ClkMux I__3982 (
            .O(N__16928),
            .I(N__16706));
    ClkMux I__3981 (
            .O(N__16927),
            .I(N__16706));
    ClkMux I__3980 (
            .O(N__16926),
            .I(N__16706));
    ClkMux I__3979 (
            .O(N__16925),
            .I(N__16706));
    ClkMux I__3978 (
            .O(N__16924),
            .I(N__16706));
    ClkMux I__3977 (
            .O(N__16923),
            .I(N__16706));
    ClkMux I__3976 (
            .O(N__16922),
            .I(N__16706));
    ClkMux I__3975 (
            .O(N__16921),
            .I(N__16706));
    ClkMux I__3974 (
            .O(N__16920),
            .I(N__16706));
    ClkMux I__3973 (
            .O(N__16919),
            .I(N__16706));
    ClkMux I__3972 (
            .O(N__16918),
            .I(N__16706));
    ClkMux I__3971 (
            .O(N__16917),
            .I(N__16706));
    ClkMux I__3970 (
            .O(N__16916),
            .I(N__16706));
    ClkMux I__3969 (
            .O(N__16915),
            .I(N__16706));
    ClkMux I__3968 (
            .O(N__16914),
            .I(N__16706));
    ClkMux I__3967 (
            .O(N__16913),
            .I(N__16706));
    ClkMux I__3966 (
            .O(N__16912),
            .I(N__16706));
    ClkMux I__3965 (
            .O(N__16911),
            .I(N__16706));
    ClkMux I__3964 (
            .O(N__16910),
            .I(N__16706));
    ClkMux I__3963 (
            .O(N__16909),
            .I(N__16706));
    ClkMux I__3962 (
            .O(N__16908),
            .I(N__16706));
    ClkMux I__3961 (
            .O(N__16907),
            .I(N__16706));
    ClkMux I__3960 (
            .O(N__16906),
            .I(N__16706));
    ClkMux I__3959 (
            .O(N__16905),
            .I(N__16706));
    ClkMux I__3958 (
            .O(N__16904),
            .I(N__16706));
    ClkMux I__3957 (
            .O(N__16903),
            .I(N__16706));
    ClkMux I__3956 (
            .O(N__16902),
            .I(N__16706));
    ClkMux I__3955 (
            .O(N__16901),
            .I(N__16706));
    ClkMux I__3954 (
            .O(N__16900),
            .I(N__16706));
    ClkMux I__3953 (
            .O(N__16899),
            .I(N__16706));
    ClkMux I__3952 (
            .O(N__16898),
            .I(N__16706));
    ClkMux I__3951 (
            .O(N__16897),
            .I(N__16706));
    GlobalMux I__3950 (
            .O(N__16706),
            .I(clk_48mhz));
    CascadeMux I__3949 (
            .O(N__16703),
            .I(N__16690));
    CascadeMux I__3948 (
            .O(N__16702),
            .I(N__16671));
    CascadeMux I__3947 (
            .O(N__16701),
            .I(N__16667));
    CascadeMux I__3946 (
            .O(N__16700),
            .I(N__16654));
    CascadeMux I__3945 (
            .O(N__16699),
            .I(N__16650));
    CascadeMux I__3944 (
            .O(N__16698),
            .I(N__16646));
    CascadeMux I__3943 (
            .O(N__16697),
            .I(N__16641));
    InMux I__3942 (
            .O(N__16696),
            .I(N__16615));
    InMux I__3941 (
            .O(N__16695),
            .I(N__16610));
    InMux I__3940 (
            .O(N__16694),
            .I(N__16610));
    InMux I__3939 (
            .O(N__16693),
            .I(N__16607));
    InMux I__3938 (
            .O(N__16690),
            .I(N__16594));
    InMux I__3937 (
            .O(N__16689),
            .I(N__16594));
    InMux I__3936 (
            .O(N__16688),
            .I(N__16594));
    InMux I__3935 (
            .O(N__16687),
            .I(N__16594));
    InMux I__3934 (
            .O(N__16686),
            .I(N__16594));
    InMux I__3933 (
            .O(N__16685),
            .I(N__16594));
    InMux I__3932 (
            .O(N__16684),
            .I(N__16589));
    InMux I__3931 (
            .O(N__16683),
            .I(N__16589));
    InMux I__3930 (
            .O(N__16682),
            .I(N__16580));
    InMux I__3929 (
            .O(N__16681),
            .I(N__16580));
    InMux I__3928 (
            .O(N__16680),
            .I(N__16580));
    InMux I__3927 (
            .O(N__16679),
            .I(N__16580));
    InMux I__3926 (
            .O(N__16678),
            .I(N__16577));
    InMux I__3925 (
            .O(N__16677),
            .I(N__16572));
    InMux I__3924 (
            .O(N__16676),
            .I(N__16572));
    InMux I__3923 (
            .O(N__16675),
            .I(N__16569));
    InMux I__3922 (
            .O(N__16674),
            .I(N__16566));
    InMux I__3921 (
            .O(N__16671),
            .I(N__16563));
    InMux I__3920 (
            .O(N__16670),
            .I(N__16560));
    InMux I__3919 (
            .O(N__16667),
            .I(N__16555));
    InMux I__3918 (
            .O(N__16666),
            .I(N__16555));
    InMux I__3917 (
            .O(N__16665),
            .I(N__16548));
    InMux I__3916 (
            .O(N__16664),
            .I(N__16548));
    InMux I__3915 (
            .O(N__16663),
            .I(N__16548));
    InMux I__3914 (
            .O(N__16662),
            .I(N__16541));
    InMux I__3913 (
            .O(N__16661),
            .I(N__16541));
    InMux I__3912 (
            .O(N__16660),
            .I(N__16541));
    InMux I__3911 (
            .O(N__16659),
            .I(N__16538));
    InMux I__3910 (
            .O(N__16658),
            .I(N__16531));
    InMux I__3909 (
            .O(N__16657),
            .I(N__16531));
    InMux I__3908 (
            .O(N__16654),
            .I(N__16531));
    InMux I__3907 (
            .O(N__16653),
            .I(N__16526));
    InMux I__3906 (
            .O(N__16650),
            .I(N__16526));
    InMux I__3905 (
            .O(N__16649),
            .I(N__16523));
    InMux I__3904 (
            .O(N__16646),
            .I(N__16518));
    InMux I__3903 (
            .O(N__16645),
            .I(N__16518));
    InMux I__3902 (
            .O(N__16644),
            .I(N__16511));
    InMux I__3901 (
            .O(N__16641),
            .I(N__16511));
    InMux I__3900 (
            .O(N__16640),
            .I(N__16511));
    InMux I__3899 (
            .O(N__16639),
            .I(N__16504));
    InMux I__3898 (
            .O(N__16638),
            .I(N__16504));
    InMux I__3897 (
            .O(N__16637),
            .I(N__16504));
    InMux I__3896 (
            .O(N__16636),
            .I(N__16497));
    InMux I__3895 (
            .O(N__16635),
            .I(N__16497));
    InMux I__3894 (
            .O(N__16634),
            .I(N__16497));
    InMux I__3893 (
            .O(N__16633),
            .I(N__16490));
    InMux I__3892 (
            .O(N__16632),
            .I(N__16490));
    InMux I__3891 (
            .O(N__16631),
            .I(N__16490));
    InMux I__3890 (
            .O(N__16630),
            .I(N__16483));
    InMux I__3889 (
            .O(N__16629),
            .I(N__16483));
    InMux I__3888 (
            .O(N__16628),
            .I(N__16483));
    InMux I__3887 (
            .O(N__16627),
            .I(N__16480));
    InMux I__3886 (
            .O(N__16626),
            .I(N__16473));
    InMux I__3885 (
            .O(N__16625),
            .I(N__16473));
    InMux I__3884 (
            .O(N__16624),
            .I(N__16473));
    InMux I__3883 (
            .O(N__16623),
            .I(N__16466));
    InMux I__3882 (
            .O(N__16622),
            .I(N__16466));
    InMux I__3881 (
            .O(N__16621),
            .I(N__16466));
    InMux I__3880 (
            .O(N__16620),
            .I(N__16459));
    InMux I__3879 (
            .O(N__16619),
            .I(N__16459));
    InMux I__3878 (
            .O(N__16618),
            .I(N__16459));
    LocalMux I__3877 (
            .O(N__16615),
            .I(N__16456));
    LocalMux I__3876 (
            .O(N__16610),
            .I(N__16450));
    LocalMux I__3875 (
            .O(N__16607),
            .I(N__16445));
    LocalMux I__3874 (
            .O(N__16594),
            .I(N__16442));
    LocalMux I__3873 (
            .O(N__16589),
            .I(N__16439));
    LocalMux I__3872 (
            .O(N__16580),
            .I(N__16433));
    LocalMux I__3871 (
            .O(N__16577),
            .I(N__16430));
    LocalMux I__3870 (
            .O(N__16572),
            .I(N__16426));
    LocalMux I__3869 (
            .O(N__16569),
            .I(N__16422));
    LocalMux I__3868 (
            .O(N__16566),
            .I(N__16410));
    LocalMux I__3867 (
            .O(N__16563),
            .I(N__16407));
    LocalMux I__3866 (
            .O(N__16560),
            .I(N__16404));
    LocalMux I__3865 (
            .O(N__16555),
            .I(N__16401));
    LocalMux I__3864 (
            .O(N__16548),
            .I(N__16398));
    LocalMux I__3863 (
            .O(N__16541),
            .I(N__16395));
    LocalMux I__3862 (
            .O(N__16538),
            .I(N__16392));
    LocalMux I__3861 (
            .O(N__16531),
            .I(N__16389));
    LocalMux I__3860 (
            .O(N__16526),
            .I(N__16386));
    LocalMux I__3859 (
            .O(N__16523),
            .I(N__16381));
    LocalMux I__3858 (
            .O(N__16518),
            .I(N__16378));
    LocalMux I__3857 (
            .O(N__16511),
            .I(N__16375));
    LocalMux I__3856 (
            .O(N__16504),
            .I(N__16372));
    LocalMux I__3855 (
            .O(N__16497),
            .I(N__16369));
    LocalMux I__3854 (
            .O(N__16490),
            .I(N__16363));
    LocalMux I__3853 (
            .O(N__16483),
            .I(N__16360));
    LocalMux I__3852 (
            .O(N__16480),
            .I(N__16352));
    LocalMux I__3851 (
            .O(N__16473),
            .I(N__16347));
    LocalMux I__3850 (
            .O(N__16466),
            .I(N__16344));
    LocalMux I__3849 (
            .O(N__16459),
            .I(N__16341));
    Glb2LocalMux I__3848 (
            .O(N__16456),
            .I(N__16217));
    SRMux I__3847 (
            .O(N__16455),
            .I(N__16217));
    SRMux I__3846 (
            .O(N__16454),
            .I(N__16217));
    SRMux I__3845 (
            .O(N__16453),
            .I(N__16217));
    Glb2LocalMux I__3844 (
            .O(N__16450),
            .I(N__16217));
    SRMux I__3843 (
            .O(N__16449),
            .I(N__16217));
    SRMux I__3842 (
            .O(N__16448),
            .I(N__16217));
    Glb2LocalMux I__3841 (
            .O(N__16445),
            .I(N__16217));
    Glb2LocalMux I__3840 (
            .O(N__16442),
            .I(N__16217));
    Glb2LocalMux I__3839 (
            .O(N__16439),
            .I(N__16217));
    SRMux I__3838 (
            .O(N__16438),
            .I(N__16217));
    SRMux I__3837 (
            .O(N__16437),
            .I(N__16217));
    SRMux I__3836 (
            .O(N__16436),
            .I(N__16217));
    Glb2LocalMux I__3835 (
            .O(N__16433),
            .I(N__16217));
    Glb2LocalMux I__3834 (
            .O(N__16430),
            .I(N__16217));
    SRMux I__3833 (
            .O(N__16429),
            .I(N__16217));
    Glb2LocalMux I__3832 (
            .O(N__16426),
            .I(N__16217));
    SRMux I__3831 (
            .O(N__16425),
            .I(N__16217));
    Glb2LocalMux I__3830 (
            .O(N__16422),
            .I(N__16217));
    SRMux I__3829 (
            .O(N__16421),
            .I(N__16217));
    SRMux I__3828 (
            .O(N__16420),
            .I(N__16217));
    SRMux I__3827 (
            .O(N__16419),
            .I(N__16217));
    SRMux I__3826 (
            .O(N__16418),
            .I(N__16217));
    SRMux I__3825 (
            .O(N__16417),
            .I(N__16217));
    SRMux I__3824 (
            .O(N__16416),
            .I(N__16217));
    SRMux I__3823 (
            .O(N__16415),
            .I(N__16217));
    SRMux I__3822 (
            .O(N__16414),
            .I(N__16217));
    SRMux I__3821 (
            .O(N__16413),
            .I(N__16217));
    Glb2LocalMux I__3820 (
            .O(N__16410),
            .I(N__16217));
    Glb2LocalMux I__3819 (
            .O(N__16407),
            .I(N__16217));
    Glb2LocalMux I__3818 (
            .O(N__16404),
            .I(N__16217));
    Glb2LocalMux I__3817 (
            .O(N__16401),
            .I(N__16217));
    Glb2LocalMux I__3816 (
            .O(N__16398),
            .I(N__16217));
    Glb2LocalMux I__3815 (
            .O(N__16395),
            .I(N__16217));
    Glb2LocalMux I__3814 (
            .O(N__16392),
            .I(N__16217));
    Glb2LocalMux I__3813 (
            .O(N__16389),
            .I(N__16217));
    Glb2LocalMux I__3812 (
            .O(N__16386),
            .I(N__16217));
    SRMux I__3811 (
            .O(N__16385),
            .I(N__16217));
    SRMux I__3810 (
            .O(N__16384),
            .I(N__16217));
    Glb2LocalMux I__3809 (
            .O(N__16381),
            .I(N__16217));
    Glb2LocalMux I__3808 (
            .O(N__16378),
            .I(N__16217));
    Glb2LocalMux I__3807 (
            .O(N__16375),
            .I(N__16217));
    Glb2LocalMux I__3806 (
            .O(N__16372),
            .I(N__16217));
    Glb2LocalMux I__3805 (
            .O(N__16369),
            .I(N__16217));
    SRMux I__3804 (
            .O(N__16368),
            .I(N__16217));
    SRMux I__3803 (
            .O(N__16367),
            .I(N__16217));
    SRMux I__3802 (
            .O(N__16366),
            .I(N__16217));
    Glb2LocalMux I__3801 (
            .O(N__16363),
            .I(N__16217));
    Glb2LocalMux I__3800 (
            .O(N__16360),
            .I(N__16217));
    SRMux I__3799 (
            .O(N__16359),
            .I(N__16217));
    SRMux I__3798 (
            .O(N__16358),
            .I(N__16217));
    SRMux I__3797 (
            .O(N__16357),
            .I(N__16217));
    SRMux I__3796 (
            .O(N__16356),
            .I(N__16217));
    SRMux I__3795 (
            .O(N__16355),
            .I(N__16217));
    Glb2LocalMux I__3794 (
            .O(N__16352),
            .I(N__16217));
    SRMux I__3793 (
            .O(N__16351),
            .I(N__16217));
    SRMux I__3792 (
            .O(N__16350),
            .I(N__16217));
    Glb2LocalMux I__3791 (
            .O(N__16347),
            .I(N__16217));
    Glb2LocalMux I__3790 (
            .O(N__16344),
            .I(N__16217));
    Glb2LocalMux I__3789 (
            .O(N__16341),
            .I(N__16217));
    SRMux I__3788 (
            .O(N__16340),
            .I(N__16217));
    GlobalMux I__3787 (
            .O(N__16217),
            .I(N__16214));
    gio2CtrlBuf I__3786 (
            .O(N__16214),
            .I(wPllLocked_i_g));
    InMux I__3785 (
            .O(N__16211),
            .I(N__16207));
    InMux I__3784 (
            .O(N__16210),
            .I(N__16204));
    LocalMux I__3783 (
            .O(N__16207),
            .I(N__16201));
    LocalMux I__3782 (
            .O(N__16204),
            .I(\uart_inst0.wRxWrData_4 ));
    Odrv4 I__3781 (
            .O(N__16201),
            .I(\uart_inst0.wRxWrData_4 ));
    InMux I__3780 (
            .O(N__16196),
            .I(N__16193));
    LocalMux I__3779 (
            .O(N__16193),
            .I(N__16189));
    InMux I__3778 (
            .O(N__16192),
            .I(N__16186));
    Span4Mux_h I__3777 (
            .O(N__16189),
            .I(N__16183));
    LocalMux I__3776 (
            .O(N__16186),
            .I(\uart_inst0.wRxWrData_1 ));
    Odrv4 I__3775 (
            .O(N__16183),
            .I(\uart_inst0.wRxWrData_1 ));
    InMux I__3774 (
            .O(N__16178),
            .I(N__16175));
    LocalMux I__3773 (
            .O(N__16175),
            .I(N__16172));
    Span4Mux_h I__3772 (
            .O(N__16172),
            .I(N__16169));
    Odrv4 I__3771 (
            .O(N__16169),
            .I(\uart_inst0.wRxWrData_0 ));
    InMux I__3770 (
            .O(N__16166),
            .I(N__16163));
    LocalMux I__3769 (
            .O(N__16163),
            .I(N__16159));
    InMux I__3768 (
            .O(N__16162),
            .I(N__16156));
    Span4Mux_v I__3767 (
            .O(N__16159),
            .I(N__16153));
    LocalMux I__3766 (
            .O(N__16156),
            .I(\uart_inst0.wRxWrData_5 ));
    Odrv4 I__3765 (
            .O(N__16153),
            .I(\uart_inst0.wRxWrData_5 ));
    InMux I__3764 (
            .O(N__16148),
            .I(N__16144));
    InMux I__3763 (
            .O(N__16147),
            .I(N__16141));
    LocalMux I__3762 (
            .O(N__16144),
            .I(N__16138));
    LocalMux I__3761 (
            .O(N__16141),
            .I(N__16134));
    Span4Mux_v I__3760 (
            .O(N__16138),
            .I(N__16131));
    InMux I__3759 (
            .O(N__16137),
            .I(N__16128));
    Span4Mux_h I__3758 (
            .O(N__16134),
            .I(N__16125));
    Odrv4 I__3757 (
            .O(N__16131),
            .I(\uart_inst0.wRxWrData_7 ));
    LocalMux I__3756 (
            .O(N__16128),
            .I(\uart_inst0.wRxWrData_7 ));
    Odrv4 I__3755 (
            .O(N__16125),
            .I(\uart_inst0.wRxWrData_7 ));
    InMux I__3754 (
            .O(N__16118),
            .I(N__16115));
    LocalMux I__3753 (
            .O(N__16115),
            .I(N__16111));
    InMux I__3752 (
            .O(N__16114),
            .I(N__16108));
    Span4Mux_h I__3751 (
            .O(N__16111),
            .I(N__16105));
    LocalMux I__3750 (
            .O(N__16108),
            .I(\uart_inst0.wRxWrData_6 ));
    Odrv4 I__3749 (
            .O(N__16105),
            .I(\uart_inst0.wRxWrData_6 ));
    InMux I__3748 (
            .O(N__16100),
            .I(N__16097));
    LocalMux I__3747 (
            .O(N__16097),
            .I(N__16093));
    InMux I__3746 (
            .O(N__16096),
            .I(N__16090));
    Span4Mux_v I__3745 (
            .O(N__16093),
            .I(N__16087));
    LocalMux I__3744 (
            .O(N__16090),
            .I(\uart_inst0.wRxWrData_3 ));
    Odrv4 I__3743 (
            .O(N__16087),
            .I(\uart_inst0.wRxWrData_3 ));
    InMux I__3742 (
            .O(N__16082),
            .I(N__16078));
    InMux I__3741 (
            .O(N__16081),
            .I(N__16075));
    LocalMux I__3740 (
            .O(N__16078),
            .I(N__16072));
    LocalMux I__3739 (
            .O(N__16075),
            .I(\uart_inst0.wRxWrData_2 ));
    Odrv4 I__3738 (
            .O(N__16072),
            .I(\uart_inst0.wRxWrData_2 ));
    CEMux I__3737 (
            .O(N__16067),
            .I(N__16063));
    CEMux I__3736 (
            .O(N__16066),
            .I(N__16060));
    LocalMux I__3735 (
            .O(N__16063),
            .I(N__16057));
    LocalMux I__3734 (
            .O(N__16060),
            .I(N__16054));
    Odrv4 I__3733 (
            .O(N__16057),
            .I(\uart_inst0.uart_inst0.rRxData_0_sqmuxa_0 ));
    Odrv4 I__3732 (
            .O(N__16054),
            .I(\uart_inst0.uart_inst0.rRxData_0_sqmuxa_0 ));
    InMux I__3731 (
            .O(N__16049),
            .I(N__16045));
    InMux I__3730 (
            .O(N__16048),
            .I(N__16041));
    LocalMux I__3729 (
            .O(N__16045),
            .I(N__16038));
    CascadeMux I__3728 (
            .O(N__16044),
            .I(N__16029));
    LocalMux I__3727 (
            .O(N__16041),
            .I(N__16026));
    Span4Mux_h I__3726 (
            .O(N__16038),
            .I(N__16023));
    InMux I__3725 (
            .O(N__16037),
            .I(N__16019));
    InMux I__3724 (
            .O(N__16036),
            .I(N__16014));
    InMux I__3723 (
            .O(N__16035),
            .I(N__16014));
    InMux I__3722 (
            .O(N__16034),
            .I(N__16009));
    InMux I__3721 (
            .O(N__16033),
            .I(N__16009));
    InMux I__3720 (
            .O(N__16032),
            .I(N__16004));
    InMux I__3719 (
            .O(N__16029),
            .I(N__16004));
    Span4Mux_v I__3718 (
            .O(N__16026),
            .I(N__16001));
    Span4Mux_v I__3717 (
            .O(N__16023),
            .I(N__15998));
    InMux I__3716 (
            .O(N__16022),
            .I(N__15995));
    LocalMux I__3715 (
            .O(N__16019),
            .I(N__15990));
    LocalMux I__3714 (
            .O(N__16014),
            .I(N__15990));
    LocalMux I__3713 (
            .O(N__16009),
            .I(N__15985));
    LocalMux I__3712 (
            .O(N__16004),
            .I(N__15985));
    Odrv4 I__3711 (
            .O(N__16001),
            .I(\uart_inst0.uart_inst0.rx_stateZ0Z_2 ));
    Odrv4 I__3710 (
            .O(N__15998),
            .I(\uart_inst0.uart_inst0.rx_stateZ0Z_2 ));
    LocalMux I__3709 (
            .O(N__15995),
            .I(\uart_inst0.uart_inst0.rx_stateZ0Z_2 ));
    Odrv4 I__3708 (
            .O(N__15990),
            .I(\uart_inst0.uart_inst0.rx_stateZ0Z_2 ));
    Odrv4 I__3707 (
            .O(N__15985),
            .I(\uart_inst0.uart_inst0.rx_stateZ0Z_2 ));
    CascadeMux I__3706 (
            .O(N__15974),
            .I(N__15970));
    CascadeMux I__3705 (
            .O(N__15973),
            .I(N__15966));
    InMux I__3704 (
            .O(N__15970),
            .I(N__15961));
    InMux I__3703 (
            .O(N__15969),
            .I(N__15958));
    InMux I__3702 (
            .O(N__15966),
            .I(N__15953));
    InMux I__3701 (
            .O(N__15965),
            .I(N__15953));
    InMux I__3700 (
            .O(N__15964),
            .I(N__15950));
    LocalMux I__3699 (
            .O(N__15961),
            .I(N__15943));
    LocalMux I__3698 (
            .O(N__15958),
            .I(N__15943));
    LocalMux I__3697 (
            .O(N__15953),
            .I(N__15943));
    LocalMux I__3696 (
            .O(N__15950),
            .I(\uart_inst0.uart_inst0.rx_bits_remainingZ0Z_0 ));
    Odrv4 I__3695 (
            .O(N__15943),
            .I(\uart_inst0.uart_inst0.rx_bits_remainingZ0Z_0 ));
    InMux I__3694 (
            .O(N__15938),
            .I(N__15934));
    InMux I__3693 (
            .O(N__15937),
            .I(N__15930));
    LocalMux I__3692 (
            .O(N__15934),
            .I(N__15927));
    InMux I__3691 (
            .O(N__15933),
            .I(N__15924));
    LocalMux I__3690 (
            .O(N__15930),
            .I(N__15913));
    Span4Mux_v I__3689 (
            .O(N__15927),
            .I(N__15913));
    LocalMux I__3688 (
            .O(N__15924),
            .I(N__15913));
    InMux I__3687 (
            .O(N__15923),
            .I(N__15910));
    InMux I__3686 (
            .O(N__15922),
            .I(N__15903));
    InMux I__3685 (
            .O(N__15921),
            .I(N__15903));
    InMux I__3684 (
            .O(N__15920),
            .I(N__15903));
    Odrv4 I__3683 (
            .O(N__15913),
            .I(\uart_inst0.uart_inst0.N_283 ));
    LocalMux I__3682 (
            .O(N__15910),
            .I(\uart_inst0.uart_inst0.N_283 ));
    LocalMux I__3681 (
            .O(N__15903),
            .I(\uart_inst0.uart_inst0.N_283 ));
    InMux I__3680 (
            .O(N__15896),
            .I(N__15892));
    InMux I__3679 (
            .O(N__15895),
            .I(N__15888));
    LocalMux I__3678 (
            .O(N__15892),
            .I(N__15885));
    InMux I__3677 (
            .O(N__15891),
            .I(N__15882));
    LocalMux I__3676 (
            .O(N__15888),
            .I(\uart_inst0.uart_inst0.rx_bits_remainingZ0Z_1 ));
    Odrv12 I__3675 (
            .O(N__15885),
            .I(\uart_inst0.uart_inst0.rx_bits_remainingZ0Z_1 ));
    LocalMux I__3674 (
            .O(N__15882),
            .I(\uart_inst0.uart_inst0.rx_bits_remainingZ0Z_1 ));
    SRMux I__3673 (
            .O(N__15875),
            .I(N__15871));
    SRMux I__3672 (
            .O(N__15874),
            .I(N__15868));
    LocalMux I__3671 (
            .O(N__15871),
            .I(N__15865));
    LocalMux I__3670 (
            .O(N__15868),
            .I(N__15861));
    Span4Mux_h I__3669 (
            .O(N__15865),
            .I(N__15858));
    InMux I__3668 (
            .O(N__15864),
            .I(N__15855));
    Odrv4 I__3667 (
            .O(N__15861),
            .I(\uart_inst0.uart_inst0.rx_state_2_sqmuxa ));
    Odrv4 I__3666 (
            .O(N__15858),
            .I(\uart_inst0.uart_inst0.rx_state_2_sqmuxa ));
    LocalMux I__3665 (
            .O(N__15855),
            .I(\uart_inst0.uart_inst0.rx_state_2_sqmuxa ));
    InMux I__3664 (
            .O(N__15848),
            .I(N__15845));
    LocalMux I__3663 (
            .O(N__15845),
            .I(N__15842));
    Span4Mux_h I__3662 (
            .O(N__15842),
            .I(N__15839));
    Odrv4 I__3661 (
            .O(N__15839),
            .I(ioFifoData_in_2));
    InMux I__3660 (
            .O(N__15836),
            .I(N__15832));
    InMux I__3659 (
            .O(N__15835),
            .I(N__15829));
    LocalMux I__3658 (
            .O(N__15832),
            .I(\fifo_inst.wRxWrData_2 ));
    LocalMux I__3657 (
            .O(N__15829),
            .I(\fifo_inst.wRxWrData_2 ));
    InMux I__3656 (
            .O(N__15824),
            .I(N__15818));
    InMux I__3655 (
            .O(N__15823),
            .I(N__15815));
    InMux I__3654 (
            .O(N__15822),
            .I(N__15812));
    InMux I__3653 (
            .O(N__15821),
            .I(N__15809));
    LocalMux I__3652 (
            .O(N__15818),
            .I(\uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7 ));
    LocalMux I__3651 (
            .O(N__15815),
            .I(\uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7 ));
    LocalMux I__3650 (
            .O(N__15812),
            .I(\uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7 ));
    LocalMux I__3649 (
            .O(N__15809),
            .I(\uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7 ));
    InMux I__3648 (
            .O(N__15800),
            .I(N__15795));
    CascadeMux I__3647 (
            .O(N__15799),
            .I(N__15791));
    CascadeMux I__3646 (
            .O(N__15798),
            .I(N__15786));
    LocalMux I__3645 (
            .O(N__15795),
            .I(N__15783));
    InMux I__3644 (
            .O(N__15794),
            .I(N__15780));
    InMux I__3643 (
            .O(N__15791),
            .I(N__15777));
    InMux I__3642 (
            .O(N__15790),
            .I(N__15774));
    CEMux I__3641 (
            .O(N__15789),
            .I(N__15771));
    InMux I__3640 (
            .O(N__15786),
            .I(N__15768));
    Odrv4 I__3639 (
            .O(N__15783),
            .I(\uart_inst0.rx_uart_fifo_inst.wRamRdEn ));
    LocalMux I__3638 (
            .O(N__15780),
            .I(\uart_inst0.rx_uart_fifo_inst.wRamRdEn ));
    LocalMux I__3637 (
            .O(N__15777),
            .I(\uart_inst0.rx_uart_fifo_inst.wRamRdEn ));
    LocalMux I__3636 (
            .O(N__15774),
            .I(\uart_inst0.rx_uart_fifo_inst.wRamRdEn ));
    LocalMux I__3635 (
            .O(N__15771),
            .I(\uart_inst0.rx_uart_fifo_inst.wRamRdEn ));
    LocalMux I__3634 (
            .O(N__15768),
            .I(\uart_inst0.rx_uart_fifo_inst.wRamRdEn ));
    InMux I__3633 (
            .O(N__15755),
            .I(N__15752));
    LocalMux I__3632 (
            .O(N__15752),
            .I(N__15748));
    InMux I__3631 (
            .O(N__15751),
            .I(N__15745));
    Odrv4 I__3630 (
            .O(N__15748),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNIO6JSZ0 ));
    LocalMux I__3629 (
            .O(N__15745),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNIO6JSZ0 ));
    CascadeMux I__3628 (
            .O(N__15740),
            .I(N__15737));
    InMux I__3627 (
            .O(N__15737),
            .I(N__15734));
    LocalMux I__3626 (
            .O(N__15734),
            .I(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_2_0 ));
    InMux I__3625 (
            .O(N__15731),
            .I(N__15727));
    InMux I__3624 (
            .O(N__15730),
            .I(N__15724));
    LocalMux I__3623 (
            .O(N__15727),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI0JNSZ0 ));
    LocalMux I__3622 (
            .O(N__15724),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI0JNSZ0 ));
    CascadeMux I__3621 (
            .O(N__15719),
            .I(N__15716));
    InMux I__3620 (
            .O(N__15716),
            .I(N__15713));
    LocalMux I__3619 (
            .O(N__15713),
            .I(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_6_0 ));
    InMux I__3618 (
            .O(N__15710),
            .I(N__15706));
    InMux I__3617 (
            .O(N__15709),
            .I(N__15703));
    LocalMux I__3616 (
            .O(N__15706),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIM3ISZ0 ));
    LocalMux I__3615 (
            .O(N__15703),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIM3ISZ0 ));
    CascadeMux I__3614 (
            .O(N__15698),
            .I(N__15695));
    InMux I__3613 (
            .O(N__15695),
            .I(N__15692));
    LocalMux I__3612 (
            .O(N__15692),
            .I(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_1_0 ));
    InMux I__3611 (
            .O(N__15689),
            .I(N__15685));
    InMux I__3610 (
            .O(N__15688),
            .I(N__15682));
    LocalMux I__3609 (
            .O(N__15685),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI2MOSZ0 ));
    LocalMux I__3608 (
            .O(N__15682),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI2MOSZ0 ));
    CascadeMux I__3607 (
            .O(N__15677),
            .I(N__15674));
    InMux I__3606 (
            .O(N__15674),
            .I(N__15671));
    LocalMux I__3605 (
            .O(N__15671),
            .I(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_7_0 ));
    InMux I__3604 (
            .O(N__15668),
            .I(N__15665));
    LocalMux I__3603 (
            .O(N__15665),
            .I(N__15662));
    Odrv4 I__3602 (
            .O(N__15662),
            .I(\uart_inst0.uart_inst0.un1_rx_bits_remaining_c1 ));
    InMux I__3601 (
            .O(N__15659),
            .I(N__15656));
    LocalMux I__3600 (
            .O(N__15656),
            .I(N__15651));
    InMux I__3599 (
            .O(N__15655),
            .I(N__15646));
    InMux I__3598 (
            .O(N__15654),
            .I(N__15646));
    Odrv4 I__3597 (
            .O(N__15651),
            .I(\uart_inst0.uart_inst0.rx_bits_remaining_2_sqmuxa ));
    LocalMux I__3596 (
            .O(N__15646),
            .I(\uart_inst0.uart_inst0.rx_bits_remaining_2_sqmuxa ));
    CascadeMux I__3595 (
            .O(N__15641),
            .I(N__15638));
    InMux I__3594 (
            .O(N__15638),
            .I(N__15634));
    InMux I__3593 (
            .O(N__15637),
            .I(N__15631));
    LocalMux I__3592 (
            .O(N__15634),
            .I(N__15626));
    LocalMux I__3591 (
            .O(N__15631),
            .I(N__15626));
    Odrv4 I__3590 (
            .O(N__15626),
            .I(\uart_inst0.uart_inst0.rx_bits_remainingZ0Z_2 ));
    InMux I__3589 (
            .O(N__15623),
            .I(N__15619));
    InMux I__3588 (
            .O(N__15622),
            .I(N__15616));
    LocalMux I__3587 (
            .O(N__15619),
            .I(N__15613));
    LocalMux I__3586 (
            .O(N__15616),
            .I(N__15610));
    Odrv4 I__3585 (
            .O(N__15613),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIQDZ0Z64 ));
    Odrv12 I__3584 (
            .O(N__15610),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIQDZ0Z64 ));
    CascadeMux I__3583 (
            .O(N__15605),
            .I(N__15602));
    InMux I__3582 (
            .O(N__15602),
            .I(N__15599));
    LocalMux I__3581 (
            .O(N__15599),
            .I(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_1 ));
    InMux I__3580 (
            .O(N__15596),
            .I(N__15592));
    InMux I__3579 (
            .O(N__15595),
            .I(N__15589));
    LocalMux I__3578 (
            .O(N__15592),
            .I(N__15586));
    LocalMux I__3577 (
            .O(N__15589),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNI0NZ0Z94 ));
    Odrv12 I__3576 (
            .O(N__15586),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNI0NZ0Z94 ));
    CascadeMux I__3575 (
            .O(N__15581),
            .I(N__15578));
    InMux I__3574 (
            .O(N__15578),
            .I(N__15575));
    LocalMux I__3573 (
            .O(N__15575),
            .I(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_4 ));
    InMux I__3572 (
            .O(N__15572),
            .I(N__15569));
    LocalMux I__3571 (
            .O(N__15569),
            .I(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_1 ));
    InMux I__3570 (
            .O(N__15566),
            .I(N__15563));
    LocalMux I__3569 (
            .O(N__15563),
            .I(N__15560));
    Odrv12 I__3568 (
            .O(N__15560),
            .I(wUartRxData_1));
    InMux I__3567 (
            .O(N__15557),
            .I(N__15554));
    LocalMux I__3566 (
            .O(N__15554),
            .I(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_2 ));
    InMux I__3565 (
            .O(N__15551),
            .I(N__15548));
    LocalMux I__3564 (
            .O(N__15548),
            .I(N__15545));
    Odrv4 I__3563 (
            .O(N__15545),
            .I(wUartRxData_2));
    InMux I__3562 (
            .O(N__15542),
            .I(N__15539));
    LocalMux I__3561 (
            .O(N__15539),
            .I(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_3 ));
    InMux I__3560 (
            .O(N__15536),
            .I(N__15533));
    LocalMux I__3559 (
            .O(N__15533),
            .I(N__15530));
    Odrv12 I__3558 (
            .O(N__15530),
            .I(wUartRxData_3));
    InMux I__3557 (
            .O(N__15527),
            .I(N__15524));
    LocalMux I__3556 (
            .O(N__15524),
            .I(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_4 ));
    InMux I__3555 (
            .O(N__15521),
            .I(N__15518));
    LocalMux I__3554 (
            .O(N__15518),
            .I(N__15515));
    Odrv4 I__3553 (
            .O(N__15515),
            .I(wUartRxData_4));
    InMux I__3552 (
            .O(N__15512),
            .I(N__15508));
    InMux I__3551 (
            .O(N__15511),
            .I(N__15505));
    LocalMux I__3550 (
            .O(N__15508),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIUFMSZ0 ));
    LocalMux I__3549 (
            .O(N__15505),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIUFMSZ0 ));
    CascadeMux I__3548 (
            .O(N__15500),
            .I(N__15497));
    InMux I__3547 (
            .O(N__15497),
            .I(N__15494));
    LocalMux I__3546 (
            .O(N__15494),
            .I(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_5_0 ));
    InMux I__3545 (
            .O(N__15491),
            .I(N__15487));
    InMux I__3544 (
            .O(N__15490),
            .I(N__15484));
    LocalMux I__3543 (
            .O(N__15487),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIQ9KSZ0 ));
    LocalMux I__3542 (
            .O(N__15484),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIQ9KSZ0 ));
    CascadeMux I__3541 (
            .O(N__15479),
            .I(N__15476));
    InMux I__3540 (
            .O(N__15476),
            .I(N__15473));
    LocalMux I__3539 (
            .O(N__15473),
            .I(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_3_0 ));
    InMux I__3538 (
            .O(N__15470),
            .I(N__15467));
    LocalMux I__3537 (
            .O(N__15467),
            .I(N__15463));
    InMux I__3536 (
            .O(N__15466),
            .I(N__15460));
    Odrv4 I__3535 (
            .O(N__15463),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNID4JC2Z0Z_0 ));
    LocalMux I__3534 (
            .O(N__15460),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNID4JC2Z0Z_0 ));
    CascadeMux I__3533 (
            .O(N__15455),
            .I(N__15452));
    InMux I__3532 (
            .O(N__15452),
            .I(N__15449));
    LocalMux I__3531 (
            .O(N__15449),
            .I(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_8 ));
    InMux I__3530 (
            .O(N__15446),
            .I(N__15442));
    InMux I__3529 (
            .O(N__15445),
            .I(N__15439));
    LocalMux I__3528 (
            .O(N__15442),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNISCLSZ0 ));
    LocalMux I__3527 (
            .O(N__15439),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNISCLSZ0 ));
    CascadeMux I__3526 (
            .O(N__15434),
            .I(N__15431));
    InMux I__3525 (
            .O(N__15431),
            .I(N__15428));
    LocalMux I__3524 (
            .O(N__15428),
            .I(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_4_0 ));
    InMux I__3523 (
            .O(N__15425),
            .I(N__15422));
    LocalMux I__3522 (
            .O(N__15422),
            .I(\fifo_inst.rx_fifo_inst.ram512x8_inst.mem_0 ));
    IoInMux I__3521 (
            .O(N__15419),
            .I(N__15416));
    LocalMux I__3520 (
            .O(N__15416),
            .I(N__15413));
    IoSpan4Mux I__3519 (
            .O(N__15413),
            .I(N__15408));
    InMux I__3518 (
            .O(N__15412),
            .I(N__15403));
    InMux I__3517 (
            .O(N__15411),
            .I(N__15403));
    Span4Mux_s3_v I__3516 (
            .O(N__15408),
            .I(N__15394));
    LocalMux I__3515 (
            .O(N__15403),
            .I(N__15391));
    InMux I__3514 (
            .O(N__15402),
            .I(N__15378));
    InMux I__3513 (
            .O(N__15401),
            .I(N__15378));
    InMux I__3512 (
            .O(N__15400),
            .I(N__15378));
    InMux I__3511 (
            .O(N__15399),
            .I(N__15378));
    InMux I__3510 (
            .O(N__15398),
            .I(N__15378));
    InMux I__3509 (
            .O(N__15397),
            .I(N__15378));
    Span4Mux_h I__3508 (
            .O(N__15394),
            .I(N__15369));
    Span4Mux_s3_v I__3507 (
            .O(N__15391),
            .I(N__15369));
    LocalMux I__3506 (
            .O(N__15378),
            .I(N__15369));
    CascadeMux I__3505 (
            .O(N__15377),
            .I(N__15358));
    InMux I__3504 (
            .O(N__15376),
            .I(N__15355));
    Span4Mux_h I__3503 (
            .O(N__15369),
            .I(N__15352));
    InMux I__3502 (
            .O(N__15368),
            .I(N__15349));
    InMux I__3501 (
            .O(N__15367),
            .I(N__15338));
    InMux I__3500 (
            .O(N__15366),
            .I(N__15338));
    InMux I__3499 (
            .O(N__15365),
            .I(N__15338));
    InMux I__3498 (
            .O(N__15364),
            .I(N__15338));
    InMux I__3497 (
            .O(N__15363),
            .I(N__15338));
    InMux I__3496 (
            .O(N__15362),
            .I(N__15331));
    InMux I__3495 (
            .O(N__15361),
            .I(N__15331));
    InMux I__3494 (
            .O(N__15358),
            .I(N__15331));
    LocalMux I__3493 (
            .O(N__15355),
            .I(P1A2_c));
    Odrv4 I__3492 (
            .O(N__15352),
            .I(P1A2_c));
    LocalMux I__3491 (
            .O(N__15349),
            .I(P1A2_c));
    LocalMux I__3490 (
            .O(N__15338),
            .I(P1A2_c));
    LocalMux I__3489 (
            .O(N__15331),
            .I(P1A2_c));
    InMux I__3488 (
            .O(N__15320),
            .I(N__15316));
    InMux I__3487 (
            .O(N__15319),
            .I(N__15313));
    LocalMux I__3486 (
            .O(N__15316),
            .I(wRxData_0));
    LocalMux I__3485 (
            .O(N__15313),
            .I(wRxData_0));
    CEMux I__3484 (
            .O(N__15308),
            .I(N__15305));
    LocalMux I__3483 (
            .O(N__15305),
            .I(N__15301));
    CEMux I__3482 (
            .O(N__15304),
            .I(N__15298));
    Span4Mux_s2_v I__3481 (
            .O(N__15301),
            .I(N__15293));
    LocalMux I__3480 (
            .O(N__15298),
            .I(N__15293));
    Odrv4 I__3479 (
            .O(N__15293),
            .I(N_84_mux_i));
    CascadeMux I__3478 (
            .O(N__15290),
            .I(N__15287));
    InMux I__3477 (
            .O(N__15287),
            .I(N__15283));
    InMux I__3476 (
            .O(N__15286),
            .I(N__15280));
    LocalMux I__3475 (
            .O(N__15283),
            .I(N__15277));
    LocalMux I__3474 (
            .O(N__15280),
            .I(N__15271));
    Span4Mux_v I__3473 (
            .O(N__15277),
            .I(N__15271));
    InMux I__3472 (
            .O(N__15276),
            .I(N__15268));
    Odrv4 I__3471 (
            .O(N__15271),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_8 ));
    LocalMux I__3470 (
            .O(N__15268),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_8 ));
    CascadeMux I__3469 (
            .O(N__15263),
            .I(N__15260));
    InMux I__3468 (
            .O(N__15260),
            .I(N__15257));
    LocalMux I__3467 (
            .O(N__15257),
            .I(N__15254));
    Span4Mux_h I__3466 (
            .O(N__15254),
            .I(N__15249));
    InMux I__3465 (
            .O(N__15253),
            .I(N__15246));
    InMux I__3464 (
            .O(N__15252),
            .I(N__15243));
    Odrv4 I__3463 (
            .O(N__15249),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_3 ));
    LocalMux I__3462 (
            .O(N__15246),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_3 ));
    LocalMux I__3461 (
            .O(N__15243),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_3 ));
    CascadeMux I__3460 (
            .O(N__15236),
            .I(N__15233));
    InMux I__3459 (
            .O(N__15233),
            .I(N__15230));
    LocalMux I__3458 (
            .O(N__15230),
            .I(N__15226));
    InMux I__3457 (
            .O(N__15229),
            .I(N__15222));
    Span4Mux_v I__3456 (
            .O(N__15226),
            .I(N__15219));
    InMux I__3455 (
            .O(N__15225),
            .I(N__15216));
    LocalMux I__3454 (
            .O(N__15222),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_2 ));
    Odrv4 I__3453 (
            .O(N__15219),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_2 ));
    LocalMux I__3452 (
            .O(N__15216),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_2 ));
    CascadeMux I__3451 (
            .O(N__15209),
            .I(N__15206));
    InMux I__3450 (
            .O(N__15206),
            .I(N__15203));
    LocalMux I__3449 (
            .O(N__15203),
            .I(N__15199));
    InMux I__3448 (
            .O(N__15202),
            .I(N__15195));
    Span4Mux_v I__3447 (
            .O(N__15199),
            .I(N__15192));
    InMux I__3446 (
            .O(N__15198),
            .I(N__15189));
    LocalMux I__3445 (
            .O(N__15195),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_1 ));
    Odrv4 I__3444 (
            .O(N__15192),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_1 ));
    LocalMux I__3443 (
            .O(N__15189),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_1 ));
    CascadeMux I__3442 (
            .O(N__15182),
            .I(\uart_inst0.rx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_0_cascade_ ));
    CascadeMux I__3441 (
            .O(N__15179),
            .I(N__15176));
    InMux I__3440 (
            .O(N__15176),
            .I(N__15173));
    LocalMux I__3439 (
            .O(N__15173),
            .I(N__15169));
    InMux I__3438 (
            .O(N__15172),
            .I(N__15165));
    Span4Mux_h I__3437 (
            .O(N__15169),
            .I(N__15162));
    InMux I__3436 (
            .O(N__15168),
            .I(N__15159));
    LocalMux I__3435 (
            .O(N__15165),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_0 ));
    Odrv4 I__3434 (
            .O(N__15162),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_0 ));
    LocalMux I__3433 (
            .O(N__15159),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_0 ));
    CascadeMux I__3432 (
            .O(N__15152),
            .I(N__15149));
    InMux I__3431 (
            .O(N__15149),
            .I(N__15145));
    InMux I__3430 (
            .O(N__15148),
            .I(N__15142));
    LocalMux I__3429 (
            .O(N__15145),
            .I(\uart_inst0.rx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_6 ));
    LocalMux I__3428 (
            .O(N__15142),
            .I(\uart_inst0.rx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_6 ));
    CascadeMux I__3427 (
            .O(N__15137),
            .I(N__15134));
    InMux I__3426 (
            .O(N__15134),
            .I(N__15131));
    LocalMux I__3425 (
            .O(N__15131),
            .I(N__15128));
    Span4Mux_v I__3424 (
            .O(N__15128),
            .I(N__15123));
    InMux I__3423 (
            .O(N__15127),
            .I(N__15120));
    InMux I__3422 (
            .O(N__15126),
            .I(N__15117));
    Odrv4 I__3421 (
            .O(N__15123),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_6 ));
    LocalMux I__3420 (
            .O(N__15120),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_6 ));
    LocalMux I__3419 (
            .O(N__15117),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_6 ));
    CascadeMux I__3418 (
            .O(N__15110),
            .I(N__15107));
    InMux I__3417 (
            .O(N__15107),
            .I(N__15104));
    LocalMux I__3416 (
            .O(N__15104),
            .I(N__15101));
    Span4Mux_v I__3415 (
            .O(N__15101),
            .I(N__15096));
    InMux I__3414 (
            .O(N__15100),
            .I(N__15093));
    InMux I__3413 (
            .O(N__15099),
            .I(N__15090));
    Odrv4 I__3412 (
            .O(N__15096),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_5 ));
    LocalMux I__3411 (
            .O(N__15093),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_5 ));
    LocalMux I__3410 (
            .O(N__15090),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_5 ));
    CascadeMux I__3409 (
            .O(N__15083),
            .I(N__15080));
    InMux I__3408 (
            .O(N__15080),
            .I(N__15076));
    CascadeMux I__3407 (
            .O(N__15079),
            .I(N__15073));
    LocalMux I__3406 (
            .O(N__15076),
            .I(N__15069));
    InMux I__3405 (
            .O(N__15073),
            .I(N__15066));
    InMux I__3404 (
            .O(N__15072),
            .I(N__15063));
    Span4Mux_v I__3403 (
            .O(N__15069),
            .I(N__15060));
    LocalMux I__3402 (
            .O(N__15066),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_7 ));
    LocalMux I__3401 (
            .O(N__15063),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_7 ));
    Odrv4 I__3400 (
            .O(N__15060),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_7 ));
    CascadeMux I__3399 (
            .O(N__15053),
            .I(N__15050));
    InMux I__3398 (
            .O(N__15050),
            .I(N__15047));
    LocalMux I__3397 (
            .O(N__15047),
            .I(N__15044));
    Span4Mux_v I__3396 (
            .O(N__15044),
            .I(N__15039));
    InMux I__3395 (
            .O(N__15043),
            .I(N__15036));
    InMux I__3394 (
            .O(N__15042),
            .I(N__15033));
    Odrv4 I__3393 (
            .O(N__15039),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_4 ));
    LocalMux I__3392 (
            .O(N__15036),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_4 ));
    LocalMux I__3391 (
            .O(N__15033),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_4 ));
    CascadeMux I__3390 (
            .O(N__15026),
            .I(N__15022));
    InMux I__3389 (
            .O(N__15025),
            .I(N__15017));
    InMux I__3388 (
            .O(N__15022),
            .I(N__15017));
    LocalMux I__3387 (
            .O(N__15017),
            .I(\uart_inst0.rx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_5 ));
    InMux I__3386 (
            .O(N__15014),
            .I(N__15011));
    LocalMux I__3385 (
            .O(N__15011),
            .I(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_5 ));
    InMux I__3384 (
            .O(N__15008),
            .I(N__15004));
    InMux I__3383 (
            .O(N__15007),
            .I(N__15001));
    LocalMux I__3382 (
            .O(N__15004),
            .I(N__14998));
    LocalMux I__3381 (
            .O(N__15001),
            .I(wUartRxData_5));
    Odrv12 I__3380 (
            .O(N__14998),
            .I(wUartRxData_5));
    CascadeMux I__3379 (
            .O(N__14993),
            .I(N__14990));
    InMux I__3378 (
            .O(N__14990),
            .I(N__14987));
    LocalMux I__3377 (
            .O(N__14987),
            .I(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_6 ));
    InMux I__3376 (
            .O(N__14984),
            .I(N__14980));
    InMux I__3375 (
            .O(N__14983),
            .I(N__14977));
    LocalMux I__3374 (
            .O(N__14980),
            .I(N__14974));
    LocalMux I__3373 (
            .O(N__14977),
            .I(wUartRxData_6));
    Odrv12 I__3372 (
            .O(N__14974),
            .I(wUartRxData_6));
    InMux I__3371 (
            .O(N__14969),
            .I(N__14966));
    LocalMux I__3370 (
            .O(N__14966),
            .I(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_7 ));
    InMux I__3369 (
            .O(N__14963),
            .I(N__14957));
    CascadeMux I__3368 (
            .O(N__14962),
            .I(N__14954));
    CascadeMux I__3367 (
            .O(N__14961),
            .I(N__14951));
    InMux I__3366 (
            .O(N__14960),
            .I(N__14940));
    LocalMux I__3365 (
            .O(N__14957),
            .I(N__14937));
    InMux I__3364 (
            .O(N__14954),
            .I(N__14934));
    InMux I__3363 (
            .O(N__14951),
            .I(N__14931));
    InMux I__3362 (
            .O(N__14950),
            .I(N__14928));
    InMux I__3361 (
            .O(N__14949),
            .I(N__14925));
    InMux I__3360 (
            .O(N__14948),
            .I(N__14918));
    InMux I__3359 (
            .O(N__14947),
            .I(N__14918));
    InMux I__3358 (
            .O(N__14946),
            .I(N__14918));
    InMux I__3357 (
            .O(N__14945),
            .I(N__14911));
    InMux I__3356 (
            .O(N__14944),
            .I(N__14911));
    InMux I__3355 (
            .O(N__14943),
            .I(N__14911));
    LocalMux I__3354 (
            .O(N__14940),
            .I(rUartRxEnZ0));
    Odrv4 I__3353 (
            .O(N__14937),
            .I(rUartRxEnZ0));
    LocalMux I__3352 (
            .O(N__14934),
            .I(rUartRxEnZ0));
    LocalMux I__3351 (
            .O(N__14931),
            .I(rUartRxEnZ0));
    LocalMux I__3350 (
            .O(N__14928),
            .I(rUartRxEnZ0));
    LocalMux I__3349 (
            .O(N__14925),
            .I(rUartRxEnZ0));
    LocalMux I__3348 (
            .O(N__14918),
            .I(rUartRxEnZ0));
    LocalMux I__3347 (
            .O(N__14911),
            .I(rUartRxEnZ0));
    InMux I__3346 (
            .O(N__14894),
            .I(N__14890));
    InMux I__3345 (
            .O(N__14893),
            .I(N__14887));
    LocalMux I__3344 (
            .O(N__14890),
            .I(N__14884));
    LocalMux I__3343 (
            .O(N__14887),
            .I(wUartRxData_7));
    Odrv4 I__3342 (
            .O(N__14884),
            .I(wUartRxData_7));
    CEMux I__3341 (
            .O(N__14879),
            .I(N__14876));
    LocalMux I__3340 (
            .O(N__14876),
            .I(N__14873));
    Odrv4 I__3339 (
            .O(N__14873),
            .I(\uart_inst0.rx_uart_fifo_inst.wUartRxEmpty_i ));
    InMux I__3338 (
            .O(N__14870),
            .I(N__14867));
    LocalMux I__3337 (
            .O(N__14867),
            .I(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_0 ));
    InMux I__3336 (
            .O(N__14864),
            .I(N__14861));
    LocalMux I__3335 (
            .O(N__14861),
            .I(N__14858));
    Odrv12 I__3334 (
            .O(N__14858),
            .I(wUartRxData_0));
    InMux I__3333 (
            .O(N__14855),
            .I(N__14852));
    LocalMux I__3332 (
            .O(N__14852),
            .I(rRamWrAddr_RNI9D19_0));
    InMux I__3331 (
            .O(N__14849),
            .I(N__14846));
    LocalMux I__3330 (
            .O(N__14846),
            .I(\uart_inst0.tx_uart_fifo_inst.N_91 ));
    CascadeMux I__3329 (
            .O(N__14843),
            .I(N__14837));
    InMux I__3328 (
            .O(N__14842),
            .I(N__14831));
    InMux I__3327 (
            .O(N__14841),
            .I(N__14831));
    InMux I__3326 (
            .O(N__14840),
            .I(N__14828));
    InMux I__3325 (
            .O(N__14837),
            .I(N__14825));
    CEMux I__3324 (
            .O(N__14836),
            .I(N__14822));
    LocalMux I__3323 (
            .O(N__14831),
            .I(N__14815));
    LocalMux I__3322 (
            .O(N__14828),
            .I(N__14815));
    LocalMux I__3321 (
            .O(N__14825),
            .I(N__14815));
    LocalMux I__3320 (
            .O(N__14822),
            .I(N__14812));
    Span4Mux_s3_v I__3319 (
            .O(N__14815),
            .I(N__14807));
    Span4Mux_h I__3318 (
            .O(N__14812),
            .I(N__14807));
    Odrv4 I__3317 (
            .O(N__14807),
            .I(fifo_inst_rx_fifo_inst_wRamWrEn));
    CascadeMux I__3316 (
            .O(N__14804),
            .I(N__14801));
    InMux I__3315 (
            .O(N__14801),
            .I(N__14798));
    LocalMux I__3314 (
            .O(N__14798),
            .I(N__14793));
    InMux I__3313 (
            .O(N__14797),
            .I(N__14790));
    InMux I__3312 (
            .O(N__14796),
            .I(N__14787));
    Odrv4 I__3311 (
            .O(N__14793),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_0));
    LocalMux I__3310 (
            .O(N__14790),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_0));
    LocalMux I__3309 (
            .O(N__14787),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_0));
    InMux I__3308 (
            .O(N__14780),
            .I(N__14777));
    LocalMux I__3307 (
            .O(N__14777),
            .I(\fifo_inst.rx_fifo_inst.ram512x8_inst.mem_4 ));
    InMux I__3306 (
            .O(N__14774),
            .I(N__14771));
    LocalMux I__3305 (
            .O(N__14771),
            .I(N__14767));
    InMux I__3304 (
            .O(N__14770),
            .I(N__14764));
    Span4Mux_v I__3303 (
            .O(N__14767),
            .I(N__14761));
    LocalMux I__3302 (
            .O(N__14764),
            .I(wRxData_4));
    Odrv4 I__3301 (
            .O(N__14761),
            .I(wRxData_4));
    InMux I__3300 (
            .O(N__14756),
            .I(N__14753));
    LocalMux I__3299 (
            .O(N__14753),
            .I(\fifo_inst.rx_fifo_inst.ram512x8_inst.mem_3 ));
    InMux I__3298 (
            .O(N__14750),
            .I(N__14746));
    InMux I__3297 (
            .O(N__14749),
            .I(N__14743));
    LocalMux I__3296 (
            .O(N__14746),
            .I(N__14740));
    LocalMux I__3295 (
            .O(N__14743),
            .I(wRxData_3));
    Odrv4 I__3294 (
            .O(N__14740),
            .I(wRxData_3));
    InMux I__3293 (
            .O(N__14735),
            .I(N__14732));
    LocalMux I__3292 (
            .O(N__14732),
            .I(\fifo_inst.rx_fifo_inst.ram512x8_inst.mem_7 ));
    InMux I__3291 (
            .O(N__14729),
            .I(N__14725));
    InMux I__3290 (
            .O(N__14728),
            .I(N__14722));
    LocalMux I__3289 (
            .O(N__14725),
            .I(wRxData_7));
    LocalMux I__3288 (
            .O(N__14722),
            .I(wRxData_7));
    InMux I__3287 (
            .O(N__14717),
            .I(N__14714));
    LocalMux I__3286 (
            .O(N__14714),
            .I(\fifo_inst.rx_fifo_inst.ram512x8_inst.mem_5 ));
    InMux I__3285 (
            .O(N__14711),
            .I(N__14707));
    InMux I__3284 (
            .O(N__14710),
            .I(N__14704));
    LocalMux I__3283 (
            .O(N__14707),
            .I(wRxData_5));
    LocalMux I__3282 (
            .O(N__14704),
            .I(wRxData_5));
    InMux I__3281 (
            .O(N__14699),
            .I(N__14696));
    LocalMux I__3280 (
            .O(N__14696),
            .I(\fifo_inst.rx_fifo_inst.ram512x8_inst.mem_1 ));
    InMux I__3279 (
            .O(N__14693),
            .I(N__14690));
    LocalMux I__3278 (
            .O(N__14690),
            .I(N__14686));
    InMux I__3277 (
            .O(N__14689),
            .I(N__14683));
    Odrv4 I__3276 (
            .O(N__14686),
            .I(wRxData_1));
    LocalMux I__3275 (
            .O(N__14683),
            .I(wRxData_1));
    InMux I__3274 (
            .O(N__14678),
            .I(N__14675));
    LocalMux I__3273 (
            .O(N__14675),
            .I(\fifo_inst.rx_fifo_inst.ram512x8_inst.mem_2 ));
    InMux I__3272 (
            .O(N__14672),
            .I(N__14668));
    InMux I__3271 (
            .O(N__14671),
            .I(N__14665));
    LocalMux I__3270 (
            .O(N__14668),
            .I(wRxData_2));
    LocalMux I__3269 (
            .O(N__14665),
            .I(wRxData_2));
    InMux I__3268 (
            .O(N__14660),
            .I(N__14657));
    LocalMux I__3267 (
            .O(N__14657),
            .I(\fifo_inst.rx_fifo_inst.ram512x8_inst.mem_6 ));
    InMux I__3266 (
            .O(N__14654),
            .I(N__14650));
    InMux I__3265 (
            .O(N__14653),
            .I(N__14647));
    LocalMux I__3264 (
            .O(N__14650),
            .I(wRxData_6));
    LocalMux I__3263 (
            .O(N__14647),
            .I(wRxData_6));
    SRMux I__3262 (
            .O(N__14642),
            .I(N__14639));
    LocalMux I__3261 (
            .O(N__14639),
            .I(N__14632));
    SRMux I__3260 (
            .O(N__14638),
            .I(N__14629));
    SRMux I__3259 (
            .O(N__14637),
            .I(N__14626));
    SRMux I__3258 (
            .O(N__14636),
            .I(N__14623));
    SRMux I__3257 (
            .O(N__14635),
            .I(N__14620));
    Span4Mux_v I__3256 (
            .O(N__14632),
            .I(N__14617));
    LocalMux I__3255 (
            .O(N__14629),
            .I(N__14614));
    LocalMux I__3254 (
            .O(N__14626),
            .I(N__14607));
    LocalMux I__3253 (
            .O(N__14623),
            .I(N__14607));
    LocalMux I__3252 (
            .O(N__14620),
            .I(N__14607));
    Odrv4 I__3251 (
            .O(N__14617),
            .I(\uart_inst0.uart_inst0.un1_rx_state49_i ));
    Odrv4 I__3250 (
            .O(N__14614),
            .I(\uart_inst0.uart_inst0.un1_rx_state49_i ));
    Odrv4 I__3249 (
            .O(N__14607),
            .I(\uart_inst0.uart_inst0.un1_rx_state49_i ));
    InMux I__3248 (
            .O(N__14600),
            .I(N__14594));
    InMux I__3247 (
            .O(N__14599),
            .I(N__14594));
    LocalMux I__3246 (
            .O(N__14594),
            .I(N__14587));
    InMux I__3245 (
            .O(N__14593),
            .I(N__14584));
    InMux I__3244 (
            .O(N__14592),
            .I(N__14581));
    InMux I__3243 (
            .O(N__14591),
            .I(N__14578));
    InMux I__3242 (
            .O(N__14590),
            .I(N__14575));
    Span4Mux_h I__3241 (
            .O(N__14587),
            .I(N__14572));
    LocalMux I__3240 (
            .O(N__14584),
            .I(N__14569));
    LocalMux I__3239 (
            .O(N__14581),
            .I(N__14566));
    LocalMux I__3238 (
            .O(N__14578),
            .I(\uart_inst0.uart_inst0.tx_countdownZ0Z_1 ));
    LocalMux I__3237 (
            .O(N__14575),
            .I(\uart_inst0.uart_inst0.tx_countdownZ0Z_1 ));
    Odrv4 I__3236 (
            .O(N__14572),
            .I(\uart_inst0.uart_inst0.tx_countdownZ0Z_1 ));
    Odrv12 I__3235 (
            .O(N__14569),
            .I(\uart_inst0.uart_inst0.tx_countdownZ0Z_1 ));
    Odrv4 I__3234 (
            .O(N__14566),
            .I(\uart_inst0.uart_inst0.tx_countdownZ0Z_1 ));
    InMux I__3233 (
            .O(N__14555),
            .I(N__14552));
    LocalMux I__3232 (
            .O(N__14552),
            .I(N__14544));
    InMux I__3231 (
            .O(N__14551),
            .I(N__14540));
    InMux I__3230 (
            .O(N__14550),
            .I(N__14537));
    InMux I__3229 (
            .O(N__14549),
            .I(N__14532));
    InMux I__3228 (
            .O(N__14548),
            .I(N__14532));
    InMux I__3227 (
            .O(N__14547),
            .I(N__14529));
    Span4Mux_h I__3226 (
            .O(N__14544),
            .I(N__14526));
    InMux I__3225 (
            .O(N__14543),
            .I(N__14523));
    LocalMux I__3224 (
            .O(N__14540),
            .I(N__14520));
    LocalMux I__3223 (
            .O(N__14537),
            .I(N__14517));
    LocalMux I__3222 (
            .O(N__14532),
            .I(\uart_inst0.uart_inst0.tx_countdownZ0Z_0 ));
    LocalMux I__3221 (
            .O(N__14529),
            .I(\uart_inst0.uart_inst0.tx_countdownZ0Z_0 ));
    Odrv4 I__3220 (
            .O(N__14526),
            .I(\uart_inst0.uart_inst0.tx_countdownZ0Z_0 ));
    LocalMux I__3219 (
            .O(N__14523),
            .I(\uart_inst0.uart_inst0.tx_countdownZ0Z_0 ));
    Odrv4 I__3218 (
            .O(N__14520),
            .I(\uart_inst0.uart_inst0.tx_countdownZ0Z_0 ));
    Odrv4 I__3217 (
            .O(N__14517),
            .I(\uart_inst0.uart_inst0.tx_countdownZ0Z_0 ));
    InMux I__3216 (
            .O(N__14504),
            .I(N__14501));
    LocalMux I__3215 (
            .O(N__14501),
            .I(N__14497));
    InMux I__3214 (
            .O(N__14500),
            .I(N__14494));
    Odrv4 I__3213 (
            .O(N__14497),
            .I(\uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_9 ));
    LocalMux I__3212 (
            .O(N__14494),
            .I(\uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_9 ));
    InMux I__3211 (
            .O(N__14489),
            .I(N__14486));
    LocalMux I__3210 (
            .O(N__14486),
            .I(N__14483));
    Odrv4 I__3209 (
            .O(N__14483),
            .I(\uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_11_3 ));
    CascadeMux I__3208 (
            .O(N__14480),
            .I(\uart_inst0.uart_inst0.tx_m5_0_2_cascade_ ));
    InMux I__3207 (
            .O(N__14477),
            .I(N__14474));
    LocalMux I__3206 (
            .O(N__14474),
            .I(N__14471));
    Span4Mux_v I__3205 (
            .O(N__14471),
            .I(N__14467));
    InMux I__3204 (
            .O(N__14470),
            .I(N__14464));
    Odrv4 I__3203 (
            .O(N__14467),
            .I(\uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_11_4 ));
    LocalMux I__3202 (
            .O(N__14464),
            .I(\uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_11_4 ));
    InMux I__3201 (
            .O(N__14459),
            .I(N__14456));
    LocalMux I__3200 (
            .O(N__14456),
            .I(N__14453));
    Odrv4 I__3199 (
            .O(N__14453),
            .I(\uart_inst0.uart_inst0.tx_N_11_mux ));
    InMux I__3198 (
            .O(N__14450),
            .I(N__14445));
    InMux I__3197 (
            .O(N__14449),
            .I(N__14442));
    InMux I__3196 (
            .O(N__14448),
            .I(N__14439));
    LocalMux I__3195 (
            .O(N__14445),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_2 ));
    LocalMux I__3194 (
            .O(N__14442),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_2 ));
    LocalMux I__3193 (
            .O(N__14439),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_2 ));
    InMux I__3192 (
            .O(N__14432),
            .I(N__14428));
    InMux I__3191 (
            .O(N__14431),
            .I(N__14425));
    LocalMux I__3190 (
            .O(N__14428),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_0 ));
    LocalMux I__3189 (
            .O(N__14425),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_0 ));
    CascadeMux I__3188 (
            .O(N__14420),
            .I(N__14415));
    InMux I__3187 (
            .O(N__14419),
            .I(N__14412));
    InMux I__3186 (
            .O(N__14418),
            .I(N__14409));
    InMux I__3185 (
            .O(N__14415),
            .I(N__14406));
    LocalMux I__3184 (
            .O(N__14412),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_3 ));
    LocalMux I__3183 (
            .O(N__14409),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_3 ));
    LocalMux I__3182 (
            .O(N__14406),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_3 ));
    InMux I__3181 (
            .O(N__14399),
            .I(N__14394));
    InMux I__3180 (
            .O(N__14398),
            .I(N__14391));
    InMux I__3179 (
            .O(N__14397),
            .I(N__14388));
    LocalMux I__3178 (
            .O(N__14394),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_1 ));
    LocalMux I__3177 (
            .O(N__14391),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_1 ));
    LocalMux I__3176 (
            .O(N__14388),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_1 ));
    InMux I__3175 (
            .O(N__14381),
            .I(N__14377));
    InMux I__3174 (
            .O(N__14380),
            .I(N__14374));
    LocalMux I__3173 (
            .O(N__14377),
            .I(N__14371));
    LocalMux I__3172 (
            .O(N__14374),
            .I(\uart_inst0.uart_inst0.tx_m5_0 ));
    Odrv4 I__3171 (
            .O(N__14371),
            .I(\uart_inst0.uart_inst0.tx_m5_0 ));
    InMux I__3170 (
            .O(N__14366),
            .I(N__14363));
    LocalMux I__3169 (
            .O(N__14363),
            .I(ioFifoData_in_5));
    InMux I__3168 (
            .O(N__14360),
            .I(N__14357));
    LocalMux I__3167 (
            .O(N__14357),
            .I(N__14353));
    InMux I__3166 (
            .O(N__14356),
            .I(N__14350));
    Span4Mux_h I__3165 (
            .O(N__14353),
            .I(N__14347));
    LocalMux I__3164 (
            .O(N__14350),
            .I(\fifo_inst.wRxWrData_5 ));
    Odrv4 I__3163 (
            .O(N__14347),
            .I(\fifo_inst.wRxWrData_5 ));
    CascadeMux I__3162 (
            .O(N__14342),
            .I(N__14339));
    InMux I__3161 (
            .O(N__14339),
            .I(N__14336));
    LocalMux I__3160 (
            .O(N__14336),
            .I(N__14333));
    Span4Mux_h I__3159 (
            .O(N__14333),
            .I(N__14328));
    InMux I__3158 (
            .O(N__14332),
            .I(N__14325));
    InMux I__3157 (
            .O(N__14331),
            .I(N__14322));
    Odrv4 I__3156 (
            .O(N__14328),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_5));
    LocalMux I__3155 (
            .O(N__14325),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_5));
    LocalMux I__3154 (
            .O(N__14322),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_5));
    CascadeMux I__3153 (
            .O(N__14315),
            .I(N__14312));
    InMux I__3152 (
            .O(N__14312),
            .I(N__14309));
    LocalMux I__3151 (
            .O(N__14309),
            .I(N__14304));
    InMux I__3150 (
            .O(N__14308),
            .I(N__14301));
    InMux I__3149 (
            .O(N__14307),
            .I(N__14298));
    Span4Mux_h I__3148 (
            .O(N__14304),
            .I(N__14295));
    LocalMux I__3147 (
            .O(N__14301),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_4));
    LocalMux I__3146 (
            .O(N__14298),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_4));
    Odrv4 I__3145 (
            .O(N__14295),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_4));
    CascadeMux I__3144 (
            .O(N__14288),
            .I(N__14284));
    CascadeMux I__3143 (
            .O(N__14287),
            .I(N__14281));
    InMux I__3142 (
            .O(N__14284),
            .I(N__14278));
    InMux I__3141 (
            .O(N__14281),
            .I(N__14275));
    LocalMux I__3140 (
            .O(N__14278),
            .I(N__14271));
    LocalMux I__3139 (
            .O(N__14275),
            .I(N__14268));
    InMux I__3138 (
            .O(N__14274),
            .I(N__14265));
    Span4Mux_v I__3137 (
            .O(N__14271),
            .I(N__14262));
    Odrv4 I__3136 (
            .O(N__14268),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_2));
    LocalMux I__3135 (
            .O(N__14265),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_2));
    Odrv4 I__3134 (
            .O(N__14262),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_2));
    CascadeMux I__3133 (
            .O(N__14255),
            .I(N__14252));
    InMux I__3132 (
            .O(N__14252),
            .I(N__14249));
    LocalMux I__3131 (
            .O(N__14249),
            .I(N__14245));
    InMux I__3130 (
            .O(N__14248),
            .I(N__14241));
    Span4Mux_h I__3129 (
            .O(N__14245),
            .I(N__14238));
    InMux I__3128 (
            .O(N__14244),
            .I(N__14235));
    LocalMux I__3127 (
            .O(N__14241),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_7));
    Odrv4 I__3126 (
            .O(N__14238),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_7));
    LocalMux I__3125 (
            .O(N__14235),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_7));
    CascadeMux I__3124 (
            .O(N__14228),
            .I(N__14225));
    InMux I__3123 (
            .O(N__14225),
            .I(N__14222));
    LocalMux I__3122 (
            .O(N__14222),
            .I(N__14219));
    Span4Mux_h I__3121 (
            .O(N__14219),
            .I(N__14214));
    InMux I__3120 (
            .O(N__14218),
            .I(N__14211));
    InMux I__3119 (
            .O(N__14217),
            .I(N__14208));
    Odrv4 I__3118 (
            .O(N__14214),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_6));
    LocalMux I__3117 (
            .O(N__14211),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_6));
    LocalMux I__3116 (
            .O(N__14208),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_6));
    CascadeMux I__3115 (
            .O(N__14201),
            .I(\uart_inst0.tx_uart_fifo_inst.m54_eZ0Z_5_cascade_ ));
    CascadeMux I__3114 (
            .O(N__14198),
            .I(\uart_inst0.tx_uart_fifo_inst.N_91_cascade_ ));
    InMux I__3113 (
            .O(N__14195),
            .I(N__14192));
    LocalMux I__3112 (
            .O(N__14192),
            .I(un1_rRamWrAddr_cry_2_c_RNIOTMG));
    CascadeMux I__3111 (
            .O(N__14189),
            .I(N__14186));
    InMux I__3110 (
            .O(N__14186),
            .I(N__14183));
    LocalMux I__3109 (
            .O(N__14183),
            .I(N__14178));
    InMux I__3108 (
            .O(N__14182),
            .I(N__14175));
    InMux I__3107 (
            .O(N__14181),
            .I(N__14172));
    Odrv4 I__3106 (
            .O(N__14178),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_3));
    LocalMux I__3105 (
            .O(N__14175),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_3));
    LocalMux I__3104 (
            .O(N__14172),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_3));
    CascadeMux I__3103 (
            .O(N__14165),
            .I(N__14162));
    InMux I__3102 (
            .O(N__14162),
            .I(N__14159));
    LocalMux I__3101 (
            .O(N__14159),
            .I(N__14156));
    Span4Mux_h I__3100 (
            .O(N__14156),
            .I(N__14151));
    InMux I__3099 (
            .O(N__14155),
            .I(N__14148));
    InMux I__3098 (
            .O(N__14154),
            .I(N__14145));
    Odrv4 I__3097 (
            .O(N__14151),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_1));
    LocalMux I__3096 (
            .O(N__14148),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_1));
    LocalMux I__3095 (
            .O(N__14145),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_1));
    CascadeMux I__3094 (
            .O(N__14138),
            .I(N__14135));
    InMux I__3093 (
            .O(N__14135),
            .I(N__14132));
    LocalMux I__3092 (
            .O(N__14132),
            .I(N__14127));
    CascadeMux I__3091 (
            .O(N__14131),
            .I(N__14124));
    InMux I__3090 (
            .O(N__14130),
            .I(N__14121));
    Span4Mux_h I__3089 (
            .O(N__14127),
            .I(N__14118));
    InMux I__3088 (
            .O(N__14124),
            .I(N__14115));
    LocalMux I__3087 (
            .O(N__14121),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_8));
    Odrv4 I__3086 (
            .O(N__14118),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_8));
    LocalMux I__3085 (
            .O(N__14115),
            .I(fifo_inst_rx_fifo_inst_rRamWrAddr_8));
    InMux I__3084 (
            .O(N__14108),
            .I(N__14105));
    LocalMux I__3083 (
            .O(N__14105),
            .I(\uart_inst0.tx_uart_fifo_inst.m54_eZ0Z_6 ));
    InMux I__3082 (
            .O(N__14102),
            .I(N__14097));
    IoInMux I__3081 (
            .O(N__14101),
            .I(N__14094));
    InMux I__3080 (
            .O(N__14100),
            .I(N__14091));
    LocalMux I__3079 (
            .O(N__14097),
            .I(N__14088));
    LocalMux I__3078 (
            .O(N__14094),
            .I(N__14085));
    LocalMux I__3077 (
            .O(N__14091),
            .I(N__14082));
    Span4Mux_h I__3076 (
            .O(N__14088),
            .I(N__14078));
    IoSpan4Mux I__3075 (
            .O(N__14085),
            .I(N__14075));
    Span4Mux_v I__3074 (
            .O(N__14082),
            .I(N__14072));
    InMux I__3073 (
            .O(N__14081),
            .I(N__14069));
    Span4Mux_h I__3072 (
            .O(N__14078),
            .I(N__14063));
    Span4Mux_s2_v I__3071 (
            .O(N__14075),
            .I(N__14063));
    Span4Mux_v I__3070 (
            .O(N__14072),
            .I(N__14058));
    LocalMux I__3069 (
            .O(N__14069),
            .I(N__14058));
    InMux I__3068 (
            .O(N__14068),
            .I(N__14055));
    Sp12to4 I__3067 (
            .O(N__14063),
            .I(N__14052));
    Span4Mux_v I__3066 (
            .O(N__14058),
            .I(N__14049));
    LocalMux I__3065 (
            .O(N__14055),
            .I(N__14046));
    Span12Mux_v I__3064 (
            .O(N__14052),
            .I(N__14039));
    Sp12to4 I__3063 (
            .O(N__14049),
            .I(N__14039));
    Sp12to4 I__3062 (
            .O(N__14046),
            .I(N__14039));
    Odrv12 I__3061 (
            .O(N__14039),
            .I(wPllLocked_i));
    InMux I__3060 (
            .O(N__14036),
            .I(N__14032));
    InMux I__3059 (
            .O(N__14035),
            .I(N__14029));
    LocalMux I__3058 (
            .O(N__14032),
            .I(\uart_inst0.uart_inst0.rRxData_0_sqmuxa ));
    LocalMux I__3057 (
            .O(N__14029),
            .I(\uart_inst0.uart_inst0.rRxData_0_sqmuxa ));
    InMux I__3056 (
            .O(N__14024),
            .I(N__14017));
    InMux I__3055 (
            .O(N__14023),
            .I(N__14006));
    InMux I__3054 (
            .O(N__14022),
            .I(N__14006));
    CascadeMux I__3053 (
            .O(N__14021),
            .I(N__14000));
    InMux I__3052 (
            .O(N__14020),
            .I(N__13995));
    LocalMux I__3051 (
            .O(N__14017),
            .I(N__13992));
    InMux I__3050 (
            .O(N__14016),
            .I(N__13987));
    InMux I__3049 (
            .O(N__14015),
            .I(N__13987));
    InMux I__3048 (
            .O(N__14014),
            .I(N__13983));
    CascadeMux I__3047 (
            .O(N__14013),
            .I(N__13980));
    CascadeMux I__3046 (
            .O(N__14012),
            .I(N__13977));
    CascadeMux I__3045 (
            .O(N__14011),
            .I(N__13974));
    LocalMux I__3044 (
            .O(N__14006),
            .I(N__13971));
    InMux I__3043 (
            .O(N__14005),
            .I(N__13968));
    InMux I__3042 (
            .O(N__14004),
            .I(N__13963));
    InMux I__3041 (
            .O(N__14003),
            .I(N__13963));
    InMux I__3040 (
            .O(N__14000),
            .I(N__13956));
    InMux I__3039 (
            .O(N__13999),
            .I(N__13956));
    InMux I__3038 (
            .O(N__13998),
            .I(N__13956));
    LocalMux I__3037 (
            .O(N__13995),
            .I(N__13953));
    Span4Mux_v I__3036 (
            .O(N__13992),
            .I(N__13950));
    LocalMux I__3035 (
            .O(N__13987),
            .I(N__13947));
    CascadeMux I__3034 (
            .O(N__13986),
            .I(N__13943));
    LocalMux I__3033 (
            .O(N__13983),
            .I(N__13940));
    InMux I__3032 (
            .O(N__13980),
            .I(N__13937));
    InMux I__3031 (
            .O(N__13977),
            .I(N__13932));
    InMux I__3030 (
            .O(N__13974),
            .I(N__13932));
    Span4Mux_v I__3029 (
            .O(N__13971),
            .I(N__13929));
    LocalMux I__3028 (
            .O(N__13968),
            .I(N__13922));
    LocalMux I__3027 (
            .O(N__13963),
            .I(N__13922));
    LocalMux I__3026 (
            .O(N__13956),
            .I(N__13922));
    Span4Mux_s3_v I__3025 (
            .O(N__13953),
            .I(N__13918));
    Span4Mux_h I__3024 (
            .O(N__13950),
            .I(N__13913));
    Span4Mux_v I__3023 (
            .O(N__13947),
            .I(N__13913));
    InMux I__3022 (
            .O(N__13946),
            .I(N__13910));
    InMux I__3021 (
            .O(N__13943),
            .I(N__13907));
    Span4Mux_v I__3020 (
            .O(N__13940),
            .I(N__13904));
    LocalMux I__3019 (
            .O(N__13937),
            .I(N__13895));
    LocalMux I__3018 (
            .O(N__13932),
            .I(N__13895));
    Span4Mux_h I__3017 (
            .O(N__13929),
            .I(N__13895));
    Span4Mux_v I__3016 (
            .O(N__13922),
            .I(N__13895));
    InMux I__3015 (
            .O(N__13921),
            .I(N__13891));
    Span4Mux_h I__3014 (
            .O(N__13918),
            .I(N__13888));
    Span4Mux_v I__3013 (
            .O(N__13913),
            .I(N__13885));
    LocalMux I__3012 (
            .O(N__13910),
            .I(N__13880));
    LocalMux I__3011 (
            .O(N__13907),
            .I(N__13880));
    Span4Mux_h I__3010 (
            .O(N__13904),
            .I(N__13875));
    Span4Mux_h I__3009 (
            .O(N__13895),
            .I(N__13875));
    InMux I__3008 (
            .O(N__13894),
            .I(N__13872));
    LocalMux I__3007 (
            .O(N__13891),
            .I(N__13869));
    Sp12to4 I__3006 (
            .O(N__13888),
            .I(N__13866));
    Sp12to4 I__3005 (
            .O(N__13885),
            .I(N__13857));
    Span12Mux_h I__3004 (
            .O(N__13880),
            .I(N__13857));
    Sp12to4 I__3003 (
            .O(N__13875),
            .I(N__13857));
    LocalMux I__3002 (
            .O(N__13872),
            .I(N__13857));
    Span4Mux_v I__3001 (
            .O(N__13869),
            .I(N__13854));
    Span12Mux_v I__3000 (
            .O(N__13866),
            .I(N__13851));
    Span12Mux_h I__2999 (
            .O(N__13857),
            .I(N__13848));
    Sp12to4 I__2998 (
            .O(N__13854),
            .I(N__13845));
    Span12Mux_h I__2997 (
            .O(N__13851),
            .I(N__13842));
    Span12Mux_v I__2996 (
            .O(N__13848),
            .I(N__13839));
    Span12Mux_v I__2995 (
            .O(N__13845),
            .I(N__13836));
    Odrv12 I__2994 (
            .O(N__13842),
            .I(wPllLocked));
    Odrv12 I__2993 (
            .O(N__13839),
            .I(wPllLocked));
    Odrv12 I__2992 (
            .O(N__13836),
            .I(wPllLocked));
    InMux I__2991 (
            .O(N__13829),
            .I(N__13826));
    LocalMux I__2990 (
            .O(N__13826),
            .I(N__13819));
    InMux I__2989 (
            .O(N__13825),
            .I(N__13814));
    InMux I__2988 (
            .O(N__13824),
            .I(N__13807));
    InMux I__2987 (
            .O(N__13823),
            .I(N__13807));
    InMux I__2986 (
            .O(N__13822),
            .I(N__13807));
    Span4Mux_h I__2985 (
            .O(N__13819),
            .I(N__13804));
    InMux I__2984 (
            .O(N__13818),
            .I(N__13799));
    InMux I__2983 (
            .O(N__13817),
            .I(N__13799));
    LocalMux I__2982 (
            .O(N__13814),
            .I(\uart_inst0.uart_inst0.N_257_0 ));
    LocalMux I__2981 (
            .O(N__13807),
            .I(\uart_inst0.uart_inst0.N_257_0 ));
    Odrv4 I__2980 (
            .O(N__13804),
            .I(\uart_inst0.uart_inst0.N_257_0 ));
    LocalMux I__2979 (
            .O(N__13799),
            .I(\uart_inst0.uart_inst0.N_257_0 ));
    CascadeMux I__2978 (
            .O(N__13790),
            .I(\uart_inst0.uart_inst0.N_273_cascade_ ));
    CascadeMux I__2977 (
            .O(N__13787),
            .I(N__13784));
    InMux I__2976 (
            .O(N__13784),
            .I(N__13781));
    LocalMux I__2975 (
            .O(N__13781),
            .I(N__13775));
    InMux I__2974 (
            .O(N__13780),
            .I(N__13772));
    InMux I__2973 (
            .O(N__13779),
            .I(N__13768));
    InMux I__2972 (
            .O(N__13778),
            .I(N__13765));
    Span4Mux_v I__2971 (
            .O(N__13775),
            .I(N__13762));
    LocalMux I__2970 (
            .O(N__13772),
            .I(N__13759));
    InMux I__2969 (
            .O(N__13771),
            .I(N__13756));
    LocalMux I__2968 (
            .O(N__13768),
            .I(N__13749));
    LocalMux I__2967 (
            .O(N__13765),
            .I(N__13749));
    Span4Mux_h I__2966 (
            .O(N__13762),
            .I(N__13749));
    Span4Mux_h I__2965 (
            .O(N__13759),
            .I(N__13746));
    LocalMux I__2964 (
            .O(N__13756),
            .I(\uart_inst0.uart_inst0.rx_stateZ0Z_3 ));
    Odrv4 I__2963 (
            .O(N__13749),
            .I(\uart_inst0.uart_inst0.rx_stateZ0Z_3 ));
    Odrv4 I__2962 (
            .O(N__13746),
            .I(\uart_inst0.uart_inst0.rx_stateZ0Z_3 ));
    InMux I__2961 (
            .O(N__13739),
            .I(N__13735));
    InMux I__2960 (
            .O(N__13738),
            .I(N__13732));
    LocalMux I__2959 (
            .O(N__13735),
            .I(N__13729));
    LocalMux I__2958 (
            .O(N__13732),
            .I(\uart_inst0.uart_inst0.rx_state_srsts_0_a5_0_0_3 ));
    Odrv4 I__2957 (
            .O(N__13729),
            .I(\uart_inst0.uart_inst0.rx_state_srsts_0_a5_0_0_3 ));
    InMux I__2956 (
            .O(N__13724),
            .I(N__13721));
    LocalMux I__2955 (
            .O(N__13721),
            .I(N__13716));
    InMux I__2954 (
            .O(N__13720),
            .I(N__13713));
    InMux I__2953 (
            .O(N__13719),
            .I(N__13710));
    Span4Mux_v I__2952 (
            .O(N__13716),
            .I(N__13707));
    LocalMux I__2951 (
            .O(N__13713),
            .I(\uart_inst0.uart_inst0.N_274_2 ));
    LocalMux I__2950 (
            .O(N__13710),
            .I(\uart_inst0.uart_inst0.N_274_2 ));
    Odrv4 I__2949 (
            .O(N__13707),
            .I(\uart_inst0.uart_inst0.N_274_2 ));
    CascadeMux I__2948 (
            .O(N__13700),
            .I(\uart_inst0.uart_inst0.un1_rx_bits_remaining_c3_cascade_ ));
    InMux I__2947 (
            .O(N__13697),
            .I(N__13693));
    InMux I__2946 (
            .O(N__13696),
            .I(N__13690));
    LocalMux I__2945 (
            .O(N__13693),
            .I(\uart_inst0.uart_inst0.rx_bits_remainingZ0Z_3 ));
    LocalMux I__2944 (
            .O(N__13690),
            .I(\uart_inst0.uart_inst0.rx_bits_remainingZ0Z_3 ));
    InMux I__2943 (
            .O(N__13685),
            .I(N__13681));
    CascadeMux I__2942 (
            .O(N__13684),
            .I(N__13676));
    LocalMux I__2941 (
            .O(N__13681),
            .I(N__13673));
    CascadeMux I__2940 (
            .O(N__13680),
            .I(N__13670));
    CascadeMux I__2939 (
            .O(N__13679),
            .I(N__13667));
    InMux I__2938 (
            .O(N__13676),
            .I(N__13664));
    Span4Mux_h I__2937 (
            .O(N__13673),
            .I(N__13661));
    InMux I__2936 (
            .O(N__13670),
            .I(N__13658));
    InMux I__2935 (
            .O(N__13667),
            .I(N__13655));
    LocalMux I__2934 (
            .O(N__13664),
            .I(N__13652));
    Odrv4 I__2933 (
            .O(N__13661),
            .I(\uart_inst0.uart_inst0.tx_countdownZ0Z_3 ));
    LocalMux I__2932 (
            .O(N__13658),
            .I(\uart_inst0.uart_inst0.tx_countdownZ0Z_3 ));
    LocalMux I__2931 (
            .O(N__13655),
            .I(\uart_inst0.uart_inst0.tx_countdownZ0Z_3 ));
    Odrv4 I__2930 (
            .O(N__13652),
            .I(\uart_inst0.uart_inst0.tx_countdownZ0Z_3 ));
    CascadeMux I__2929 (
            .O(N__13643),
            .I(N__13640));
    InMux I__2928 (
            .O(N__13640),
            .I(N__13637));
    LocalMux I__2927 (
            .O(N__13637),
            .I(\uart_inst0.uart_inst0.tx_N_2 ));
    InMux I__2926 (
            .O(N__13634),
            .I(N__13631));
    LocalMux I__2925 (
            .O(N__13631),
            .I(N__13625));
    InMux I__2924 (
            .O(N__13630),
            .I(N__13622));
    InMux I__2923 (
            .O(N__13629),
            .I(N__13619));
    InMux I__2922 (
            .O(N__13628),
            .I(N__13616));
    Span4Mux_v I__2921 (
            .O(N__13625),
            .I(N__13611));
    LocalMux I__2920 (
            .O(N__13622),
            .I(N__13611));
    LocalMux I__2919 (
            .O(N__13619),
            .I(\uart_inst0.uart_inst0.tx_countdownZ0Z_2 ));
    LocalMux I__2918 (
            .O(N__13616),
            .I(\uart_inst0.uart_inst0.tx_countdownZ0Z_2 ));
    Odrv4 I__2917 (
            .O(N__13611),
            .I(\uart_inst0.uart_inst0.tx_countdownZ0Z_2 ));
    SRMux I__2916 (
            .O(N__13604),
            .I(N__13562));
    SRMux I__2915 (
            .O(N__13603),
            .I(N__13562));
    SRMux I__2914 (
            .O(N__13602),
            .I(N__13562));
    SRMux I__2913 (
            .O(N__13601),
            .I(N__13562));
    SRMux I__2912 (
            .O(N__13600),
            .I(N__13562));
    SRMux I__2911 (
            .O(N__13599),
            .I(N__13562));
    SRMux I__2910 (
            .O(N__13598),
            .I(N__13562));
    SRMux I__2909 (
            .O(N__13597),
            .I(N__13562));
    SRMux I__2908 (
            .O(N__13596),
            .I(N__13562));
    SRMux I__2907 (
            .O(N__13595),
            .I(N__13562));
    SRMux I__2906 (
            .O(N__13594),
            .I(N__13562));
    SRMux I__2905 (
            .O(N__13593),
            .I(N__13562));
    SRMux I__2904 (
            .O(N__13592),
            .I(N__13562));
    SRMux I__2903 (
            .O(N__13591),
            .I(N__13562));
    GlobalMux I__2902 (
            .O(N__13562),
            .I(N__13559));
    gio2CtrlBuf I__2901 (
            .O(N__13559),
            .I(N_292_g));
    CascadeMux I__2900 (
            .O(N__13556),
            .I(N__13551));
    InMux I__2899 (
            .O(N__13555),
            .I(N__13538));
    InMux I__2898 (
            .O(N__13554),
            .I(N__13529));
    InMux I__2897 (
            .O(N__13551),
            .I(N__13529));
    InMux I__2896 (
            .O(N__13550),
            .I(N__13529));
    InMux I__2895 (
            .O(N__13549),
            .I(N__13529));
    InMux I__2894 (
            .O(N__13548),
            .I(N__13526));
    InMux I__2893 (
            .O(N__13547),
            .I(N__13511));
    InMux I__2892 (
            .O(N__13546),
            .I(N__13511));
    InMux I__2891 (
            .O(N__13545),
            .I(N__13511));
    InMux I__2890 (
            .O(N__13544),
            .I(N__13511));
    InMux I__2889 (
            .O(N__13543),
            .I(N__13511));
    InMux I__2888 (
            .O(N__13542),
            .I(N__13511));
    InMux I__2887 (
            .O(N__13541),
            .I(N__13511));
    LocalMux I__2886 (
            .O(N__13538),
            .I(N__13505));
    LocalMux I__2885 (
            .O(N__13529),
            .I(N__13505));
    LocalMux I__2884 (
            .O(N__13526),
            .I(N__13500));
    LocalMux I__2883 (
            .O(N__13511),
            .I(N__13500));
    InMux I__2882 (
            .O(N__13510),
            .I(N__13497));
    Odrv4 I__2881 (
            .O(N__13505),
            .I(\uart_inst0.uart_inst0.N_147_0_i ));
    Odrv4 I__2880 (
            .O(N__13500),
            .I(\uart_inst0.uart_inst0.N_147_0_i ));
    LocalMux I__2879 (
            .O(N__13497),
            .I(\uart_inst0.uart_inst0.N_147_0_i ));
    InMux I__2878 (
            .O(N__13490),
            .I(N__13487));
    LocalMux I__2877 (
            .O(N__13487),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_2_s1_THRU_CO ));
    InMux I__2876 (
            .O(N__13484),
            .I(N__13480));
    InMux I__2875 (
            .O(N__13483),
            .I(N__13477));
    LocalMux I__2874 (
            .O(N__13480),
            .I(N__13472));
    LocalMux I__2873 (
            .O(N__13477),
            .I(N__13472));
    Odrv4 I__2872 (
            .O(N__13472),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIOAZ0Z54 ));
    CascadeMux I__2871 (
            .O(N__13469),
            .I(N__13466));
    InMux I__2870 (
            .O(N__13466),
            .I(N__13463));
    LocalMux I__2869 (
            .O(N__13463),
            .I(N__13460));
    Odrv4 I__2868 (
            .O(N__13460),
            .I(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_0 ));
    CascadeMux I__2867 (
            .O(N__13457),
            .I(N__13453));
    InMux I__2866 (
            .O(N__13456),
            .I(N__13450));
    InMux I__2865 (
            .O(N__13453),
            .I(N__13447));
    LocalMux I__2864 (
            .O(N__13450),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_6 ));
    LocalMux I__2863 (
            .O(N__13447),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_6 ));
    InMux I__2862 (
            .O(N__13442),
            .I(N__13438));
    InMux I__2861 (
            .O(N__13441),
            .I(N__13435));
    LocalMux I__2860 (
            .O(N__13438),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_5 ));
    LocalMux I__2859 (
            .O(N__13435),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_5 ));
    CascadeMux I__2858 (
            .O(N__13430),
            .I(N__13427));
    InMux I__2857 (
            .O(N__13427),
            .I(N__13423));
    InMux I__2856 (
            .O(N__13426),
            .I(N__13420));
    LocalMux I__2855 (
            .O(N__13423),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_7 ));
    LocalMux I__2854 (
            .O(N__13420),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_7 ));
    InMux I__2853 (
            .O(N__13415),
            .I(N__13411));
    InMux I__2852 (
            .O(N__13414),
            .I(N__13408));
    LocalMux I__2851 (
            .O(N__13411),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_4 ));
    LocalMux I__2850 (
            .O(N__13408),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_4 ));
    CascadeMux I__2849 (
            .O(N__13403),
            .I(N__13400));
    InMux I__2848 (
            .O(N__13400),
            .I(N__13397));
    LocalMux I__2847 (
            .O(N__13397),
            .I(\uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_5 ));
    InMux I__2846 (
            .O(N__13394),
            .I(N__13388));
    InMux I__2845 (
            .O(N__13393),
            .I(N__13388));
    LocalMux I__2844 (
            .O(N__13388),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_8 ));
    InMux I__2843 (
            .O(N__13385),
            .I(N__13382));
    LocalMux I__2842 (
            .O(N__13382),
            .I(\uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_4 ));
    CascadeMux I__2841 (
            .O(N__13379),
            .I(N__13376));
    InMux I__2840 (
            .O(N__13376),
            .I(N__13373));
    LocalMux I__2839 (
            .O(N__13373),
            .I(N__13367));
    InMux I__2838 (
            .O(N__13372),
            .I(N__13364));
    InMux I__2837 (
            .O(N__13371),
            .I(N__13359));
    InMux I__2836 (
            .O(N__13370),
            .I(N__13359));
    Odrv12 I__2835 (
            .O(N__13367),
            .I(wUartRxEmpty));
    LocalMux I__2834 (
            .O(N__13364),
            .I(wUartRxEmpty));
    LocalMux I__2833 (
            .O(N__13359),
            .I(wUartRxEmpty));
    InMux I__2832 (
            .O(N__13352),
            .I(N__13348));
    InMux I__2831 (
            .O(N__13351),
            .I(N__13345));
    LocalMux I__2830 (
            .O(N__13348),
            .I(N__13342));
    LocalMux I__2829 (
            .O(N__13345),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_0 ));
    Odrv4 I__2828 (
            .O(N__13342),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_0 ));
    CascadeMux I__2827 (
            .O(N__13337),
            .I(N__13334));
    InMux I__2826 (
            .O(N__13334),
            .I(N__13330));
    InMux I__2825 (
            .O(N__13333),
            .I(N__13327));
    LocalMux I__2824 (
            .O(N__13330),
            .I(N__13324));
    LocalMux I__2823 (
            .O(N__13327),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_3 ));
    Odrv4 I__2822 (
            .O(N__13324),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_3 ));
    CascadeMux I__2821 (
            .O(N__13319),
            .I(N__13312));
    InMux I__2820 (
            .O(N__13318),
            .I(N__13309));
    InMux I__2819 (
            .O(N__13317),
            .I(N__13304));
    InMux I__2818 (
            .O(N__13316),
            .I(N__13304));
    InMux I__2817 (
            .O(N__13315),
            .I(N__13299));
    InMux I__2816 (
            .O(N__13312),
            .I(N__13299));
    LocalMux I__2815 (
            .O(N__13309),
            .I(N__13291));
    LocalMux I__2814 (
            .O(N__13304),
            .I(N__13291));
    LocalMux I__2813 (
            .O(N__13299),
            .I(N__13291));
    InMux I__2812 (
            .O(N__13298),
            .I(N__13287));
    Span4Mux_v I__2811 (
            .O(N__13291),
            .I(N__13284));
    InMux I__2810 (
            .O(N__13290),
            .I(N__13281));
    LocalMux I__2809 (
            .O(N__13287),
            .I(N__13274));
    Sp12to4 I__2808 (
            .O(N__13284),
            .I(N__13274));
    LocalMux I__2807 (
            .O(N__13281),
            .I(N__13274));
    Span12Mux_h I__2806 (
            .O(N__13274),
            .I(N__13271));
    Span12Mux_v I__2805 (
            .O(N__13271),
            .I(N__13268));
    Odrv12 I__2804 (
            .O(N__13268),
            .I(P1A1_c));
    InMux I__2803 (
            .O(N__13265),
            .I(N__13260));
    CascadeMux I__2802 (
            .O(N__13264),
            .I(N__13255));
    CascadeMux I__2801 (
            .O(N__13263),
            .I(N__13251));
    LocalMux I__2800 (
            .O(N__13260),
            .I(N__13247));
    InMux I__2799 (
            .O(N__13259),
            .I(N__13242));
    InMux I__2798 (
            .O(N__13258),
            .I(N__13242));
    InMux I__2797 (
            .O(N__13255),
            .I(N__13239));
    InMux I__2796 (
            .O(N__13254),
            .I(N__13236));
    InMux I__2795 (
            .O(N__13251),
            .I(N__13231));
    InMux I__2794 (
            .O(N__13250),
            .I(N__13231));
    Span4Mux_h I__2793 (
            .O(N__13247),
            .I(N__13226));
    LocalMux I__2792 (
            .O(N__13242),
            .I(N__13226));
    LocalMux I__2791 (
            .O(N__13239),
            .I(\uart_inst0.uart_inst0.rx_stateZ0Z_1 ));
    LocalMux I__2790 (
            .O(N__13236),
            .I(\uart_inst0.uart_inst0.rx_stateZ0Z_1 ));
    LocalMux I__2789 (
            .O(N__13231),
            .I(\uart_inst0.uart_inst0.rx_stateZ0Z_1 ));
    Odrv4 I__2788 (
            .O(N__13226),
            .I(\uart_inst0.uart_inst0.rx_stateZ0Z_1 ));
    InMux I__2787 (
            .O(N__13217),
            .I(N__13213));
    InMux I__2786 (
            .O(N__13216),
            .I(N__13210));
    LocalMux I__2785 (
            .O(N__13213),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIK0HSZ0 ));
    LocalMux I__2784 (
            .O(N__13210),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIK0HSZ0 ));
    InMux I__2783 (
            .O(N__13205),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_0 ));
    InMux I__2782 (
            .O(N__13202),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_1 ));
    InMux I__2781 (
            .O(N__13199),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_2 ));
    InMux I__2780 (
            .O(N__13196),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_3 ));
    InMux I__2779 (
            .O(N__13193),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_4 ));
    InMux I__2778 (
            .O(N__13190),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_5 ));
    InMux I__2777 (
            .O(N__13187),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_6 ));
    InMux I__2776 (
            .O(N__13184),
            .I(bfn_17_11_0_));
    InMux I__2775 (
            .O(N__13181),
            .I(N__13177));
    InMux I__2774 (
            .O(N__13180),
            .I(N__13174));
    LocalMux I__2773 (
            .O(N__13177),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_1 ));
    LocalMux I__2772 (
            .O(N__13174),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_1 ));
    InMux I__2771 (
            .O(N__13169),
            .I(N__13165));
    InMux I__2770 (
            .O(N__13168),
            .I(N__13162));
    LocalMux I__2769 (
            .O(N__13165),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_2 ));
    LocalMux I__2768 (
            .O(N__13162),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_2 ));
    CascadeMux I__2767 (
            .O(N__13157),
            .I(N__13151));
    CascadeMux I__2766 (
            .O(N__13156),
            .I(N__13148));
    CEMux I__2765 (
            .O(N__13155),
            .I(N__13143));
    InMux I__2764 (
            .O(N__13154),
            .I(N__13137));
    InMux I__2763 (
            .O(N__13151),
            .I(N__13134));
    InMux I__2762 (
            .O(N__13148),
            .I(N__13131));
    InMux I__2761 (
            .O(N__13147),
            .I(N__13126));
    InMux I__2760 (
            .O(N__13146),
            .I(N__13126));
    LocalMux I__2759 (
            .O(N__13143),
            .I(N__13123));
    InMux I__2758 (
            .O(N__13142),
            .I(N__13118));
    InMux I__2757 (
            .O(N__13141),
            .I(N__13118));
    InMux I__2756 (
            .O(N__13140),
            .I(N__13115));
    LocalMux I__2755 (
            .O(N__13137),
            .I(N__13110));
    LocalMux I__2754 (
            .O(N__13134),
            .I(N__13110));
    LocalMux I__2753 (
            .O(N__13131),
            .I(N__13103));
    LocalMux I__2752 (
            .O(N__13126),
            .I(N__13103));
    Span4Mux_h I__2751 (
            .O(N__13123),
            .I(N__13103));
    LocalMux I__2750 (
            .O(N__13118),
            .I(\uart_inst0.rx_uart_fifo_inst.wRamWrEn ));
    LocalMux I__2749 (
            .O(N__13115),
            .I(\uart_inst0.rx_uart_fifo_inst.wRamWrEn ));
    Odrv4 I__2748 (
            .O(N__13110),
            .I(\uart_inst0.rx_uart_fifo_inst.wRamWrEn ));
    Odrv4 I__2747 (
            .O(N__13103),
            .I(\uart_inst0.rx_uart_fifo_inst.wRamWrEn ));
    InMux I__2746 (
            .O(N__13094),
            .I(N__13085));
    InMux I__2745 (
            .O(N__13093),
            .I(N__13082));
    InMux I__2744 (
            .O(N__13092),
            .I(N__13075));
    InMux I__2743 (
            .O(N__13091),
            .I(N__13075));
    InMux I__2742 (
            .O(N__13090),
            .I(N__13075));
    InMux I__2741 (
            .O(N__13089),
            .I(N__13070));
    InMux I__2740 (
            .O(N__13088),
            .I(N__13070));
    LocalMux I__2739 (
            .O(N__13085),
            .I(\uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_0 ));
    LocalMux I__2738 (
            .O(N__13082),
            .I(\uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_0 ));
    LocalMux I__2737 (
            .O(N__13075),
            .I(\uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_0 ));
    LocalMux I__2736 (
            .O(N__13070),
            .I(\uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_0 ));
    CascadeMux I__2735 (
            .O(N__13061),
            .I(\uart_inst0.rx_uart_fifo_inst.rDataCount_RNI3V391Z0Z_2_cascade_ ));
    InMux I__2734 (
            .O(N__13058),
            .I(N__13055));
    LocalMux I__2733 (
            .O(N__13055),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rDataCount15_2_0_0_0 ));
    CascadeMux I__2732 (
            .O(N__13052),
            .I(\uart_inst0.rx_uart_fifo_inst.wRamRdEn_cascade_ ));
    InMux I__2731 (
            .O(N__13049),
            .I(N__13046));
    LocalMux I__2730 (
            .O(N__13046),
            .I(N__13043));
    Span12Mux_s7_v I__2729 (
            .O(N__13043),
            .I(N__13037));
    InMux I__2728 (
            .O(N__13042),
            .I(N__13034));
    InMux I__2727 (
            .O(N__13041),
            .I(N__13031));
    InMux I__2726 (
            .O(N__13040),
            .I(N__13028));
    Odrv12 I__2725 (
            .O(N__13037),
            .I(rUartRxStateZ0Z_0));
    LocalMux I__2724 (
            .O(N__13034),
            .I(rUartRxStateZ0Z_0));
    LocalMux I__2723 (
            .O(N__13031),
            .I(rUartRxStateZ0Z_0));
    LocalMux I__2722 (
            .O(N__13028),
            .I(rUartRxStateZ0Z_0));
    InMux I__2721 (
            .O(N__13019),
            .I(N__13016));
    LocalMux I__2720 (
            .O(N__13016),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rDataCount_c2 ));
    InMux I__2719 (
            .O(N__13013),
            .I(N__13007));
    InMux I__2718 (
            .O(N__13012),
            .I(N__13007));
    LocalMux I__2717 (
            .O(N__13007),
            .I(\uart_inst0.rx_uart_fifo_inst.rDataCount_0_sqmuxa ));
    CascadeMux I__2716 (
            .O(N__13004),
            .I(N__12997));
    CascadeMux I__2715 (
            .O(N__13003),
            .I(N__12994));
    InMux I__2714 (
            .O(N__13002),
            .I(N__12991));
    InMux I__2713 (
            .O(N__13001),
            .I(N__12986));
    InMux I__2712 (
            .O(N__13000),
            .I(N__12986));
    InMux I__2711 (
            .O(N__12997),
            .I(N__12981));
    InMux I__2710 (
            .O(N__12994),
            .I(N__12981));
    LocalMux I__2709 (
            .O(N__12991),
            .I(\uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_2 ));
    LocalMux I__2708 (
            .O(N__12986),
            .I(\uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_2 ));
    LocalMux I__2707 (
            .O(N__12981),
            .I(\uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_2 ));
    InMux I__2706 (
            .O(N__12974),
            .I(N__12971));
    LocalMux I__2705 (
            .O(N__12971),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rDataCount_axbxc3_1_1 ));
    CascadeMux I__2704 (
            .O(N__12968),
            .I(N__12963));
    CascadeMux I__2703 (
            .O(N__12967),
            .I(N__12959));
    InMux I__2702 (
            .O(N__12966),
            .I(N__12954));
    InMux I__2701 (
            .O(N__12963),
            .I(N__12949));
    InMux I__2700 (
            .O(N__12962),
            .I(N__12949));
    InMux I__2699 (
            .O(N__12959),
            .I(N__12942));
    InMux I__2698 (
            .O(N__12958),
            .I(N__12942));
    InMux I__2697 (
            .O(N__12957),
            .I(N__12942));
    LocalMux I__2696 (
            .O(N__12954),
            .I(\uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_1 ));
    LocalMux I__2695 (
            .O(N__12949),
            .I(\uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_1 ));
    LocalMux I__2694 (
            .O(N__12942),
            .I(\uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_1 ));
    CascadeMux I__2693 (
            .O(N__12935),
            .I(N__12931));
    InMux I__2692 (
            .O(N__12934),
            .I(N__12922));
    InMux I__2691 (
            .O(N__12931),
            .I(N__12922));
    InMux I__2690 (
            .O(N__12930),
            .I(N__12917));
    InMux I__2689 (
            .O(N__12929),
            .I(N__12917));
    InMux I__2688 (
            .O(N__12928),
            .I(N__12912));
    InMux I__2687 (
            .O(N__12927),
            .I(N__12912));
    LocalMux I__2686 (
            .O(N__12922),
            .I(\uart_inst0.wRxWrFull_0 ));
    LocalMux I__2685 (
            .O(N__12917),
            .I(\uart_inst0.wRxWrFull_0 ));
    LocalMux I__2684 (
            .O(N__12912),
            .I(\uart_inst0.wRxWrFull_0 ));
    InMux I__2683 (
            .O(N__12905),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_5 ));
    InMux I__2682 (
            .O(N__12902),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_6 ));
    InMux I__2681 (
            .O(N__12899),
            .I(bfn_17_7_0_));
    InMux I__2680 (
            .O(N__12896),
            .I(N__12893));
    LocalMux I__2679 (
            .O(N__12893),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNO_0_0_3 ));
    InMux I__2678 (
            .O(N__12890),
            .I(N__12887));
    LocalMux I__2677 (
            .O(N__12887),
            .I(\uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNO_0_0_0 ));
    CascadeMux I__2676 (
            .O(N__12884),
            .I(wUartRxEmpty_cascade_));
    InMux I__2675 (
            .O(N__12881),
            .I(N__12878));
    LocalMux I__2674 (
            .O(N__12878),
            .I(N__12875));
    Odrv4 I__2673 (
            .O(N__12875),
            .I(rRxDataZ0Z_0));
    InMux I__2672 (
            .O(N__12872),
            .I(N__12869));
    LocalMux I__2671 (
            .O(N__12869),
            .I(N__12866));
    Span4Mux_h I__2670 (
            .O(N__12866),
            .I(N__12863));
    Odrv4 I__2669 (
            .O(N__12863),
            .I(rRxDataZ0Z_5));
    InMux I__2668 (
            .O(N__12860),
            .I(N__12857));
    LocalMux I__2667 (
            .O(N__12857),
            .I(N__12854));
    Odrv4 I__2666 (
            .O(N__12854),
            .I(rRxDataZ0Z_7));
    CEMux I__2665 (
            .O(N__12851),
            .I(N__12847));
    CEMux I__2664 (
            .O(N__12850),
            .I(N__12844));
    LocalMux I__2663 (
            .O(N__12847),
            .I(N__12841));
    LocalMux I__2662 (
            .O(N__12844),
            .I(N__12838));
    Span4Mux_h I__2661 (
            .O(N__12841),
            .I(N__12835));
    Span4Mux_h I__2660 (
            .O(N__12838),
            .I(N__12832));
    Odrv4 I__2659 (
            .O(N__12835),
            .I(N_27_0));
    Odrv4 I__2658 (
            .O(N__12832),
            .I(N_27_0));
    InMux I__2657 (
            .O(N__12827),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_0 ));
    InMux I__2656 (
            .O(N__12824),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_1 ));
    InMux I__2655 (
            .O(N__12821),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_2 ));
    InMux I__2654 (
            .O(N__12818),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_3 ));
    InMux I__2653 (
            .O(N__12815),
            .I(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_4 ));
    InMux I__2652 (
            .O(N__12812),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_5 ));
    InMux I__2651 (
            .O(N__12809),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_6 ));
    InMux I__2650 (
            .O(N__12806),
            .I(bfn_17_3_0_));
    CascadeMux I__2649 (
            .O(N__12803),
            .I(N__12800));
    InMux I__2648 (
            .O(N__12800),
            .I(N__12797));
    LocalMux I__2647 (
            .O(N__12797),
            .I(N__12793));
    InMux I__2646 (
            .O(N__12796),
            .I(N__12790));
    Span4Mux_s2_v I__2645 (
            .O(N__12793),
            .I(N__12787));
    LocalMux I__2644 (
            .O(N__12790),
            .I(N__12784));
    Odrv4 I__2643 (
            .O(N__12787),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIGAUPZ0 ));
    Odrv4 I__2642 (
            .O(N__12784),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIGAUPZ0 ));
    InMux I__2641 (
            .O(N__12779),
            .I(N__12776));
    LocalMux I__2640 (
            .O(N__12776),
            .I(N__12772));
    InMux I__2639 (
            .O(N__12775),
            .I(N__12769));
    Odrv4 I__2638 (
            .O(N__12772),
            .I(fifo_inst_tx_fifo_inst_rRamRdAddr_2));
    LocalMux I__2637 (
            .O(N__12769),
            .I(fifo_inst_tx_fifo_inst_rRamRdAddr_2));
    InMux I__2636 (
            .O(N__12764),
            .I(N__12759));
    InMux I__2635 (
            .O(N__12763),
            .I(N__12751));
    InMux I__2634 (
            .O(N__12762),
            .I(N__12746));
    LocalMux I__2633 (
            .O(N__12759),
            .I(N__12743));
    InMux I__2632 (
            .O(N__12758),
            .I(N__12732));
    InMux I__2631 (
            .O(N__12757),
            .I(N__12732));
    InMux I__2630 (
            .O(N__12756),
            .I(N__12732));
    InMux I__2629 (
            .O(N__12755),
            .I(N__12732));
    InMux I__2628 (
            .O(N__12754),
            .I(N__12732));
    LocalMux I__2627 (
            .O(N__12751),
            .I(N__12729));
    InMux I__2626 (
            .O(N__12750),
            .I(N__12726));
    InMux I__2625 (
            .O(N__12749),
            .I(N__12722));
    LocalMux I__2624 (
            .O(N__12746),
            .I(N__12719));
    Span4Mux_h I__2623 (
            .O(N__12743),
            .I(N__12712));
    LocalMux I__2622 (
            .O(N__12732),
            .I(N__12712));
    Span4Mux_v I__2621 (
            .O(N__12729),
            .I(N__12712));
    LocalMux I__2620 (
            .O(N__12726),
            .I(N__12709));
    InMux I__2619 (
            .O(N__12725),
            .I(N__12706));
    LocalMux I__2618 (
            .O(N__12722),
            .I(fifo_inst_wRxWrFull));
    Odrv12 I__2617 (
            .O(N__12719),
            .I(fifo_inst_wRxWrFull));
    Odrv4 I__2616 (
            .O(N__12712),
            .I(fifo_inst_wRxWrFull));
    Odrv4 I__2615 (
            .O(N__12709),
            .I(fifo_inst_wRxWrFull));
    LocalMux I__2614 (
            .O(N__12706),
            .I(fifo_inst_wRxWrFull));
    InMux I__2613 (
            .O(N__12695),
            .I(N__12692));
    LocalMux I__2612 (
            .O(N__12692),
            .I(N__12683));
    InMux I__2611 (
            .O(N__12691),
            .I(N__12680));
    InMux I__2610 (
            .O(N__12690),
            .I(N__12675));
    InMux I__2609 (
            .O(N__12689),
            .I(N__12675));
    InMux I__2608 (
            .O(N__12688),
            .I(N__12668));
    InMux I__2607 (
            .O(N__12687),
            .I(N__12668));
    InMux I__2606 (
            .O(N__12686),
            .I(N__12668));
    Span4Mux_h I__2605 (
            .O(N__12683),
            .I(N__12665));
    LocalMux I__2604 (
            .O(N__12680),
            .I(fifo_inst_rx_fifo_inst_rDataCount_2));
    LocalMux I__2603 (
            .O(N__12675),
            .I(fifo_inst_rx_fifo_inst_rDataCount_2));
    LocalMux I__2602 (
            .O(N__12668),
            .I(fifo_inst_rx_fifo_inst_rDataCount_2));
    Odrv4 I__2601 (
            .O(N__12665),
            .I(fifo_inst_rx_fifo_inst_rDataCount_2));
    CascadeMux I__2600 (
            .O(N__12656),
            .I(N__12653));
    InMux I__2599 (
            .O(N__12653),
            .I(N__12647));
    CascadeMux I__2598 (
            .O(N__12652),
            .I(N__12642));
    CascadeMux I__2597 (
            .O(N__12651),
            .I(N__12638));
    CascadeMux I__2596 (
            .O(N__12650),
            .I(N__12634));
    LocalMux I__2595 (
            .O(N__12647),
            .I(N__12631));
    InMux I__2594 (
            .O(N__12646),
            .I(N__12628));
    InMux I__2593 (
            .O(N__12645),
            .I(N__12625));
    InMux I__2592 (
            .O(N__12642),
            .I(N__12618));
    InMux I__2591 (
            .O(N__12641),
            .I(N__12618));
    InMux I__2590 (
            .O(N__12638),
            .I(N__12618));
    InMux I__2589 (
            .O(N__12637),
            .I(N__12613));
    InMux I__2588 (
            .O(N__12634),
            .I(N__12613));
    Span4Mux_h I__2587 (
            .O(N__12631),
            .I(N__12610));
    LocalMux I__2586 (
            .O(N__12628),
            .I(fifo_inst_rx_fifo_inst_rDataCount_0));
    LocalMux I__2585 (
            .O(N__12625),
            .I(fifo_inst_rx_fifo_inst_rDataCount_0));
    LocalMux I__2584 (
            .O(N__12618),
            .I(fifo_inst_rx_fifo_inst_rDataCount_0));
    LocalMux I__2583 (
            .O(N__12613),
            .I(fifo_inst_rx_fifo_inst_rDataCount_0));
    Odrv4 I__2582 (
            .O(N__12610),
            .I(fifo_inst_rx_fifo_inst_rDataCount_0));
    InMux I__2581 (
            .O(N__12599),
            .I(N__12595));
    CascadeMux I__2580 (
            .O(N__12598),
            .I(N__12589));
    LocalMux I__2579 (
            .O(N__12595),
            .I(N__12583));
    InMux I__2578 (
            .O(N__12594),
            .I(N__12580));
    InMux I__2577 (
            .O(N__12593),
            .I(N__12577));
    InMux I__2576 (
            .O(N__12592),
            .I(N__12574));
    InMux I__2575 (
            .O(N__12589),
            .I(N__12567));
    InMux I__2574 (
            .O(N__12588),
            .I(N__12567));
    InMux I__2573 (
            .O(N__12587),
            .I(N__12567));
    InMux I__2572 (
            .O(N__12586),
            .I(N__12564));
    Span4Mux_v I__2571 (
            .O(N__12583),
            .I(N__12561));
    LocalMux I__2570 (
            .O(N__12580),
            .I(fifo_inst_rx_fifo_inst_rDataCount_1));
    LocalMux I__2569 (
            .O(N__12577),
            .I(fifo_inst_rx_fifo_inst_rDataCount_1));
    LocalMux I__2568 (
            .O(N__12574),
            .I(fifo_inst_rx_fifo_inst_rDataCount_1));
    LocalMux I__2567 (
            .O(N__12567),
            .I(fifo_inst_rx_fifo_inst_rDataCount_1));
    LocalMux I__2566 (
            .O(N__12564),
            .I(fifo_inst_rx_fifo_inst_rDataCount_1));
    Odrv4 I__2565 (
            .O(N__12561),
            .I(fifo_inst_rx_fifo_inst_rDataCount_1));
    InMux I__2564 (
            .O(N__12548),
            .I(N__12545));
    LocalMux I__2563 (
            .O(N__12545),
            .I(N__12542));
    Span4Mux_h I__2562 (
            .O(N__12542),
            .I(N__12539));
    Odrv4 I__2561 (
            .O(N__12539),
            .I(rRxDataZ0Z_6));
    InMux I__2560 (
            .O(N__12536),
            .I(N__12533));
    LocalMux I__2559 (
            .O(N__12533),
            .I(N__12530));
    Span4Mux_h I__2558 (
            .O(N__12530),
            .I(N__12527));
    Odrv4 I__2557 (
            .O(N__12527),
            .I(rRxDataZ0Z_1));
    CascadeMux I__2556 (
            .O(N__12524),
            .I(N__12521));
    InMux I__2555 (
            .O(N__12521),
            .I(N__12518));
    LocalMux I__2554 (
            .O(N__12518),
            .I(N__12515));
    Odrv4 I__2553 (
            .O(N__12515),
            .I(rRxDataZ0Z_2));
    InMux I__2552 (
            .O(N__12512),
            .I(N__12509));
    LocalMux I__2551 (
            .O(N__12509),
            .I(N__12506));
    Odrv4 I__2550 (
            .O(N__12506),
            .I(rRxDataZ0Z_3));
    InMux I__2549 (
            .O(N__12503),
            .I(N__12498));
    InMux I__2548 (
            .O(N__12502),
            .I(N__12495));
    InMux I__2547 (
            .O(N__12501),
            .I(N__12492));
    LocalMux I__2546 (
            .O(N__12498),
            .I(N__12487));
    LocalMux I__2545 (
            .O(N__12495),
            .I(N__12487));
    LocalMux I__2544 (
            .O(N__12492),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_12 ));
    Odrv4 I__2543 (
            .O(N__12487),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_12 ));
    InMux I__2542 (
            .O(N__12482),
            .I(N__12479));
    LocalMux I__2541 (
            .O(N__12479),
            .I(N__12476));
    Odrv4 I__2540 (
            .O(N__12476),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_11_s1_THRU_CO ));
    InMux I__2539 (
            .O(N__12473),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_11_s1 ));
    IoInMux I__2538 (
            .O(N__12470),
            .I(N__12467));
    LocalMux I__2537 (
            .O(N__12467),
            .I(N__12464));
    IoSpan4Mux I__2536 (
            .O(N__12464),
            .I(N__12461));
    Span4Mux_s2_v I__2535 (
            .O(N__12461),
            .I(N__12446));
    CascadeMux I__2534 (
            .O(N__12460),
            .I(N__12443));
    CascadeMux I__2533 (
            .O(N__12459),
            .I(N__12440));
    CascadeMux I__2532 (
            .O(N__12458),
            .I(N__12436));
    CascadeMux I__2531 (
            .O(N__12457),
            .I(N__12433));
    CascadeMux I__2530 (
            .O(N__12456),
            .I(N__12430));
    CascadeMux I__2529 (
            .O(N__12455),
            .I(N__12427));
    CascadeMux I__2528 (
            .O(N__12454),
            .I(N__12424));
    CascadeMux I__2527 (
            .O(N__12453),
            .I(N__12421));
    CascadeMux I__2526 (
            .O(N__12452),
            .I(N__12418));
    CascadeMux I__2525 (
            .O(N__12451),
            .I(N__12415));
    CascadeMux I__2524 (
            .O(N__12450),
            .I(N__12412));
    CascadeMux I__2523 (
            .O(N__12449),
            .I(N__12409));
    Span4Mux_v I__2522 (
            .O(N__12446),
            .I(N__12399));
    InMux I__2521 (
            .O(N__12443),
            .I(N__12390));
    InMux I__2520 (
            .O(N__12440),
            .I(N__12390));
    InMux I__2519 (
            .O(N__12439),
            .I(N__12390));
    InMux I__2518 (
            .O(N__12436),
            .I(N__12390));
    InMux I__2517 (
            .O(N__12433),
            .I(N__12385));
    InMux I__2516 (
            .O(N__12430),
            .I(N__12385));
    InMux I__2515 (
            .O(N__12427),
            .I(N__12378));
    InMux I__2514 (
            .O(N__12424),
            .I(N__12378));
    InMux I__2513 (
            .O(N__12421),
            .I(N__12378));
    InMux I__2512 (
            .O(N__12418),
            .I(N__12369));
    InMux I__2511 (
            .O(N__12415),
            .I(N__12369));
    InMux I__2510 (
            .O(N__12412),
            .I(N__12369));
    InMux I__2509 (
            .O(N__12409),
            .I(N__12369));
    CascadeMux I__2508 (
            .O(N__12408),
            .I(N__12366));
    CascadeMux I__2507 (
            .O(N__12407),
            .I(N__12363));
    CascadeMux I__2506 (
            .O(N__12406),
            .I(N__12360));
    CascadeMux I__2505 (
            .O(N__12405),
            .I(N__12357));
    CascadeMux I__2504 (
            .O(N__12404),
            .I(N__12353));
    CascadeMux I__2503 (
            .O(N__12403),
            .I(N__12349));
    CascadeMux I__2502 (
            .O(N__12402),
            .I(N__12345));
    Span4Mux_v I__2501 (
            .O(N__12399),
            .I(N__12327));
    LocalMux I__2500 (
            .O(N__12390),
            .I(N__12327));
    LocalMux I__2499 (
            .O(N__12385),
            .I(N__12327));
    LocalMux I__2498 (
            .O(N__12378),
            .I(N__12327));
    LocalMux I__2497 (
            .O(N__12369),
            .I(N__12327));
    InMux I__2496 (
            .O(N__12366),
            .I(N__12322));
    InMux I__2495 (
            .O(N__12363),
            .I(N__12322));
    InMux I__2494 (
            .O(N__12360),
            .I(N__12317));
    InMux I__2493 (
            .O(N__12357),
            .I(N__12317));
    InMux I__2492 (
            .O(N__12356),
            .I(N__12300));
    InMux I__2491 (
            .O(N__12353),
            .I(N__12300));
    InMux I__2490 (
            .O(N__12352),
            .I(N__12300));
    InMux I__2489 (
            .O(N__12349),
            .I(N__12300));
    InMux I__2488 (
            .O(N__12348),
            .I(N__12300));
    InMux I__2487 (
            .O(N__12345),
            .I(N__12300));
    CascadeMux I__2486 (
            .O(N__12344),
            .I(N__12297));
    CascadeMux I__2485 (
            .O(N__12343),
            .I(N__12294));
    CascadeMux I__2484 (
            .O(N__12342),
            .I(N__12291));
    CascadeMux I__2483 (
            .O(N__12341),
            .I(N__12288));
    CascadeMux I__2482 (
            .O(N__12340),
            .I(N__12285));
    CascadeMux I__2481 (
            .O(N__12339),
            .I(N__12282));
    CascadeMux I__2480 (
            .O(N__12338),
            .I(N__12279));
    Span4Mux_v I__2479 (
            .O(N__12327),
            .I(N__12271));
    LocalMux I__2478 (
            .O(N__12322),
            .I(N__12271));
    LocalMux I__2477 (
            .O(N__12317),
            .I(N__12271));
    SRMux I__2476 (
            .O(N__12316),
            .I(N__12268));
    SRMux I__2475 (
            .O(N__12315),
            .I(N__12264));
    SRMux I__2474 (
            .O(N__12314),
            .I(N__12261));
    SRMux I__2473 (
            .O(N__12313),
            .I(N__12258));
    LocalMux I__2472 (
            .O(N__12300),
            .I(N__12253));
    InMux I__2471 (
            .O(N__12297),
            .I(N__12246));
    InMux I__2470 (
            .O(N__12294),
            .I(N__12246));
    InMux I__2469 (
            .O(N__12291),
            .I(N__12246));
    InMux I__2468 (
            .O(N__12288),
            .I(N__12237));
    InMux I__2467 (
            .O(N__12285),
            .I(N__12237));
    InMux I__2466 (
            .O(N__12282),
            .I(N__12237));
    InMux I__2465 (
            .O(N__12279),
            .I(N__12237));
    SRMux I__2464 (
            .O(N__12278),
            .I(N__12234));
    Span4Mux_v I__2463 (
            .O(N__12271),
            .I(N__12229));
    LocalMux I__2462 (
            .O(N__12268),
            .I(N__12229));
    SRMux I__2461 (
            .O(N__12267),
            .I(N__12226));
    LocalMux I__2460 (
            .O(N__12264),
            .I(N__12223));
    LocalMux I__2459 (
            .O(N__12261),
            .I(N__12218));
    LocalMux I__2458 (
            .O(N__12258),
            .I(N__12218));
    SRMux I__2457 (
            .O(N__12257),
            .I(N__12215));
    SRMux I__2456 (
            .O(N__12256),
            .I(N__12212));
    Span4Mux_v I__2455 (
            .O(N__12253),
            .I(N__12205));
    LocalMux I__2454 (
            .O(N__12246),
            .I(N__12205));
    LocalMux I__2453 (
            .O(N__12237),
            .I(N__12205));
    LocalMux I__2452 (
            .O(N__12234),
            .I(N__12202));
    Span4Mux_h I__2451 (
            .O(N__12229),
            .I(N__12197));
    LocalMux I__2450 (
            .O(N__12226),
            .I(N__12197));
    Span4Mux_s3_v I__2449 (
            .O(N__12223),
            .I(N__12192));
    Span4Mux_s3_v I__2448 (
            .O(N__12218),
            .I(N__12192));
    LocalMux I__2447 (
            .O(N__12215),
            .I(N__12189));
    LocalMux I__2446 (
            .O(N__12212),
            .I(N__12186));
    Span4Mux_h I__2445 (
            .O(N__12205),
            .I(N__12183));
    Span4Mux_h I__2444 (
            .O(N__12202),
            .I(N__12180));
    Span4Mux_v I__2443 (
            .O(N__12197),
            .I(N__12177));
    Span4Mux_v I__2442 (
            .O(N__12192),
            .I(N__12172));
    Span4Mux_v I__2441 (
            .O(N__12189),
            .I(N__12172));
    Span12Mux_h I__2440 (
            .O(N__12186),
            .I(N__12169));
    Span4Mux_v I__2439 (
            .O(N__12183),
            .I(N__12166));
    Span4Mux_h I__2438 (
            .O(N__12180),
            .I(N__12163));
    Span4Mux_h I__2437 (
            .O(N__12177),
            .I(N__12158));
    Span4Mux_h I__2436 (
            .O(N__12172),
            .I(N__12158));
    Odrv12 I__2435 (
            .O(N__12169),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2434 (
            .O(N__12166),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2433 (
            .O(N__12163),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__2432 (
            .O(N__12158),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__2431 (
            .O(N__12149),
            .I(N__12145));
    CascadeMux I__2430 (
            .O(N__12148),
            .I(N__12141));
    InMux I__2429 (
            .O(N__12145),
            .I(N__12138));
    InMux I__2428 (
            .O(N__12144),
            .I(N__12133));
    InMux I__2427 (
            .O(N__12141),
            .I(N__12133));
    LocalMux I__2426 (
            .O(N__12138),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_13 ));
    LocalMux I__2425 (
            .O(N__12133),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_13 ));
    InMux I__2424 (
            .O(N__12128),
            .I(N__12125));
    LocalMux I__2423 (
            .O(N__12125),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_12_s1_THRU_CO ));
    InMux I__2422 (
            .O(N__12122),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_12_s1 ));
    InMux I__2421 (
            .O(N__12119),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_13_s1 ));
    InMux I__2420 (
            .O(N__12116),
            .I(N__12112));
    InMux I__2419 (
            .O(N__12115),
            .I(N__12109));
    LocalMux I__2418 (
            .O(N__12112),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_14 ));
    LocalMux I__2417 (
            .O(N__12109),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_14 ));
    CEMux I__2416 (
            .O(N__12104),
            .I(N__12101));
    LocalMux I__2415 (
            .O(N__12101),
            .I(N__12098));
    Span4Mux_h I__2414 (
            .O(N__12098),
            .I(N__12095));
    Odrv4 I__2413 (
            .O(N__12095),
            .I(\uart_inst0.uart_inst0.N_147_0_i_0 ));
    InMux I__2412 (
            .O(N__12092),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_0 ));
    InMux I__2411 (
            .O(N__12089),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_1 ));
    InMux I__2410 (
            .O(N__12086),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_2 ));
    InMux I__2409 (
            .O(N__12083),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_3 ));
    InMux I__2408 (
            .O(N__12080),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_4 ));
    CascadeMux I__2407 (
            .O(N__12077),
            .I(N__12072));
    InMux I__2406 (
            .O(N__12076),
            .I(N__12069));
    InMux I__2405 (
            .O(N__12075),
            .I(N__12066));
    InMux I__2404 (
            .O(N__12072),
            .I(N__12063));
    LocalMux I__2403 (
            .O(N__12069),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_5 ));
    LocalMux I__2402 (
            .O(N__12066),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_5 ));
    LocalMux I__2401 (
            .O(N__12063),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_5 ));
    InMux I__2400 (
            .O(N__12056),
            .I(N__12053));
    LocalMux I__2399 (
            .O(N__12053),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_4_s1_THRU_CO ));
    InMux I__2398 (
            .O(N__12050),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_4_s1 ));
    InMux I__2397 (
            .O(N__12047),
            .I(N__12042));
    InMux I__2396 (
            .O(N__12046),
            .I(N__12039));
    InMux I__2395 (
            .O(N__12045),
            .I(N__12036));
    LocalMux I__2394 (
            .O(N__12042),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_6 ));
    LocalMux I__2393 (
            .O(N__12039),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_6 ));
    LocalMux I__2392 (
            .O(N__12036),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_6 ));
    InMux I__2391 (
            .O(N__12029),
            .I(N__12026));
    LocalMux I__2390 (
            .O(N__12026),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_5_s1_THRU_CO ));
    InMux I__2389 (
            .O(N__12023),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_5_s1 ));
    InMux I__2388 (
            .O(N__12020),
            .I(N__12015));
    InMux I__2387 (
            .O(N__12019),
            .I(N__12012));
    InMux I__2386 (
            .O(N__12018),
            .I(N__12009));
    LocalMux I__2385 (
            .O(N__12015),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_7 ));
    LocalMux I__2384 (
            .O(N__12012),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_7 ));
    LocalMux I__2383 (
            .O(N__12009),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_7 ));
    InMux I__2382 (
            .O(N__12002),
            .I(N__11999));
    LocalMux I__2381 (
            .O(N__11999),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_6_s1_THRU_CO ));
    InMux I__2380 (
            .O(N__11996),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_6_s1 ));
    InMux I__2379 (
            .O(N__11993),
            .I(N__11989));
    InMux I__2378 (
            .O(N__11992),
            .I(N__11985));
    LocalMux I__2377 (
            .O(N__11989),
            .I(N__11982));
    InMux I__2376 (
            .O(N__11988),
            .I(N__11979));
    LocalMux I__2375 (
            .O(N__11985),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_8 ));
    Odrv4 I__2374 (
            .O(N__11982),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_8 ));
    LocalMux I__2373 (
            .O(N__11979),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_8 ));
    InMux I__2372 (
            .O(N__11972),
            .I(N__11969));
    LocalMux I__2371 (
            .O(N__11969),
            .I(N__11966));
    Odrv4 I__2370 (
            .O(N__11966),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_7_s1_THRU_CO ));
    InMux I__2369 (
            .O(N__11963),
            .I(bfn_16_19_0_));
    InMux I__2368 (
            .O(N__11960),
            .I(N__11956));
    InMux I__2367 (
            .O(N__11959),
            .I(N__11952));
    LocalMux I__2366 (
            .O(N__11956),
            .I(N__11949));
    InMux I__2365 (
            .O(N__11955),
            .I(N__11946));
    LocalMux I__2364 (
            .O(N__11952),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_9 ));
    Odrv4 I__2363 (
            .O(N__11949),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_9 ));
    LocalMux I__2362 (
            .O(N__11946),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_9 ));
    InMux I__2361 (
            .O(N__11939),
            .I(N__11936));
    LocalMux I__2360 (
            .O(N__11936),
            .I(N__11933));
    Odrv4 I__2359 (
            .O(N__11933),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_8_s1_THRU_CO ));
    InMux I__2358 (
            .O(N__11930),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_8_s1 ));
    InMux I__2357 (
            .O(N__11927),
            .I(N__11922));
    InMux I__2356 (
            .O(N__11926),
            .I(N__11917));
    InMux I__2355 (
            .O(N__11925),
            .I(N__11917));
    LocalMux I__2354 (
            .O(N__11922),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_10 ));
    LocalMux I__2353 (
            .O(N__11917),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_10 ));
    InMux I__2352 (
            .O(N__11912),
            .I(N__11909));
    LocalMux I__2351 (
            .O(N__11909),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_9_s1_THRU_CO ));
    InMux I__2350 (
            .O(N__11906),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_9_s1 ));
    InMux I__2349 (
            .O(N__11903),
            .I(N__11898));
    InMux I__2348 (
            .O(N__11902),
            .I(N__11893));
    InMux I__2347 (
            .O(N__11901),
            .I(N__11893));
    LocalMux I__2346 (
            .O(N__11898),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_11 ));
    LocalMux I__2345 (
            .O(N__11893),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_11 ));
    InMux I__2344 (
            .O(N__11888),
            .I(N__11885));
    LocalMux I__2343 (
            .O(N__11885),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_10_s1_THRU_CO ));
    InMux I__2342 (
            .O(N__11882),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_10_s1 ));
    CascadeMux I__2341 (
            .O(N__11879),
            .I(N__11876));
    InMux I__2340 (
            .O(N__11876),
            .I(N__11868));
    InMux I__2339 (
            .O(N__11875),
            .I(N__11868));
    InMux I__2338 (
            .O(N__11874),
            .I(N__11865));
    InMux I__2337 (
            .O(N__11873),
            .I(N__11862));
    LocalMux I__2336 (
            .O(N__11868),
            .I(N__11850));
    LocalMux I__2335 (
            .O(N__11865),
            .I(N__11845));
    LocalMux I__2334 (
            .O(N__11862),
            .I(N__11845));
    InMux I__2333 (
            .O(N__11861),
            .I(N__11840));
    InMux I__2332 (
            .O(N__11860),
            .I(N__11840));
    InMux I__2331 (
            .O(N__11859),
            .I(N__11831));
    InMux I__2330 (
            .O(N__11858),
            .I(N__11831));
    InMux I__2329 (
            .O(N__11857),
            .I(N__11831));
    InMux I__2328 (
            .O(N__11856),
            .I(N__11831));
    InMux I__2327 (
            .O(N__11855),
            .I(N__11824));
    InMux I__2326 (
            .O(N__11854),
            .I(N__11824));
    InMux I__2325 (
            .O(N__11853),
            .I(N__11824));
    Odrv4 I__2324 (
            .O(N__11850),
            .I(\uart_inst0.uart_inst0.N_147_0 ));
    Odrv4 I__2323 (
            .O(N__11845),
            .I(\uart_inst0.uart_inst0.N_147_0 ));
    LocalMux I__2322 (
            .O(N__11840),
            .I(\uart_inst0.uart_inst0.N_147_0 ));
    LocalMux I__2321 (
            .O(N__11831),
            .I(\uart_inst0.uart_inst0.N_147_0 ));
    LocalMux I__2320 (
            .O(N__11824),
            .I(\uart_inst0.uart_inst0.N_147_0 ));
    CascadeMux I__2319 (
            .O(N__11813),
            .I(N__11810));
    InMux I__2318 (
            .O(N__11810),
            .I(N__11807));
    LocalMux I__2317 (
            .O(N__11807),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_0_s1_THRU_CO ));
    InMux I__2316 (
            .O(N__11804),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_0_s1 ));
    InMux I__2315 (
            .O(N__11801),
            .I(N__11798));
    LocalMux I__2314 (
            .O(N__11798),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_1_s1_THRU_CO ));
    InMux I__2313 (
            .O(N__11795),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_1_s1 ));
    InMux I__2312 (
            .O(N__11792),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_2_s1 ));
    InMux I__2311 (
            .O(N__11789),
            .I(N__11784));
    InMux I__2310 (
            .O(N__11788),
            .I(N__11781));
    InMux I__2309 (
            .O(N__11787),
            .I(N__11778));
    LocalMux I__2308 (
            .O(N__11784),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_4 ));
    LocalMux I__2307 (
            .O(N__11781),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_4 ));
    LocalMux I__2306 (
            .O(N__11778),
            .I(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_4 ));
    InMux I__2305 (
            .O(N__11771),
            .I(N__11768));
    LocalMux I__2304 (
            .O(N__11768),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_3_s1_THRU_CO ));
    InMux I__2303 (
            .O(N__11765),
            .I(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_3_s1 ));
    InMux I__2302 (
            .O(N__11762),
            .I(N__11759));
    LocalMux I__2301 (
            .O(N__11759),
            .I(\uart_inst0.uart_inst0.rx_countdown_cry_3_THRU_CO ));
    InMux I__2300 (
            .O(N__11756),
            .I(\uart_inst0.uart_inst0.rx_countdown_cry_3 ));
    InMux I__2299 (
            .O(N__11753),
            .I(N__11745));
    InMux I__2298 (
            .O(N__11752),
            .I(N__11734));
    InMux I__2297 (
            .O(N__11751),
            .I(N__11734));
    InMux I__2296 (
            .O(N__11750),
            .I(N__11734));
    InMux I__2295 (
            .O(N__11749),
            .I(N__11734));
    InMux I__2294 (
            .O(N__11748),
            .I(N__11734));
    LocalMux I__2293 (
            .O(N__11745),
            .I(\uart_inst0.uart_inst0.N_252_0_i ));
    LocalMux I__2292 (
            .O(N__11734),
            .I(\uart_inst0.uart_inst0.N_252_0_i ));
    InMux I__2291 (
            .O(N__11729),
            .I(\uart_inst0.uart_inst0.rx_countdown_cry_4 ));
    CascadeMux I__2290 (
            .O(N__11726),
            .I(N__11722));
    InMux I__2289 (
            .O(N__11725),
            .I(N__11719));
    InMux I__2288 (
            .O(N__11722),
            .I(N__11716));
    LocalMux I__2287 (
            .O(N__11719),
            .I(\uart_inst0.uart_inst0.rx_countdownZ0Z_5 ));
    LocalMux I__2286 (
            .O(N__11716),
            .I(\uart_inst0.uart_inst0.rx_countdownZ0Z_5 ));
    CEMux I__2285 (
            .O(N__11711),
            .I(N__11707));
    CEMux I__2284 (
            .O(N__11710),
            .I(N__11704));
    LocalMux I__2283 (
            .O(N__11707),
            .I(N__11701));
    LocalMux I__2282 (
            .O(N__11704),
            .I(N__11698));
    Odrv4 I__2281 (
            .O(N__11701),
            .I(\uart_inst0.uart_inst0.rx_countdowne_0_i ));
    Odrv4 I__2280 (
            .O(N__11698),
            .I(\uart_inst0.uart_inst0.rx_countdowne_0_i ));
    InMux I__2279 (
            .O(N__11693),
            .I(N__11688));
    InMux I__2278 (
            .O(N__11692),
            .I(N__11685));
    InMux I__2277 (
            .O(N__11691),
            .I(N__11682));
    LocalMux I__2276 (
            .O(N__11688),
            .I(N__11675));
    LocalMux I__2275 (
            .O(N__11685),
            .I(N__11675));
    LocalMux I__2274 (
            .O(N__11682),
            .I(N__11675));
    Odrv4 I__2273 (
            .O(N__11675),
            .I(\uart_inst0.uart_inst0.N_258_0 ));
    CascadeMux I__2272 (
            .O(N__11672),
            .I(\uart_inst0.uart_inst0.N_276_cascade_ ));
    InMux I__2271 (
            .O(N__11669),
            .I(N__11666));
    LocalMux I__2270 (
            .O(N__11666),
            .I(N__11662));
    InMux I__2269 (
            .O(N__11665),
            .I(N__11655));
    Span4Mux_h I__2268 (
            .O(N__11662),
            .I(N__11645));
    InMux I__2267 (
            .O(N__11661),
            .I(N__11640));
    InMux I__2266 (
            .O(N__11660),
            .I(N__11640));
    InMux I__2265 (
            .O(N__11659),
            .I(N__11637));
    InMux I__2264 (
            .O(N__11658),
            .I(N__11634));
    LocalMux I__2263 (
            .O(N__11655),
            .I(N__11631));
    InMux I__2262 (
            .O(N__11654),
            .I(N__11628));
    InMux I__2261 (
            .O(N__11653),
            .I(N__11625));
    InMux I__2260 (
            .O(N__11652),
            .I(N__11620));
    InMux I__2259 (
            .O(N__11651),
            .I(N__11620));
    InMux I__2258 (
            .O(N__11650),
            .I(N__11613));
    InMux I__2257 (
            .O(N__11649),
            .I(N__11613));
    InMux I__2256 (
            .O(N__11648),
            .I(N__11613));
    Span4Mux_v I__2255 (
            .O(N__11645),
            .I(N__11606));
    LocalMux I__2254 (
            .O(N__11640),
            .I(N__11606));
    LocalMux I__2253 (
            .O(N__11637),
            .I(N__11606));
    LocalMux I__2252 (
            .O(N__11634),
            .I(\uart_inst0.uart_inst0.tx_stateZ0Z_0 ));
    Odrv4 I__2251 (
            .O(N__11631),
            .I(\uart_inst0.uart_inst0.tx_stateZ0Z_0 ));
    LocalMux I__2250 (
            .O(N__11628),
            .I(\uart_inst0.uart_inst0.tx_stateZ0Z_0 ));
    LocalMux I__2249 (
            .O(N__11625),
            .I(\uart_inst0.uart_inst0.tx_stateZ0Z_0 ));
    LocalMux I__2248 (
            .O(N__11620),
            .I(\uart_inst0.uart_inst0.tx_stateZ0Z_0 ));
    LocalMux I__2247 (
            .O(N__11613),
            .I(\uart_inst0.uart_inst0.tx_stateZ0Z_0 ));
    Odrv4 I__2246 (
            .O(N__11606),
            .I(\uart_inst0.uart_inst0.tx_stateZ0Z_0 ));
    InMux I__2245 (
            .O(N__11591),
            .I(N__11588));
    LocalMux I__2244 (
            .O(N__11588),
            .I(N__11584));
    InMux I__2243 (
            .O(N__11587),
            .I(N__11576));
    Span4Mux_h I__2242 (
            .O(N__11584),
            .I(N__11572));
    CascadeMux I__2241 (
            .O(N__11583),
            .I(N__11569));
    CascadeMux I__2240 (
            .O(N__11582),
            .I(N__11566));
    CascadeMux I__2239 (
            .O(N__11581),
            .I(N__11562));
    CascadeMux I__2238 (
            .O(N__11580),
            .I(N__11557));
    CascadeMux I__2237 (
            .O(N__11579),
            .I(N__11553));
    LocalMux I__2236 (
            .O(N__11576),
            .I(N__11549));
    InMux I__2235 (
            .O(N__11575),
            .I(N__11546));
    Span4Mux_v I__2234 (
            .O(N__11572),
            .I(N__11543));
    InMux I__2233 (
            .O(N__11569),
            .I(N__11540));
    InMux I__2232 (
            .O(N__11566),
            .I(N__11535));
    InMux I__2231 (
            .O(N__11565),
            .I(N__11535));
    InMux I__2230 (
            .O(N__11562),
            .I(N__11528));
    InMux I__2229 (
            .O(N__11561),
            .I(N__11528));
    InMux I__2228 (
            .O(N__11560),
            .I(N__11528));
    InMux I__2227 (
            .O(N__11557),
            .I(N__11521));
    InMux I__2226 (
            .O(N__11556),
            .I(N__11521));
    InMux I__2225 (
            .O(N__11553),
            .I(N__11521));
    InMux I__2224 (
            .O(N__11552),
            .I(N__11518));
    Odrv12 I__2223 (
            .O(N__11549),
            .I(\uart_inst0.uart_inst0.tx_stateZ0Z_1 ));
    LocalMux I__2222 (
            .O(N__11546),
            .I(\uart_inst0.uart_inst0.tx_stateZ0Z_1 ));
    Odrv4 I__2221 (
            .O(N__11543),
            .I(\uart_inst0.uart_inst0.tx_stateZ0Z_1 ));
    LocalMux I__2220 (
            .O(N__11540),
            .I(\uart_inst0.uart_inst0.tx_stateZ0Z_1 ));
    LocalMux I__2219 (
            .O(N__11535),
            .I(\uart_inst0.uart_inst0.tx_stateZ0Z_1 ));
    LocalMux I__2218 (
            .O(N__11528),
            .I(\uart_inst0.uart_inst0.tx_stateZ0Z_1 ));
    LocalMux I__2217 (
            .O(N__11521),
            .I(\uart_inst0.uart_inst0.tx_stateZ0Z_1 ));
    LocalMux I__2216 (
            .O(N__11518),
            .I(\uart_inst0.uart_inst0.tx_stateZ0Z_1 ));
    InMux I__2215 (
            .O(N__11501),
            .I(N__11498));
    LocalMux I__2214 (
            .O(N__11498),
            .I(N__11495));
    Odrv4 I__2213 (
            .O(N__11495),
            .I(\uart_inst0.uart_inst0.un1_m3_0_a2_0 ));
    InMux I__2212 (
            .O(N__11492),
            .I(N__11489));
    LocalMux I__2211 (
            .O(N__11489),
            .I(\uart_inst0.uart_inst0.N_275 ));
    CascadeMux I__2210 (
            .O(N__11486),
            .I(\uart_inst0.uart_inst0.N_283_cascade_ ));
    InMux I__2209 (
            .O(N__11483),
            .I(N__11479));
    InMux I__2208 (
            .O(N__11482),
            .I(N__11476));
    LocalMux I__2207 (
            .O(N__11479),
            .I(N__11473));
    LocalMux I__2206 (
            .O(N__11476),
            .I(N__11470));
    Odrv12 I__2205 (
            .O(N__11473),
            .I(\uart_inst0.uart_inst0.rx_stateZ0Z_6 ));
    Odrv4 I__2204 (
            .O(N__11470),
            .I(\uart_inst0.uart_inst0.rx_stateZ0Z_6 ));
    InMux I__2203 (
            .O(N__11465),
            .I(N__11459));
    InMux I__2202 (
            .O(N__11464),
            .I(N__11459));
    LocalMux I__2201 (
            .O(N__11459),
            .I(\uart_inst0.uart_inst0.rx_state_srsts_0_o2_3_3 ));
    InMux I__2200 (
            .O(N__11456),
            .I(N__11452));
    InMux I__2199 (
            .O(N__11455),
            .I(N__11449));
    LocalMux I__2198 (
            .O(N__11452),
            .I(\uart_inst0.uart_inst0.rx_countdown_2_sqmuxa_i_1 ));
    LocalMux I__2197 (
            .O(N__11449),
            .I(\uart_inst0.uart_inst0.rx_countdown_2_sqmuxa_i_1 ));
    InMux I__2196 (
            .O(N__11444),
            .I(N__11441));
    LocalMux I__2195 (
            .O(N__11441),
            .I(N__11438));
    Odrv12 I__2194 (
            .O(N__11438),
            .I(\uart_inst0.uart_inst0.un1_rx_clk_divider_0 ));
    CascadeMux I__2193 (
            .O(N__11435),
            .I(\uart_inst0.uart_inst0.N_258_0_cascade_ ));
    InMux I__2192 (
            .O(N__11432),
            .I(N__11425));
    InMux I__2191 (
            .O(N__11431),
            .I(N__11422));
    InMux I__2190 (
            .O(N__11430),
            .I(N__11419));
    InMux I__2189 (
            .O(N__11429),
            .I(N__11414));
    InMux I__2188 (
            .O(N__11428),
            .I(N__11414));
    LocalMux I__2187 (
            .O(N__11425),
            .I(\uart_inst0.uart_inst0.rx_countdownZ0Z_0 ));
    LocalMux I__2186 (
            .O(N__11422),
            .I(\uart_inst0.uart_inst0.rx_countdownZ0Z_0 ));
    LocalMux I__2185 (
            .O(N__11419),
            .I(\uart_inst0.uart_inst0.rx_countdownZ0Z_0 ));
    LocalMux I__2184 (
            .O(N__11414),
            .I(\uart_inst0.uart_inst0.rx_countdownZ0Z_0 ));
    InMux I__2183 (
            .O(N__11405),
            .I(N__11399));
    InMux I__2182 (
            .O(N__11404),
            .I(N__11396));
    InMux I__2181 (
            .O(N__11403),
            .I(N__11391));
    InMux I__2180 (
            .O(N__11402),
            .I(N__11391));
    LocalMux I__2179 (
            .O(N__11399),
            .I(\uart_inst0.uart_inst0.rx_countdownZ0Z_1 ));
    LocalMux I__2178 (
            .O(N__11396),
            .I(\uart_inst0.uart_inst0.rx_countdownZ0Z_1 ));
    LocalMux I__2177 (
            .O(N__11391),
            .I(\uart_inst0.uart_inst0.rx_countdownZ0Z_1 ));
    InMux I__2176 (
            .O(N__11384),
            .I(N__11381));
    LocalMux I__2175 (
            .O(N__11381),
            .I(\uart_inst0.uart_inst0.rx_countdown_s_1 ));
    InMux I__2174 (
            .O(N__11378),
            .I(\uart_inst0.uart_inst0.rx_countdown_cry_0 ));
    InMux I__2173 (
            .O(N__11375),
            .I(N__11371));
    InMux I__2172 (
            .O(N__11374),
            .I(N__11368));
    LocalMux I__2171 (
            .O(N__11371),
            .I(\uart_inst0.uart_inst0.rx_countdownZ0Z_2 ));
    LocalMux I__2170 (
            .O(N__11368),
            .I(\uart_inst0.uart_inst0.rx_countdownZ0Z_2 ));
    InMux I__2169 (
            .O(N__11363),
            .I(N__11360));
    LocalMux I__2168 (
            .O(N__11360),
            .I(\uart_inst0.uart_inst0.rx_countdown_s_2 ));
    InMux I__2167 (
            .O(N__11357),
            .I(\uart_inst0.uart_inst0.rx_countdown_cry_1 ));
    InMux I__2166 (
            .O(N__11354),
            .I(N__11350));
    InMux I__2165 (
            .O(N__11353),
            .I(N__11347));
    LocalMux I__2164 (
            .O(N__11350),
            .I(\uart_inst0.uart_inst0.rx_countdownZ0Z_3 ));
    LocalMux I__2163 (
            .O(N__11347),
            .I(\uart_inst0.uart_inst0.rx_countdownZ0Z_3 ));
    InMux I__2162 (
            .O(N__11342),
            .I(N__11339));
    LocalMux I__2161 (
            .O(N__11339),
            .I(\uart_inst0.uart_inst0.rx_countdown_s_3 ));
    InMux I__2160 (
            .O(N__11336),
            .I(\uart_inst0.uart_inst0.rx_countdown_cry_2 ));
    InMux I__2159 (
            .O(N__11333),
            .I(N__11328));
    InMux I__2158 (
            .O(N__11332),
            .I(N__11325));
    InMux I__2157 (
            .O(N__11331),
            .I(N__11322));
    LocalMux I__2156 (
            .O(N__11328),
            .I(\uart_inst0.uart_inst0.rx_countdownZ0Z_4 ));
    LocalMux I__2155 (
            .O(N__11325),
            .I(\uart_inst0.uart_inst0.rx_countdownZ0Z_4 ));
    LocalMux I__2154 (
            .O(N__11322),
            .I(\uart_inst0.uart_inst0.rx_countdownZ0Z_4 ));
    InMux I__2153 (
            .O(N__11315),
            .I(N__11311));
    InMux I__2152 (
            .O(N__11314),
            .I(N__11308));
    LocalMux I__2151 (
            .O(N__11311),
            .I(N__11305));
    LocalMux I__2150 (
            .O(N__11308),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ1Z_1 ));
    Odrv4 I__2149 (
            .O(N__11305),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ1Z_1 ));
    CascadeMux I__2148 (
            .O(N__11300),
            .I(N__11297));
    InMux I__2147 (
            .O(N__11297),
            .I(N__11293));
    InMux I__2146 (
            .O(N__11296),
            .I(N__11290));
    LocalMux I__2145 (
            .O(N__11293),
            .I(N__11287));
    LocalMux I__2144 (
            .O(N__11290),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ0Z_2 ));
    Odrv4 I__2143 (
            .O(N__11287),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ0Z_2 ));
    CascadeMux I__2142 (
            .O(N__11282),
            .I(N__11279));
    InMux I__2141 (
            .O(N__11279),
            .I(N__11276));
    LocalMux I__2140 (
            .O(N__11276),
            .I(N__11270));
    InMux I__2139 (
            .O(N__11275),
            .I(N__11267));
    InMux I__2138 (
            .O(N__11274),
            .I(N__11262));
    InMux I__2137 (
            .O(N__11273),
            .I(N__11262));
    Odrv4 I__2136 (
            .O(N__11270),
            .I(\uart_inst0.uart_inst0.rx_stateZ0Z_5 ));
    LocalMux I__2135 (
            .O(N__11267),
            .I(\uart_inst0.uart_inst0.rx_stateZ0Z_5 ));
    LocalMux I__2134 (
            .O(N__11262),
            .I(\uart_inst0.uart_inst0.rx_stateZ0Z_5 ));
    InMux I__2133 (
            .O(N__11255),
            .I(N__11252));
    LocalMux I__2132 (
            .O(N__11252),
            .I(N__11249));
    Odrv4 I__2131 (
            .O(N__11249),
            .I(rUartRxDataZ0Z_0));
    InMux I__2130 (
            .O(N__11246),
            .I(N__11231));
    InMux I__2129 (
            .O(N__11245),
            .I(N__11231));
    InMux I__2128 (
            .O(N__11244),
            .I(N__11231));
    InMux I__2127 (
            .O(N__11243),
            .I(N__11231));
    InMux I__2126 (
            .O(N__11242),
            .I(N__11231));
    LocalMux I__2125 (
            .O(N__11231),
            .I(N__11225));
    InMux I__2124 (
            .O(N__11230),
            .I(N__11218));
    InMux I__2123 (
            .O(N__11229),
            .I(N__11218));
    InMux I__2122 (
            .O(N__11228),
            .I(N__11218));
    Span4Mux_h I__2121 (
            .O(N__11225),
            .I(N__11211));
    LocalMux I__2120 (
            .O(N__11218),
            .I(N__11211));
    InMux I__2119 (
            .O(N__11217),
            .I(N__11208));
    InMux I__2118 (
            .O(N__11216),
            .I(N__11205));
    Odrv4 I__2117 (
            .O(N__11211),
            .I(rUartRxFlagZ0));
    LocalMux I__2116 (
            .O(N__11208),
            .I(rUartRxFlagZ0));
    LocalMux I__2115 (
            .O(N__11205),
            .I(rUartRxFlagZ0));
    InMux I__2114 (
            .O(N__11198),
            .I(N__11195));
    LocalMux I__2113 (
            .O(N__11195),
            .I(N__11192));
    Span4Mux_v I__2112 (
            .O(N__11192),
            .I(N__11189));
    Span4Mux_h I__2111 (
            .O(N__11189),
            .I(N__11186));
    Odrv4 I__2110 (
            .O(N__11186),
            .I(rUartTxDataZ0Z_0));
    CEMux I__2109 (
            .O(N__11183),
            .I(N__11180));
    LocalMux I__2108 (
            .O(N__11180),
            .I(N__11176));
    CEMux I__2107 (
            .O(N__11179),
            .I(N__11173));
    Odrv12 I__2106 (
            .O(N__11176),
            .I(rUartTxEn_4_0));
    LocalMux I__2105 (
            .O(N__11173),
            .I(rUartTxEn_4_0));
    CEMux I__2104 (
            .O(N__11168),
            .I(N__11164));
    CEMux I__2103 (
            .O(N__11167),
            .I(N__11161));
    LocalMux I__2102 (
            .O(N__11164),
            .I(rUartRxState_0_0));
    LocalMux I__2101 (
            .O(N__11161),
            .I(rUartRxState_0_0));
    InMux I__2100 (
            .O(N__11156),
            .I(N__11152));
    InMux I__2099 (
            .O(N__11155),
            .I(N__11148));
    LocalMux I__2098 (
            .O(N__11152),
            .I(N__11145));
    InMux I__2097 (
            .O(N__11151),
            .I(N__11142));
    LocalMux I__2096 (
            .O(N__11148),
            .I(N__11139));
    Span4Mux_v I__2095 (
            .O(N__11145),
            .I(N__11136));
    LocalMux I__2094 (
            .O(N__11142),
            .I(N__11131));
    Span4Mux_h I__2093 (
            .O(N__11139),
            .I(N__11131));
    Span4Mux_v I__2092 (
            .O(N__11136),
            .I(N__11123));
    Span4Mux_h I__2091 (
            .O(N__11131),
            .I(N__11123));
    InMux I__2090 (
            .O(N__11130),
            .I(N__11118));
    InMux I__2089 (
            .O(N__11129),
            .I(N__11118));
    InMux I__2088 (
            .O(N__11128),
            .I(N__11115));
    Odrv4 I__2087 (
            .O(N__11123),
            .I(\uart_inst0.uart_inst0.rx_stateZ0Z_0 ));
    LocalMux I__2086 (
            .O(N__11118),
            .I(\uart_inst0.uart_inst0.rx_stateZ0Z_0 ));
    LocalMux I__2085 (
            .O(N__11115),
            .I(\uart_inst0.uart_inst0.rx_stateZ0Z_0 ));
    CascadeMux I__2084 (
            .O(N__11108),
            .I(N__11105));
    InMux I__2083 (
            .O(N__11105),
            .I(N__11096));
    InMux I__2082 (
            .O(N__11104),
            .I(N__11096));
    InMux I__2081 (
            .O(N__11103),
            .I(N__11096));
    LocalMux I__2080 (
            .O(N__11096),
            .I(\uart_inst0.wRxWrEn_0 ));
    CascadeMux I__2079 (
            .O(N__11093),
            .I(N__11090));
    InMux I__2078 (
            .O(N__11090),
            .I(N__11087));
    LocalMux I__2077 (
            .O(N__11087),
            .I(N__11084));
    Span4Mux_h I__2076 (
            .O(N__11084),
            .I(N__11081));
    Odrv4 I__2075 (
            .O(N__11081),
            .I(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_0_0 ));
    InMux I__2074 (
            .O(N__11078),
            .I(N__11074));
    InMux I__2073 (
            .O(N__11077),
            .I(N__11071));
    LocalMux I__2072 (
            .O(N__11074),
            .I(N__11068));
    LocalMux I__2071 (
            .O(N__11071),
            .I(fifo_inst_rx_fifo_inst_rRamRdAddr_5));
    Odrv4 I__2070 (
            .O(N__11068),
            .I(fifo_inst_rx_fifo_inst_rRamRdAddr_5));
    InMux I__2069 (
            .O(N__11063),
            .I(N__11059));
    InMux I__2068 (
            .O(N__11062),
            .I(N__11056));
    LocalMux I__2067 (
            .O(N__11059),
            .I(fifo_inst_rx_fifo_inst_rRamRdAddr_4));
    LocalMux I__2066 (
            .O(N__11056),
            .I(fifo_inst_rx_fifo_inst_rRamRdAddr_4));
    InMux I__2065 (
            .O(N__11051),
            .I(N__11048));
    LocalMux I__2064 (
            .O(N__11048),
            .I(N__11045));
    Span4Mux_h I__2063 (
            .O(N__11045),
            .I(N__11041));
    InMux I__2062 (
            .O(N__11044),
            .I(N__11038));
    Odrv4 I__2061 (
            .O(N__11041),
            .I(fifo_inst_rx_fifo_inst_rRamRdAddr_2));
    LocalMux I__2060 (
            .O(N__11038),
            .I(fifo_inst_rx_fifo_inst_rRamRdAddr_2));
    InMux I__2059 (
            .O(N__11033),
            .I(N__11029));
    InMux I__2058 (
            .O(N__11032),
            .I(N__11026));
    LocalMux I__2057 (
            .O(N__11029),
            .I(N__11023));
    LocalMux I__2056 (
            .O(N__11026),
            .I(fifo_inst_rx_fifo_inst_rRamRdAddr_7));
    Odrv4 I__2055 (
            .O(N__11023),
            .I(fifo_inst_rx_fifo_inst_rRamRdAddr_7));
    InMux I__2054 (
            .O(N__11018),
            .I(N__11014));
    InMux I__2053 (
            .O(N__11017),
            .I(N__11011));
    LocalMux I__2052 (
            .O(N__11014),
            .I(N__11008));
    LocalMux I__2051 (
            .O(N__11011),
            .I(fifo_inst_rx_fifo_inst_rRamRdAddr_6));
    Odrv4 I__2050 (
            .O(N__11008),
            .I(fifo_inst_rx_fifo_inst_rRamRdAddr_6));
    CascadeMux I__2049 (
            .O(N__11003),
            .I(\uart_inst0.tx_uart_fifo_inst.m58_eZ0Z_5_cascade_ ));
    InMux I__2048 (
            .O(N__11000),
            .I(N__10997));
    LocalMux I__2047 (
            .O(N__10997),
            .I(\uart_inst0.tx_uart_fifo_inst.m58_eZ0Z_6 ));
    InMux I__2046 (
            .O(N__10994),
            .I(N__10989));
    InMux I__2045 (
            .O(N__10993),
            .I(N__10986));
    InMux I__2044 (
            .O(N__10992),
            .I(N__10983));
    LocalMux I__2043 (
            .O(N__10989),
            .I(\uart_inst0.tx_uart_fifo_inst.N_99 ));
    LocalMux I__2042 (
            .O(N__10986),
            .I(\uart_inst0.tx_uart_fifo_inst.N_99 ));
    LocalMux I__2041 (
            .O(N__10983),
            .I(\uart_inst0.tx_uart_fifo_inst.N_99 ));
    InMux I__2040 (
            .O(N__10976),
            .I(N__10970));
    InMux I__2039 (
            .O(N__10975),
            .I(N__10970));
    LocalMux I__2038 (
            .O(N__10970),
            .I(rRamRdAddr_RNI0S8U_0));
    CascadeMux I__2037 (
            .O(N__10967),
            .I(N__10963));
    InMux I__2036 (
            .O(N__10966),
            .I(N__10958));
    InMux I__2035 (
            .O(N__10963),
            .I(N__10955));
    InMux I__2034 (
            .O(N__10962),
            .I(N__10951));
    InMux I__2033 (
            .O(N__10961),
            .I(N__10948));
    LocalMux I__2032 (
            .O(N__10958),
            .I(N__10943));
    LocalMux I__2031 (
            .O(N__10955),
            .I(N__10943));
    CascadeMux I__2030 (
            .O(N__10954),
            .I(N__10939));
    LocalMux I__2029 (
            .O(N__10951),
            .I(N__10934));
    LocalMux I__2028 (
            .O(N__10948),
            .I(N__10934));
    Span4Mux_h I__2027 (
            .O(N__10943),
            .I(N__10931));
    InMux I__2026 (
            .O(N__10942),
            .I(N__10928));
    InMux I__2025 (
            .O(N__10939),
            .I(N__10925));
    Odrv4 I__2024 (
            .O(N__10934),
            .I(fifo_inst_rx_fifo_inst_wRamRdEn));
    Odrv4 I__2023 (
            .O(N__10931),
            .I(fifo_inst_rx_fifo_inst_wRamRdEn));
    LocalMux I__2022 (
            .O(N__10928),
            .I(fifo_inst_rx_fifo_inst_wRamRdEn));
    LocalMux I__2021 (
            .O(N__10925),
            .I(fifo_inst_rx_fifo_inst_wRamRdEn));
    CascadeMux I__2020 (
            .O(N__10916),
            .I(\uart_inst0.tx_uart_fifo_inst.N_99_cascade_ ));
    InMux I__2019 (
            .O(N__10913),
            .I(N__10909));
    InMux I__2018 (
            .O(N__10912),
            .I(N__10906));
    LocalMux I__2017 (
            .O(N__10909),
            .I(fifo_inst_rx_fifo_inst_rRamRdAddr_0));
    LocalMux I__2016 (
            .O(N__10906),
            .I(fifo_inst_rx_fifo_inst_rRamRdAddr_0));
    InMux I__2015 (
            .O(N__10901),
            .I(N__10898));
    LocalMux I__2014 (
            .O(N__10898),
            .I(N__10895));
    Odrv4 I__2013 (
            .O(N__10895),
            .I(rUartRxDataZ0Z_3));
    InMux I__2012 (
            .O(N__10892),
            .I(N__10889));
    LocalMux I__2011 (
            .O(N__10889),
            .I(N__10886));
    Span4Mux_v I__2010 (
            .O(N__10886),
            .I(N__10883));
    Span4Mux_h I__2009 (
            .O(N__10883),
            .I(N__10880));
    Odrv4 I__2008 (
            .O(N__10880),
            .I(rUartTxDataZ0Z_3));
    CascadeMux I__2007 (
            .O(N__10877),
            .I(N__10874));
    InMux I__2006 (
            .O(N__10874),
            .I(N__10871));
    LocalMux I__2005 (
            .O(N__10871),
            .I(N__10868));
    Odrv4 I__2004 (
            .O(N__10868),
            .I(rUartRxDataZ0Z_4));
    InMux I__2003 (
            .O(N__10865),
            .I(N__10862));
    LocalMux I__2002 (
            .O(N__10862),
            .I(rRxDataZ0Z_4));
    InMux I__2001 (
            .O(N__10859),
            .I(N__10856));
    LocalMux I__2000 (
            .O(N__10856),
            .I(N__10853));
    Span4Mux_v I__1999 (
            .O(N__10853),
            .I(N__10850));
    Odrv4 I__1998 (
            .O(N__10850),
            .I(rUartTxDataZ0Z_4));
    CascadeMux I__1997 (
            .O(N__10847),
            .I(N__10844));
    InMux I__1996 (
            .O(N__10844),
            .I(N__10841));
    LocalMux I__1995 (
            .O(N__10841),
            .I(rUartRxDataZ0Z_7));
    InMux I__1994 (
            .O(N__10838),
            .I(N__10835));
    LocalMux I__1993 (
            .O(N__10835),
            .I(N__10832));
    Span4Mux_v I__1992 (
            .O(N__10832),
            .I(N__10829));
    Odrv4 I__1991 (
            .O(N__10829),
            .I(rUartTxDataZ0Z_7));
    InMux I__1990 (
            .O(N__10826),
            .I(N__10823));
    LocalMux I__1989 (
            .O(N__10823),
            .I(N__10820));
    Odrv4 I__1988 (
            .O(N__10820),
            .I(rUartRxDataZ0Z_2));
    InMux I__1987 (
            .O(N__10817),
            .I(N__10814));
    LocalMux I__1986 (
            .O(N__10814),
            .I(N__10811));
    Span4Mux_v I__1985 (
            .O(N__10811),
            .I(N__10808));
    Span4Mux_h I__1984 (
            .O(N__10808),
            .I(N__10805));
    Odrv4 I__1983 (
            .O(N__10805),
            .I(rUartTxDataZ0Z_2));
    CascadeMux I__1982 (
            .O(N__10802),
            .I(N__10799));
    InMux I__1981 (
            .O(N__10799),
            .I(N__10796));
    LocalMux I__1980 (
            .O(N__10796),
            .I(N__10793));
    Span4Mux_h I__1979 (
            .O(N__10793),
            .I(N__10789));
    InMux I__1978 (
            .O(N__10792),
            .I(N__10786));
    Odrv4 I__1977 (
            .O(N__10789),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIM36CZ0 ));
    LocalMux I__1976 (
            .O(N__10786),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIM36CZ0 ));
    CascadeMux I__1975 (
            .O(N__10781),
            .I(N__10778));
    InMux I__1974 (
            .O(N__10778),
            .I(N__10775));
    LocalMux I__1973 (
            .O(N__10775),
            .I(N__10772));
    Span4Mux_s2_v I__1972 (
            .O(N__10772),
            .I(N__10769));
    Span4Mux_h I__1971 (
            .O(N__10769),
            .I(N__10765));
    InMux I__1970 (
            .O(N__10768),
            .I(N__10762));
    Odrv4 I__1969 (
            .O(N__10765),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIAHVBZ0 ));
    LocalMux I__1968 (
            .O(N__10762),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIAHVBZ0 ));
    InMux I__1967 (
            .O(N__10757),
            .I(N__10751));
    InMux I__1966 (
            .O(N__10756),
            .I(N__10751));
    LocalMux I__1965 (
            .O(N__10751),
            .I(un1_rRamRdAddr_cry_2_c_RNII9N9));
    CascadeMux I__1964 (
            .O(N__10748),
            .I(N__10745));
    InMux I__1963 (
            .O(N__10745),
            .I(N__10742));
    LocalMux I__1962 (
            .O(N__10742),
            .I(N__10739));
    Span4Mux_h I__1961 (
            .O(N__10739),
            .I(N__10736));
    Odrv4 I__1960 (
            .O(N__10736),
            .I(m60));
    CascadeMux I__1959 (
            .O(N__10733),
            .I(N__10730));
    InMux I__1958 (
            .O(N__10730),
            .I(N__10727));
    LocalMux I__1957 (
            .O(N__10727),
            .I(N__10724));
    Span4Mux_h I__1956 (
            .O(N__10724),
            .I(N__10720));
    InMux I__1955 (
            .O(N__10723),
            .I(N__10717));
    Odrv4 I__1954 (
            .O(N__10720),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIGQ2CZ0 ));
    LocalMux I__1953 (
            .O(N__10717),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIGQ2CZ0 ));
    InMux I__1952 (
            .O(N__10712),
            .I(N__10708));
    InMux I__1951 (
            .O(N__10711),
            .I(N__10705));
    LocalMux I__1950 (
            .O(N__10708),
            .I(fifo_inst_rx_fifo_inst_rRamRdAddr_3));
    LocalMux I__1949 (
            .O(N__10705),
            .I(fifo_inst_rx_fifo_inst_rRamRdAddr_3));
    InMux I__1948 (
            .O(N__10700),
            .I(N__10696));
    InMux I__1947 (
            .O(N__10699),
            .I(N__10693));
    LocalMux I__1946 (
            .O(N__10696),
            .I(fifo_inst_rx_fifo_inst_rRamRdAddr_1));
    LocalMux I__1945 (
            .O(N__10693),
            .I(fifo_inst_rx_fifo_inst_rRamRdAddr_1));
    CascadeMux I__1944 (
            .O(N__10688),
            .I(N__10684));
    InMux I__1943 (
            .O(N__10687),
            .I(N__10681));
    InMux I__1942 (
            .O(N__10684),
            .I(N__10678));
    LocalMux I__1941 (
            .O(N__10681),
            .I(fifo_inst_rx_fifo_inst_rRamRdAddr_8));
    LocalMux I__1940 (
            .O(N__10678),
            .I(fifo_inst_rx_fifo_inst_rRamRdAddr_8));
    InMux I__1939 (
            .O(N__10673),
            .I(N__10669));
    InMux I__1938 (
            .O(N__10672),
            .I(N__10666));
    LocalMux I__1937 (
            .O(N__10669),
            .I(N__10663));
    LocalMux I__1936 (
            .O(N__10666),
            .I(N_101));
    Odrv4 I__1935 (
            .O(N__10663),
            .I(N_101));
    InMux I__1934 (
            .O(N__10658),
            .I(N__10653));
    InMux I__1933 (
            .O(N__10657),
            .I(N__10649));
    InMux I__1932 (
            .O(N__10656),
            .I(N__10646));
    LocalMux I__1931 (
            .O(N__10653),
            .I(N__10643));
    InMux I__1930 (
            .O(N__10652),
            .I(N__10640));
    LocalMux I__1929 (
            .O(N__10649),
            .I(N__10637));
    LocalMux I__1928 (
            .O(N__10646),
            .I(N__10633));
    Span4Mux_v I__1927 (
            .O(N__10643),
            .I(N__10628));
    LocalMux I__1926 (
            .O(N__10640),
            .I(N__10628));
    Span4Mux_v I__1925 (
            .O(N__10637),
            .I(N__10625));
    InMux I__1924 (
            .O(N__10636),
            .I(N__10622));
    Odrv4 I__1923 (
            .O(N__10633),
            .I(N_97));
    Odrv4 I__1922 (
            .O(N__10628),
            .I(N_97));
    Odrv4 I__1921 (
            .O(N__10625),
            .I(N_97));
    LocalMux I__1920 (
            .O(N__10622),
            .I(N_97));
    CascadeMux I__1919 (
            .O(N__10613),
            .I(N__10610));
    InMux I__1918 (
            .O(N__10610),
            .I(N__10604));
    InMux I__1917 (
            .O(N__10609),
            .I(N__10601));
    InMux I__1916 (
            .O(N__10608),
            .I(N__10597));
    InMux I__1915 (
            .O(N__10607),
            .I(N__10594));
    LocalMux I__1914 (
            .O(N__10604),
            .I(N__10588));
    LocalMux I__1913 (
            .O(N__10601),
            .I(N__10588));
    InMux I__1912 (
            .O(N__10600),
            .I(N__10585));
    LocalMux I__1911 (
            .O(N__10597),
            .I(N__10582));
    LocalMux I__1910 (
            .O(N__10594),
            .I(N__10579));
    CascadeMux I__1909 (
            .O(N__10593),
            .I(N__10576));
    Span4Mux_v I__1908 (
            .O(N__10588),
            .I(N__10571));
    LocalMux I__1907 (
            .O(N__10585),
            .I(N__10571));
    Span4Mux_v I__1906 (
            .O(N__10582),
            .I(N__10566));
    Span4Mux_v I__1905 (
            .O(N__10579),
            .I(N__10566));
    InMux I__1904 (
            .O(N__10576),
            .I(N__10563));
    Span4Mux_v I__1903 (
            .O(N__10571),
            .I(N__10560));
    Sp12to4 I__1902 (
            .O(N__10566),
            .I(N__10555));
    LocalMux I__1901 (
            .O(N__10563),
            .I(N__10555));
    Span4Mux_h I__1900 (
            .O(N__10560),
            .I(N__10552));
    Span12Mux_h I__1899 (
            .O(N__10555),
            .I(N__10549));
    Sp12to4 I__1898 (
            .O(N__10552),
            .I(N__10546));
    Span12Mux_v I__1897 (
            .O(N__10549),
            .I(N__10543));
    Span12Mux_v I__1896 (
            .O(N__10546),
            .I(N__10540));
    Span12Mux_v I__1895 (
            .O(N__10543),
            .I(N__10537));
    Odrv12 I__1894 (
            .O(N__10540),
            .I(iTxE_n_c));
    Odrv12 I__1893 (
            .O(N__10537),
            .I(iTxE_n_c));
    InMux I__1892 (
            .O(N__10532),
            .I(N__10527));
    InMux I__1891 (
            .O(N__10531),
            .I(N__10520));
    InMux I__1890 (
            .O(N__10530),
            .I(N__10517));
    LocalMux I__1889 (
            .O(N__10527),
            .I(N__10514));
    InMux I__1888 (
            .O(N__10526),
            .I(N__10511));
    InMux I__1887 (
            .O(N__10525),
            .I(N__10508));
    InMux I__1886 (
            .O(N__10524),
            .I(N__10503));
    InMux I__1885 (
            .O(N__10523),
            .I(N__10503));
    LocalMux I__1884 (
            .O(N__10520),
            .I(N__10500));
    LocalMux I__1883 (
            .O(N__10517),
            .I(N__10496));
    Span4Mux_h I__1882 (
            .O(N__10514),
            .I(N__10491));
    LocalMux I__1881 (
            .O(N__10511),
            .I(N__10491));
    LocalMux I__1880 (
            .O(N__10508),
            .I(N__10484));
    LocalMux I__1879 (
            .O(N__10503),
            .I(N__10484));
    Span4Mux_h I__1878 (
            .O(N__10500),
            .I(N__10484));
    InMux I__1877 (
            .O(N__10499),
            .I(N__10481));
    Odrv4 I__1876 (
            .O(N__10496),
            .I(N_8_0));
    Odrv4 I__1875 (
            .O(N__10491),
            .I(N_8_0));
    Odrv4 I__1874 (
            .O(N__10484),
            .I(N_8_0));
    LocalMux I__1873 (
            .O(N__10481),
            .I(N_8_0));
    CascadeMux I__1872 (
            .O(N__10472),
            .I(fifo_inst_ft2232h_inst_un1_rFifoState_1_sqmuxa_0_i_cascade_));
    CEMux I__1871 (
            .O(N__10469),
            .I(N__10466));
    LocalMux I__1870 (
            .O(N__10466),
            .I(N__10463));
    Odrv4 I__1869 (
            .O(N__10463),
            .I(\fifo_inst.ft2232h_inst.un1_rFifoState_1_sqmuxa_0_i_0 ));
    CascadeMux I__1868 (
            .O(N__10460),
            .I(N__10457));
    InMux I__1867 (
            .O(N__10457),
            .I(N__10454));
    LocalMux I__1866 (
            .O(N__10454),
            .I(N__10451));
    Span4Mux_h I__1865 (
            .O(N__10451),
            .I(N__10448));
    Odrv4 I__1864 (
            .O(N__10448),
            .I(m59));
    CascadeMux I__1863 (
            .O(N__10445),
            .I(N__10442));
    InMux I__1862 (
            .O(N__10442),
            .I(N__10436));
    InMux I__1861 (
            .O(N__10441),
            .I(N__10436));
    LocalMux I__1860 (
            .O(N__10436),
            .I(un1_rRamRdAddr_cry_2_c_RNIMVKN));
    CascadeMux I__1859 (
            .O(N__10433),
            .I(N__10430));
    InMux I__1858 (
            .O(N__10430),
            .I(N__10427));
    LocalMux I__1857 (
            .O(N__10427),
            .I(N__10424));
    Span4Mux_s2_v I__1856 (
            .O(N__10424),
            .I(N__10421));
    Odrv4 I__1855 (
            .O(N__10421),
            .I(m74));
    InMux I__1854 (
            .O(N__10418),
            .I(N__10414));
    InMux I__1853 (
            .O(N__10417),
            .I(N__10411));
    LocalMux I__1852 (
            .O(N__10414),
            .I(fifo_inst_tx_fifo_inst_rRamRdAddr_5));
    LocalMux I__1851 (
            .O(N__10411),
            .I(fifo_inst_tx_fifo_inst_rRamRdAddr_5));
    InMux I__1850 (
            .O(N__10406),
            .I(N__10402));
    InMux I__1849 (
            .O(N__10405),
            .I(N__10399));
    LocalMux I__1848 (
            .O(N__10402),
            .I(fifo_inst_tx_fifo_inst_rRamRdAddr_7));
    LocalMux I__1847 (
            .O(N__10399),
            .I(fifo_inst_tx_fifo_inst_rRamRdAddr_7));
    InMux I__1846 (
            .O(N__10394),
            .I(N__10390));
    InMux I__1845 (
            .O(N__10393),
            .I(N__10387));
    LocalMux I__1844 (
            .O(N__10390),
            .I(fifo_inst_tx_fifo_inst_rRamRdAddr_6));
    LocalMux I__1843 (
            .O(N__10387),
            .I(fifo_inst_tx_fifo_inst_rRamRdAddr_6));
    CascadeMux I__1842 (
            .O(N__10382),
            .I(\uart_inst0.tx_uart_fifo_inst.m72_eZ0Z_5_cascade_ ));
    CascadeMux I__1841 (
            .O(N__10379),
            .I(\uart_inst0.tx_uart_fifo_inst.N_100_cascade_ ));
    CascadeMux I__1840 (
            .O(N__10376),
            .I(N__10373));
    InMux I__1839 (
            .O(N__10373),
            .I(N__10370));
    LocalMux I__1838 (
            .O(N__10370),
            .I(N__10367));
    Span4Mux_s2_v I__1837 (
            .O(N__10367),
            .I(N__10364));
    Odrv4 I__1836 (
            .O(N__10364),
            .I(m73));
    InMux I__1835 (
            .O(N__10361),
            .I(N__10357));
    InMux I__1834 (
            .O(N__10360),
            .I(N__10354));
    LocalMux I__1833 (
            .O(N__10357),
            .I(fifo_inst_tx_fifo_inst_rRamRdAddr_3));
    LocalMux I__1832 (
            .O(N__10354),
            .I(fifo_inst_tx_fifo_inst_rRamRdAddr_3));
    InMux I__1831 (
            .O(N__10349),
            .I(N__10345));
    InMux I__1830 (
            .O(N__10348),
            .I(N__10342));
    LocalMux I__1829 (
            .O(N__10345),
            .I(fifo_inst_tx_fifo_inst_rRamRdAddr_1));
    LocalMux I__1828 (
            .O(N__10342),
            .I(fifo_inst_tx_fifo_inst_rRamRdAddr_1));
    CascadeMux I__1827 (
            .O(N__10337),
            .I(N__10334));
    InMux I__1826 (
            .O(N__10334),
            .I(N__10330));
    InMux I__1825 (
            .O(N__10333),
            .I(N__10327));
    LocalMux I__1824 (
            .O(N__10330),
            .I(N__10324));
    LocalMux I__1823 (
            .O(N__10327),
            .I(fifo_inst_tx_fifo_inst_rRamRdAddr_8));
    Odrv4 I__1822 (
            .O(N__10324),
            .I(fifo_inst_tx_fifo_inst_rRamRdAddr_8));
    InMux I__1821 (
            .O(N__10319),
            .I(N__10316));
    LocalMux I__1820 (
            .O(N__10316),
            .I(\uart_inst0.tx_uart_fifo_inst.m72_eZ0Z_6 ));
    CascadeMux I__1819 (
            .O(N__10313),
            .I(N__10310));
    InMux I__1818 (
            .O(N__10310),
            .I(N__10307));
    LocalMux I__1817 (
            .O(N__10307),
            .I(N__10304));
    Span4Mux_s2_v I__1816 (
            .O(N__10304),
            .I(N__10300));
    InMux I__1815 (
            .O(N__10303),
            .I(N__10297));
    Odrv4 I__1814 (
            .O(N__10300),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIKG0QZ0 ));
    LocalMux I__1813 (
            .O(N__10297),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIKG0QZ0 ));
    InMux I__1812 (
            .O(N__10292),
            .I(N__10288));
    InMux I__1811 (
            .O(N__10291),
            .I(N__10285));
    LocalMux I__1810 (
            .O(N__10288),
            .I(fifo_inst_tx_fifo_inst_rRamRdAddr_4));
    LocalMux I__1809 (
            .O(N__10285),
            .I(fifo_inst_tx_fifo_inst_rRamRdAddr_4));
    InMux I__1808 (
            .O(N__10280),
            .I(N__10266));
    InMux I__1807 (
            .O(N__10279),
            .I(N__10266));
    InMux I__1806 (
            .O(N__10278),
            .I(N__10266));
    InMux I__1805 (
            .O(N__10277),
            .I(N__10266));
    CEMux I__1804 (
            .O(N__10276),
            .I(N__10262));
    CascadeMux I__1803 (
            .O(N__10275),
            .I(N__10259));
    LocalMux I__1802 (
            .O(N__10266),
            .I(N__10256));
    InMux I__1801 (
            .O(N__10265),
            .I(N__10253));
    LocalMux I__1800 (
            .O(N__10262),
            .I(N__10250));
    InMux I__1799 (
            .O(N__10259),
            .I(N__10247));
    Odrv4 I__1798 (
            .O(N__10256),
            .I(fifo_inst_tx_fifo_inst_wRamRdEn));
    LocalMux I__1797 (
            .O(N__10253),
            .I(fifo_inst_tx_fifo_inst_wRamRdEn));
    Odrv4 I__1796 (
            .O(N__10250),
            .I(fifo_inst_tx_fifo_inst_wRamRdEn));
    LocalMux I__1795 (
            .O(N__10247),
            .I(fifo_inst_tx_fifo_inst_wRamRdEn));
    CascadeMux I__1794 (
            .O(N__10238),
            .I(N__10235));
    InMux I__1793 (
            .O(N__10235),
            .I(N__10229));
    InMux I__1792 (
            .O(N__10234),
            .I(N__10229));
    LocalMux I__1791 (
            .O(N__10229),
            .I(rRamRdAddr_RNI9KL42_0));
    InMux I__1790 (
            .O(N__10226),
            .I(N__10217));
    InMux I__1789 (
            .O(N__10225),
            .I(N__10217));
    InMux I__1788 (
            .O(N__10224),
            .I(N__10217));
    LocalMux I__1787 (
            .O(N__10217),
            .I(\uart_inst0.tx_uart_fifo_inst.N_100 ));
    InMux I__1786 (
            .O(N__10214),
            .I(N__10210));
    InMux I__1785 (
            .O(N__10213),
            .I(N__10207));
    LocalMux I__1784 (
            .O(N__10210),
            .I(fifo_inst_tx_fifo_inst_rRamRdAddr_0));
    LocalMux I__1783 (
            .O(N__10207),
            .I(fifo_inst_tx_fifo_inst_rRamRdAddr_0));
    CascadeMux I__1782 (
            .O(N__10202),
            .I(\uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_11_3_cascade_ ));
    InMux I__1781 (
            .O(N__10199),
            .I(N__10191));
    InMux I__1780 (
            .O(N__10198),
            .I(N__10191));
    InMux I__1779 (
            .O(N__10197),
            .I(N__10188));
    InMux I__1778 (
            .O(N__10196),
            .I(N__10185));
    LocalMux I__1777 (
            .O(N__10191),
            .I(\uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13 ));
    LocalMux I__1776 (
            .O(N__10188),
            .I(\uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13 ));
    LocalMux I__1775 (
            .O(N__10185),
            .I(\uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13 ));
    CascadeMux I__1774 (
            .O(N__10178),
            .I(N__10175));
    InMux I__1773 (
            .O(N__10175),
            .I(N__10170));
    InMux I__1772 (
            .O(N__10174),
            .I(N__10167));
    InMux I__1771 (
            .O(N__10173),
            .I(N__10164));
    LocalMux I__1770 (
            .O(N__10170),
            .I(N__10157));
    LocalMux I__1769 (
            .O(N__10167),
            .I(N__10154));
    LocalMux I__1768 (
            .O(N__10164),
            .I(N__10151));
    InMux I__1767 (
            .O(N__10163),
            .I(N__10148));
    CascadeMux I__1766 (
            .O(N__10162),
            .I(N__10144));
    InMux I__1765 (
            .O(N__10161),
            .I(N__10138));
    InMux I__1764 (
            .O(N__10160),
            .I(N__10138));
    Span4Mux_h I__1763 (
            .O(N__10157),
            .I(N__10135));
    Span12Mux_h I__1762 (
            .O(N__10154),
            .I(N__10132));
    Span4Mux_h I__1761 (
            .O(N__10151),
            .I(N__10127));
    LocalMux I__1760 (
            .O(N__10148),
            .I(N__10127));
    InMux I__1759 (
            .O(N__10147),
            .I(N__10122));
    InMux I__1758 (
            .O(N__10144),
            .I(N__10122));
    InMux I__1757 (
            .O(N__10143),
            .I(N__10119));
    LocalMux I__1756 (
            .O(N__10138),
            .I(wTxFull));
    Odrv4 I__1755 (
            .O(N__10135),
            .I(wTxFull));
    Odrv12 I__1754 (
            .O(N__10132),
            .I(wTxFull));
    Odrv4 I__1753 (
            .O(N__10127),
            .I(wTxFull));
    LocalMux I__1752 (
            .O(N__10122),
            .I(wTxFull));
    LocalMux I__1751 (
            .O(N__10119),
            .I(wTxFull));
    InMux I__1750 (
            .O(N__10106),
            .I(N__10103));
    LocalMux I__1749 (
            .O(N__10103),
            .I(N__10099));
    InMux I__1748 (
            .O(N__10102),
            .I(N__10096));
    Span12Mux_v I__1747 (
            .O(N__10099),
            .I(N__10093));
    LocalMux I__1746 (
            .O(N__10096),
            .I(rTxDataZ0Z_0));
    Odrv12 I__1745 (
            .O(N__10093),
            .I(rTxDataZ0Z_0));
    IoInMux I__1744 (
            .O(N__10088),
            .I(N__10084));
    IoInMux I__1743 (
            .O(N__10087),
            .I(N__10081));
    LocalMux I__1742 (
            .O(N__10084),
            .I(N__10076));
    LocalMux I__1741 (
            .O(N__10081),
            .I(N__10076));
    IoSpan4Mux I__1740 (
            .O(N__10076),
            .I(N__10072));
    IoInMux I__1739 (
            .O(N__10075),
            .I(N__10069));
    Span4Mux_s3_v I__1738 (
            .O(N__10072),
            .I(N__10065));
    LocalMux I__1737 (
            .O(N__10069),
            .I(N__10061));
    IoInMux I__1736 (
            .O(N__10068),
            .I(N__10058));
    Sp12to4 I__1735 (
            .O(N__10065),
            .I(N__10052));
    IoInMux I__1734 (
            .O(N__10064),
            .I(N__10049));
    IoSpan4Mux I__1733 (
            .O(N__10061),
            .I(N__10044));
    LocalMux I__1732 (
            .O(N__10058),
            .I(N__10044));
    IoInMux I__1731 (
            .O(N__10057),
            .I(N__10041));
    IoInMux I__1730 (
            .O(N__10056),
            .I(N__10038));
    IoInMux I__1729 (
            .O(N__10055),
            .I(N__10035));
    Span12Mux_v I__1728 (
            .O(N__10052),
            .I(N__10032));
    LocalMux I__1727 (
            .O(N__10049),
            .I(N__10029));
    IoSpan4Mux I__1726 (
            .O(N__10044),
            .I(N__10024));
    LocalMux I__1725 (
            .O(N__10041),
            .I(N__10024));
    LocalMux I__1724 (
            .O(N__10038),
            .I(N__10021));
    LocalMux I__1723 (
            .O(N__10035),
            .I(N__10018));
    Span12Mux_v I__1722 (
            .O(N__10032),
            .I(N__10015));
    Span4Mux_s1_v I__1721 (
            .O(N__10029),
            .I(N__10012));
    Span4Mux_s1_v I__1720 (
            .O(N__10024),
            .I(N__10009));
    Span4Mux_s1_v I__1719 (
            .O(N__10021),
            .I(N__10004));
    Span4Mux_s1_v I__1718 (
            .O(N__10018),
            .I(N__10004));
    Odrv12 I__1717 (
            .O(N__10015),
            .I(rTxBusReady));
    Odrv4 I__1716 (
            .O(N__10012),
            .I(rTxBusReady));
    Odrv4 I__1715 (
            .O(N__10009),
            .I(rTxBusReady));
    Odrv4 I__1714 (
            .O(N__10004),
            .I(rTxBusReady));
    CascadeMux I__1713 (
            .O(N__9995),
            .I(\uart_inst0.uart_inst0.tx_state_ns_0_0_0_cascade_ ));
    InMux I__1712 (
            .O(N__9992),
            .I(N__9989));
    LocalMux I__1711 (
            .O(N__9989),
            .I(N__9985));
    InMux I__1710 (
            .O(N__9988),
            .I(N__9982));
    Odrv4 I__1709 (
            .O(N__9985),
            .I(\uart_inst0.uart_inst0.tx_state_1_sqmuxa_1_0_a3_0 ));
    LocalMux I__1708 (
            .O(N__9982),
            .I(\uart_inst0.uart_inst0.tx_state_1_sqmuxa_1_0_a3_0 ));
    SRMux I__1707 (
            .O(N__9977),
            .I(N__9974));
    LocalMux I__1706 (
            .O(N__9974),
            .I(N__9971));
    Span4Mux_h I__1705 (
            .O(N__9971),
            .I(N__9967));
    InMux I__1704 (
            .O(N__9970),
            .I(N__9964));
    Odrv4 I__1703 (
            .O(N__9967),
            .I(\uart_inst0.uart_inst0.tx_state_RNI1319Z0Z_0 ));
    LocalMux I__1702 (
            .O(N__9964),
            .I(\uart_inst0.uart_inst0.tx_state_RNI1319Z0Z_0 ));
    InMux I__1701 (
            .O(N__9959),
            .I(N__9952));
    InMux I__1700 (
            .O(N__9958),
            .I(N__9947));
    InMux I__1699 (
            .O(N__9957),
            .I(N__9947));
    InMux I__1698 (
            .O(N__9956),
            .I(N__9944));
    InMux I__1697 (
            .O(N__9955),
            .I(N__9941));
    LocalMux I__1696 (
            .O(N__9952),
            .I(N__9938));
    LocalMux I__1695 (
            .O(N__9947),
            .I(\uart_inst0.uart_inst0.tx_bits_remainingZ0Z_1 ));
    LocalMux I__1694 (
            .O(N__9944),
            .I(\uart_inst0.uart_inst0.tx_bits_remainingZ0Z_1 ));
    LocalMux I__1693 (
            .O(N__9941),
            .I(\uart_inst0.uart_inst0.tx_bits_remainingZ0Z_1 ));
    Odrv4 I__1692 (
            .O(N__9938),
            .I(\uart_inst0.uart_inst0.tx_bits_remainingZ0Z_1 ));
    InMux I__1691 (
            .O(N__9929),
            .I(N__9918));
    InMux I__1690 (
            .O(N__9928),
            .I(N__9918));
    InMux I__1689 (
            .O(N__9927),
            .I(N__9918));
    InMux I__1688 (
            .O(N__9926),
            .I(N__9915));
    InMux I__1687 (
            .O(N__9925),
            .I(N__9912));
    LocalMux I__1686 (
            .O(N__9918),
            .I(\uart_inst0.uart_inst0.tx_bits_remainingZ0Z_0 ));
    LocalMux I__1685 (
            .O(N__9915),
            .I(\uart_inst0.uart_inst0.tx_bits_remainingZ0Z_0 ));
    LocalMux I__1684 (
            .O(N__9912),
            .I(\uart_inst0.uart_inst0.tx_bits_remainingZ0Z_0 ));
    CascadeMux I__1683 (
            .O(N__9905),
            .I(\uart_inst0.uart_inst0.un1_tx_bits_remaining_ac0_1_a0_0_cascade_ ));
    InMux I__1682 (
            .O(N__9902),
            .I(N__9899));
    LocalMux I__1681 (
            .O(N__9899),
            .I(\uart_inst0.uart_inst0.un1_tx_bits_remaining_ac0_1 ));
    CascadeMux I__1680 (
            .O(N__9896),
            .I(\uart_inst0.uart_inst0.un1_rx_state49_i_cascade_ ));
    CascadeMux I__1679 (
            .O(N__9893),
            .I(\uart_inst0.uart_inst0.tx_countdown_RNO_0Z0Z_3_cascade_ ));
    CascadeMux I__1678 (
            .O(N__9890),
            .I(\uart_inst0.uart_inst0.N_147_0_cascade_ ));
    CascadeMux I__1677 (
            .O(N__9887),
            .I(\uart_inst0.uart_inst0.N_277_cascade_ ));
    InMux I__1676 (
            .O(N__9884),
            .I(N__9881));
    LocalMux I__1675 (
            .O(N__9881),
            .I(\uart_inst0.uart_inst0.rx_state_srsts_0_a5_1_0 ));
    CascadeMux I__1674 (
            .O(N__9878),
            .I(\uart_inst0.uart_inst0.N_280_cascade_ ));
    InMux I__1673 (
            .O(N__9875),
            .I(N__9870));
    InMux I__1672 (
            .O(N__9874),
            .I(N__9865));
    InMux I__1671 (
            .O(N__9873),
            .I(N__9865));
    LocalMux I__1670 (
            .O(N__9870),
            .I(\uart_inst0.uart_inst0.rx_stateZ0Z_4 ));
    LocalMux I__1669 (
            .O(N__9865),
            .I(\uart_inst0.uart_inst0.rx_stateZ0Z_4 ));
    InMux I__1668 (
            .O(N__9860),
            .I(N__9857));
    LocalMux I__1667 (
            .O(N__9857),
            .I(\uart_inst0.uart_inst0.N_261_0 ));
    InMux I__1666 (
            .O(N__9854),
            .I(N__9851));
    LocalMux I__1665 (
            .O(N__9851),
            .I(N__9845));
    CascadeMux I__1664 (
            .O(N__9850),
            .I(N__9842));
    InMux I__1663 (
            .O(N__9849),
            .I(N__9839));
    CascadeMux I__1662 (
            .O(N__9848),
            .I(N__9836));
    Span4Mux_h I__1661 (
            .O(N__9845),
            .I(N__9833));
    InMux I__1660 (
            .O(N__9842),
            .I(N__9829));
    LocalMux I__1659 (
            .O(N__9839),
            .I(N__9826));
    InMux I__1658 (
            .O(N__9836),
            .I(N__9823));
    Span4Mux_v I__1657 (
            .O(N__9833),
            .I(N__9820));
    InMux I__1656 (
            .O(N__9832),
            .I(N__9817));
    LocalMux I__1655 (
            .O(N__9829),
            .I(N__9814));
    Odrv4 I__1654 (
            .O(N__9826),
            .I(\uart_inst0.wTxRdEmpty ));
    LocalMux I__1653 (
            .O(N__9823),
            .I(\uart_inst0.wTxRdEmpty ));
    Odrv4 I__1652 (
            .O(N__9820),
            .I(\uart_inst0.wTxRdEmpty ));
    LocalMux I__1651 (
            .O(N__9817),
            .I(\uart_inst0.wTxRdEmpty ));
    Odrv12 I__1650 (
            .O(N__9814),
            .I(\uart_inst0.wTxRdEmpty ));
    CascadeMux I__1649 (
            .O(N__9803),
            .I(\uart_inst0.uart_inst0.rx_state_srsts_0_o2_3_3_cascade_ ));
    CascadeMux I__1648 (
            .O(N__9800),
            .I(\uart_inst0.uart_inst0.N_257_0_cascade_ ));
    CascadeMux I__1647 (
            .O(N__9797),
            .I(N__9793));
    InMux I__1646 (
            .O(N__9796),
            .I(N__9789));
    InMux I__1645 (
            .O(N__9793),
            .I(N__9786));
    InMux I__1644 (
            .O(N__9792),
            .I(N__9783));
    LocalMux I__1643 (
            .O(N__9789),
            .I(N__9780));
    LocalMux I__1642 (
            .O(N__9786),
            .I(\uart_inst0.uart_inst0.tx_bits_remainingZ0Z_2 ));
    LocalMux I__1641 (
            .O(N__9783),
            .I(\uart_inst0.uart_inst0.tx_bits_remainingZ0Z_2 ));
    Odrv4 I__1640 (
            .O(N__9780),
            .I(\uart_inst0.uart_inst0.tx_bits_remainingZ0Z_2 ));
    CascadeMux I__1639 (
            .O(N__9773),
            .I(N__9770));
    InMux I__1638 (
            .O(N__9770),
            .I(N__9767));
    LocalMux I__1637 (
            .O(N__9767),
            .I(N__9763));
    InMux I__1636 (
            .O(N__9766),
            .I(N__9760));
    Span4Mux_h I__1635 (
            .O(N__9763),
            .I(N__9757));
    LocalMux I__1634 (
            .O(N__9760),
            .I(\uart_inst0.uart_inst0.tx_bits_remainingZ0Z_3 ));
    Odrv4 I__1633 (
            .O(N__9757),
            .I(\uart_inst0.uart_inst0.tx_bits_remainingZ0Z_3 ));
    CascadeMux I__1632 (
            .O(N__9752),
            .I(N__9749));
    InMux I__1631 (
            .O(N__9749),
            .I(N__9743));
    InMux I__1630 (
            .O(N__9748),
            .I(N__9743));
    LocalMux I__1629 (
            .O(N__9743),
            .I(\uart_inst0.uart_inst0.N_157 ));
    CascadeMux I__1628 (
            .O(N__9740),
            .I(\uart_inst0.uart_inst0.N_157_cascade_ ));
    CascadeMux I__1627 (
            .O(N__9737),
            .I(N__9734));
    InMux I__1626 (
            .O(N__9734),
            .I(N__9731));
    LocalMux I__1625 (
            .O(N__9731),
            .I(N__9728));
    Odrv12 I__1624 (
            .O(N__9728),
            .I(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_3 ));
    InMux I__1623 (
            .O(N__9725),
            .I(N__9721));
    InMux I__1622 (
            .O(N__9724),
            .I(N__9718));
    LocalMux I__1621 (
            .O(N__9721),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIUJZ0Z84 ));
    LocalMux I__1620 (
            .O(N__9718),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIUJZ0Z84 ));
    InMux I__1619 (
            .O(N__9713),
            .I(N__9710));
    LocalMux I__1618 (
            .O(N__9710),
            .I(N__9706));
    InMux I__1617 (
            .O(N__9709),
            .I(N__9703));
    Odrv4 I__1616 (
            .O(N__9706),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_4 ));
    LocalMux I__1615 (
            .O(N__9703),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_4 ));
    InMux I__1614 (
            .O(N__9698),
            .I(N__9695));
    LocalMux I__1613 (
            .O(N__9695),
            .I(N__9691));
    InMux I__1612 (
            .O(N__9694),
            .I(N__9688));
    Odrv4 I__1611 (
            .O(N__9691),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_5 ));
    LocalMux I__1610 (
            .O(N__9688),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_5 ));
    InMux I__1609 (
            .O(N__9683),
            .I(N__9679));
    InMux I__1608 (
            .O(N__9682),
            .I(N__9676));
    LocalMux I__1607 (
            .O(N__9679),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNI2QAZ0Z4 ));
    LocalMux I__1606 (
            .O(N__9676),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNI2QAZ0Z4 ));
    InMux I__1605 (
            .O(N__9671),
            .I(N__9668));
    LocalMux I__1604 (
            .O(N__9668),
            .I(N__9664));
    InMux I__1603 (
            .O(N__9667),
            .I(N__9661));
    Odrv4 I__1602 (
            .O(N__9664),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_6 ));
    LocalMux I__1601 (
            .O(N__9661),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_6 ));
    InMux I__1600 (
            .O(N__9656),
            .I(N__9652));
    InMux I__1599 (
            .O(N__9655),
            .I(N__9649));
    LocalMux I__1598 (
            .O(N__9652),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI4TBZ0Z4 ));
    LocalMux I__1597 (
            .O(N__9649),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI4TBZ0Z4 ));
    CascadeMux I__1596 (
            .O(N__9644),
            .I(N__9641));
    InMux I__1595 (
            .O(N__9641),
            .I(N__9638));
    LocalMux I__1594 (
            .O(N__9638),
            .I(N__9635));
    Span4Mux_v I__1593 (
            .O(N__9635),
            .I(N__9631));
    InMux I__1592 (
            .O(N__9634),
            .I(N__9628));
    Odrv4 I__1591 (
            .O(N__9631),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_7 ));
    LocalMux I__1590 (
            .O(N__9628),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_7 ));
    InMux I__1589 (
            .O(N__9623),
            .I(N__9619));
    InMux I__1588 (
            .O(N__9622),
            .I(N__9616));
    LocalMux I__1587 (
            .O(N__9619),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI60DZ0Z4 ));
    LocalMux I__1586 (
            .O(N__9616),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI60DZ0Z4 ));
    InMux I__1585 (
            .O(N__9611),
            .I(N__9607));
    InMux I__1584 (
            .O(N__9610),
            .I(N__9604));
    LocalMux I__1583 (
            .O(N__9607),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_8 ));
    LocalMux I__1582 (
            .O(N__9604),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_8 ));
    CascadeMux I__1581 (
            .O(N__9599),
            .I(\uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_5_cascade_ ));
    CascadeMux I__1580 (
            .O(N__9596),
            .I(\uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7_cascade_ ));
    CEMux I__1579 (
            .O(N__9593),
            .I(N__9584));
    CascadeMux I__1578 (
            .O(N__9592),
            .I(N__9581));
    InMux I__1577 (
            .O(N__9591),
            .I(N__9578));
    InMux I__1576 (
            .O(N__9590),
            .I(N__9571));
    InMux I__1575 (
            .O(N__9589),
            .I(N__9571));
    InMux I__1574 (
            .O(N__9588),
            .I(N__9571));
    InMux I__1573 (
            .O(N__9587),
            .I(N__9568));
    LocalMux I__1572 (
            .O(N__9584),
            .I(N__9565));
    InMux I__1571 (
            .O(N__9581),
            .I(N__9562));
    LocalMux I__1570 (
            .O(N__9578),
            .I(\uart_inst0.tx_uart_fifo_inst.wRamRdEn_1 ));
    LocalMux I__1569 (
            .O(N__9571),
            .I(\uart_inst0.tx_uart_fifo_inst.wRamRdEn_1 ));
    LocalMux I__1568 (
            .O(N__9568),
            .I(\uart_inst0.tx_uart_fifo_inst.wRamRdEn_1 ));
    Odrv4 I__1567 (
            .O(N__9565),
            .I(\uart_inst0.tx_uart_fifo_inst.wRamRdEn_1 ));
    LocalMux I__1566 (
            .O(N__9562),
            .I(\uart_inst0.tx_uart_fifo_inst.wRamRdEn_1 ));
    CascadeMux I__1565 (
            .O(N__9551),
            .I(N__9548));
    InMux I__1564 (
            .O(N__9548),
            .I(N__9545));
    LocalMux I__1563 (
            .O(N__9545),
            .I(N__9542));
    Span4Mux_v I__1562 (
            .O(N__9542),
            .I(N__9539));
    Odrv4 I__1561 (
            .O(N__9539),
            .I(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0 ));
    InMux I__1560 (
            .O(N__9536),
            .I(N__9530));
    InMux I__1559 (
            .O(N__9535),
            .I(N__9530));
    LocalMux I__1558 (
            .O(N__9530),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIBDOK2Z0Z_0 ));
    CascadeMux I__1557 (
            .O(N__9527),
            .I(N__9523));
    InMux I__1556 (
            .O(N__9526),
            .I(N__9519));
    InMux I__1555 (
            .O(N__9523),
            .I(N__9514));
    InMux I__1554 (
            .O(N__9522),
            .I(N__9514));
    LocalMux I__1553 (
            .O(N__9519),
            .I(\uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7 ));
    LocalMux I__1552 (
            .O(N__9514),
            .I(\uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7 ));
    InMux I__1551 (
            .O(N__9509),
            .I(N__9501));
    InMux I__1550 (
            .O(N__9508),
            .I(N__9501));
    InMux I__1549 (
            .O(N__9507),
            .I(N__9496));
    CascadeMux I__1548 (
            .O(N__9506),
            .I(N__9493));
    LocalMux I__1547 (
            .O(N__9501),
            .I(N__9490));
    InMux I__1546 (
            .O(N__9500),
            .I(N__9484));
    InMux I__1545 (
            .O(N__9499),
            .I(N__9481));
    LocalMux I__1544 (
            .O(N__9496),
            .I(N__9478));
    InMux I__1543 (
            .O(N__9493),
            .I(N__9475));
    Span4Mux_v I__1542 (
            .O(N__9490),
            .I(N__9472));
    InMux I__1541 (
            .O(N__9489),
            .I(N__9465));
    InMux I__1540 (
            .O(N__9488),
            .I(N__9465));
    InMux I__1539 (
            .O(N__9487),
            .I(N__9465));
    LocalMux I__1538 (
            .O(N__9484),
            .I(\uart_inst0.wTxRdEn_0 ));
    LocalMux I__1537 (
            .O(N__9481),
            .I(\uart_inst0.wTxRdEn_0 ));
    Odrv4 I__1536 (
            .O(N__9478),
            .I(\uart_inst0.wTxRdEn_0 ));
    LocalMux I__1535 (
            .O(N__9475),
            .I(\uart_inst0.wTxRdEn_0 ));
    Odrv4 I__1534 (
            .O(N__9472),
            .I(\uart_inst0.wTxRdEn_0 ));
    LocalMux I__1533 (
            .O(N__9465),
            .I(\uart_inst0.wTxRdEn_0 ));
    CascadeMux I__1532 (
            .O(N__9452),
            .I(N__9449));
    InMux I__1531 (
            .O(N__9449),
            .I(N__9446));
    LocalMux I__1530 (
            .O(N__9446),
            .I(N__9443));
    Odrv12 I__1529 (
            .O(N__9443),
            .I(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_5 ));
    CascadeMux I__1528 (
            .O(N__9440),
            .I(N__9437));
    InMux I__1527 (
            .O(N__9437),
            .I(N__9434));
    LocalMux I__1526 (
            .O(N__9434),
            .I(N__9431));
    Odrv12 I__1525 (
            .O(N__9431),
            .I(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_6 ));
    CascadeMux I__1524 (
            .O(N__9428),
            .I(N__9425));
    InMux I__1523 (
            .O(N__9425),
            .I(N__9422));
    LocalMux I__1522 (
            .O(N__9422),
            .I(N__9419));
    Odrv12 I__1521 (
            .O(N__9419),
            .I(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_7 ));
    InMux I__1520 (
            .O(N__9416),
            .I(N__9412));
    InMux I__1519 (
            .O(N__9415),
            .I(N__9409));
    LocalMux I__1518 (
            .O(N__9412),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_0 ));
    LocalMux I__1517 (
            .O(N__9409),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_0 ));
    InMux I__1516 (
            .O(N__9404),
            .I(N__9400));
    InMux I__1515 (
            .O(N__9403),
            .I(N__9397));
    LocalMux I__1514 (
            .O(N__9400),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_3 ));
    LocalMux I__1513 (
            .O(N__9397),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_3 ));
    InMux I__1512 (
            .O(N__9392),
            .I(N__9389));
    LocalMux I__1511 (
            .O(N__9389),
            .I(\uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_4 ));
    InMux I__1510 (
            .O(N__9386),
            .I(N__9383));
    LocalMux I__1509 (
            .O(N__9383),
            .I(rUartRxDataZ0Z_5));
    InMux I__1508 (
            .O(N__9380),
            .I(N__9377));
    LocalMux I__1507 (
            .O(N__9377),
            .I(rUartRxDataZ0Z_6));
    InMux I__1506 (
            .O(N__9374),
            .I(N__9371));
    LocalMux I__1505 (
            .O(N__9371),
            .I(N__9368));
    Odrv4 I__1504 (
            .O(N__9368),
            .I(rUartRxDataZ0Z_1));
    CascadeMux I__1503 (
            .O(N__9365),
            .I(N__9362));
    InMux I__1502 (
            .O(N__9362),
            .I(N__9359));
    LocalMux I__1501 (
            .O(N__9359),
            .I(N__9356));
    Span4Mux_h I__1500 (
            .O(N__9356),
            .I(N__9353));
    Odrv4 I__1499 (
            .O(N__9353),
            .I(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_2 ));
    CascadeMux I__1498 (
            .O(N__9350),
            .I(N__9346));
    InMux I__1497 (
            .O(N__9349),
            .I(N__9341));
    InMux I__1496 (
            .O(N__9346),
            .I(N__9341));
    LocalMux I__1495 (
            .O(N__9341),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNISGZ0Z74 ));
    InMux I__1494 (
            .O(N__9338),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_6 ));
    InMux I__1493 (
            .O(N__9335),
            .I(bfn_15_6_0_));
    CascadeMux I__1492 (
            .O(N__9332),
            .I(N__9329));
    InMux I__1491 (
            .O(N__9329),
            .I(N__9326));
    LocalMux I__1490 (
            .O(N__9326),
            .I(N__9323));
    Span4Mux_h I__1489 (
            .O(N__9323),
            .I(N__9319));
    InMux I__1488 (
            .O(N__9322),
            .I(N__9316));
    Odrv4 I__1487 (
            .O(N__9319),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIIT3CZ0 ));
    LocalMux I__1486 (
            .O(N__9316),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIIT3CZ0 ));
    InMux I__1485 (
            .O(N__9311),
            .I(N__9307));
    InMux I__1484 (
            .O(N__9310),
            .I(N__9304));
    LocalMux I__1483 (
            .O(N__9307),
            .I(N__9299));
    LocalMux I__1482 (
            .O(N__9304),
            .I(N__9296));
    InMux I__1481 (
            .O(N__9303),
            .I(N__9292));
    InMux I__1480 (
            .O(N__9302),
            .I(N__9289));
    Span4Mux_v I__1479 (
            .O(N__9299),
            .I(N__9283));
    Span4Mux_v I__1478 (
            .O(N__9296),
            .I(N__9283));
    InMux I__1477 (
            .O(N__9295),
            .I(N__9280));
    LocalMux I__1476 (
            .O(N__9292),
            .I(N__9275));
    LocalMux I__1475 (
            .O(N__9289),
            .I(N__9275));
    InMux I__1474 (
            .O(N__9288),
            .I(N__9272));
    Odrv4 I__1473 (
            .O(N__9283),
            .I(rTxEnZ0));
    LocalMux I__1472 (
            .O(N__9280),
            .I(rTxEnZ0));
    Odrv4 I__1471 (
            .O(N__9275),
            .I(rTxEnZ0));
    LocalMux I__1470 (
            .O(N__9272),
            .I(rTxEnZ0));
    CascadeMux I__1469 (
            .O(N__9263),
            .I(N__9260));
    InMux I__1468 (
            .O(N__9260),
            .I(N__9254));
    CascadeMux I__1467 (
            .O(N__9259),
            .I(N__9248));
    InMux I__1466 (
            .O(N__9258),
            .I(N__9243));
    InMux I__1465 (
            .O(N__9257),
            .I(N__9243));
    LocalMux I__1464 (
            .O(N__9254),
            .I(N__9240));
    InMux I__1463 (
            .O(N__9253),
            .I(N__9232));
    InMux I__1462 (
            .O(N__9252),
            .I(N__9232));
    InMux I__1461 (
            .O(N__9251),
            .I(N__9227));
    InMux I__1460 (
            .O(N__9248),
            .I(N__9227));
    LocalMux I__1459 (
            .O(N__9243),
            .I(N__9222));
    Span4Mux_v I__1458 (
            .O(N__9240),
            .I(N__9222));
    InMux I__1457 (
            .O(N__9239),
            .I(N__9219));
    InMux I__1456 (
            .O(N__9238),
            .I(N__9214));
    InMux I__1455 (
            .O(N__9237),
            .I(N__9214));
    LocalMux I__1454 (
            .O(N__9232),
            .I(fifo_inst_wTxRdEn));
    LocalMux I__1453 (
            .O(N__9227),
            .I(fifo_inst_wTxRdEn));
    Odrv4 I__1452 (
            .O(N__9222),
            .I(fifo_inst_wTxRdEn));
    LocalMux I__1451 (
            .O(N__9219),
            .I(fifo_inst_wTxRdEn));
    LocalMux I__1450 (
            .O(N__9214),
            .I(fifo_inst_wTxRdEn));
    InMux I__1449 (
            .O(N__9203),
            .I(N__9197));
    InMux I__1448 (
            .O(N__9202),
            .I(N__9197));
    LocalMux I__1447 (
            .O(N__9197),
            .I(N__9194));
    Span4Mux_v I__1446 (
            .O(N__9194),
            .I(N__9191));
    Odrv4 I__1445 (
            .O(N__9191),
            .I(fifo_inst_tx_fifo_inst_rDataCount_0_sqmuxa));
    CascadeMux I__1444 (
            .O(N__9188),
            .I(N__9184));
    InMux I__1443 (
            .O(N__9187),
            .I(N__9180));
    InMux I__1442 (
            .O(N__9184),
            .I(N__9174));
    InMux I__1441 (
            .O(N__9183),
            .I(N__9174));
    LocalMux I__1440 (
            .O(N__9180),
            .I(N__9171));
    InMux I__1439 (
            .O(N__9179),
            .I(N__9168));
    LocalMux I__1438 (
            .O(N__9174),
            .I(fifo_inst_ft2232h_inst_rWrDelay));
    Odrv4 I__1437 (
            .O(N__9171),
            .I(fifo_inst_ft2232h_inst_rWrDelay));
    LocalMux I__1436 (
            .O(N__9168),
            .I(fifo_inst_ft2232h_inst_rWrDelay));
    InMux I__1435 (
            .O(N__9161),
            .I(N__9156));
    InMux I__1434 (
            .O(N__9160),
            .I(N__9150));
    InMux I__1433 (
            .O(N__9159),
            .I(N__9150));
    LocalMux I__1432 (
            .O(N__9156),
            .I(N__9147));
    InMux I__1431 (
            .O(N__9155),
            .I(N__9144));
    LocalMux I__1430 (
            .O(N__9150),
            .I(fifo_inst_ft2232h_inst_rFifoState_4));
    Odrv4 I__1429 (
            .O(N__9147),
            .I(fifo_inst_ft2232h_inst_rFifoState_4));
    LocalMux I__1428 (
            .O(N__9144),
            .I(fifo_inst_ft2232h_inst_rFifoState_4));
    CascadeMux I__1427 (
            .O(N__9137),
            .I(N__9134));
    InMux I__1426 (
            .O(N__9134),
            .I(N__9131));
    LocalMux I__1425 (
            .O(N__9131),
            .I(N__9128));
    Span4Mux_h I__1424 (
            .O(N__9128),
            .I(N__9124));
    InMux I__1423 (
            .O(N__9127),
            .I(N__9121));
    Odrv4 I__1422 (
            .O(N__9124),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNIO67CZ0 ));
    LocalMux I__1421 (
            .O(N__9121),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNIO67CZ0 ));
    InMux I__1420 (
            .O(N__9116),
            .I(N__9113));
    LocalMux I__1419 (
            .O(N__9113),
            .I(N__9110));
    Span4Mux_v I__1418 (
            .O(N__9110),
            .I(N__9107));
    Odrv4 I__1417 (
            .O(N__9107),
            .I(rUartTxDataZ0Z_6));
    InMux I__1416 (
            .O(N__9104),
            .I(N__9101));
    LocalMux I__1415 (
            .O(N__9101),
            .I(N__9098));
    Span4Mux_v I__1414 (
            .O(N__9098),
            .I(N__9095));
    Odrv4 I__1413 (
            .O(N__9095),
            .I(rUartTxDataZ0Z_5));
    InMux I__1412 (
            .O(N__9092),
            .I(N__9089));
    LocalMux I__1411 (
            .O(N__9089),
            .I(N__9086));
    Span4Mux_v I__1410 (
            .O(N__9086),
            .I(N__9083));
    Span4Mux_h I__1409 (
            .O(N__9083),
            .I(N__9080));
    Odrv4 I__1408 (
            .O(N__9080),
            .I(rUartTxDataZ0Z_1));
    InMux I__1407 (
            .O(N__9077),
            .I(N__9066));
    InMux I__1406 (
            .O(N__9076),
            .I(N__9066));
    InMux I__1405 (
            .O(N__9075),
            .I(N__9061));
    InMux I__1404 (
            .O(N__9074),
            .I(N__9061));
    InMux I__1403 (
            .O(N__9073),
            .I(N__9056));
    InMux I__1402 (
            .O(N__9072),
            .I(N__9056));
    InMux I__1401 (
            .O(N__9071),
            .I(N__9053));
    LocalMux I__1400 (
            .O(N__9066),
            .I(fifo_inst_wRxWrEn));
    LocalMux I__1399 (
            .O(N__9061),
            .I(fifo_inst_wRxWrEn));
    LocalMux I__1398 (
            .O(N__9056),
            .I(fifo_inst_wRxWrEn));
    LocalMux I__1397 (
            .O(N__9053),
            .I(fifo_inst_wRxWrEn));
    InMux I__1396 (
            .O(N__9044),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_0 ));
    CascadeMux I__1395 (
            .O(N__9041),
            .I(N__9038));
    InMux I__1394 (
            .O(N__9038),
            .I(N__9035));
    LocalMux I__1393 (
            .O(N__9035),
            .I(N__9032));
    Span4Mux_v I__1392 (
            .O(N__9032),
            .I(N__9028));
    InMux I__1391 (
            .O(N__9031),
            .I(N__9025));
    Odrv4 I__1390 (
            .O(N__9028),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNICK0CZ0 ));
    LocalMux I__1389 (
            .O(N__9025),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNICK0CZ0 ));
    InMux I__1388 (
            .O(N__9020),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_1 ));
    InMux I__1387 (
            .O(N__9017),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_2 ));
    InMux I__1386 (
            .O(N__9014),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_3 ));
    InMux I__1385 (
            .O(N__9011),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_4 ));
    CascadeMux I__1384 (
            .O(N__9008),
            .I(N__9005));
    InMux I__1383 (
            .O(N__9005),
            .I(N__9002));
    LocalMux I__1382 (
            .O(N__9002),
            .I(N__8999));
    Span4Mux_s2_v I__1381 (
            .O(N__8999),
            .I(N__8996));
    Span4Mux_h I__1380 (
            .O(N__8996),
            .I(N__8992));
    InMux I__1379 (
            .O(N__8995),
            .I(N__8989));
    Odrv4 I__1378 (
            .O(N__8992),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIK05CZ0 ));
    LocalMux I__1377 (
            .O(N__8989),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIK05CZ0 ));
    InMux I__1376 (
            .O(N__8984),
            .I(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_5 ));
    InMux I__1375 (
            .O(N__8981),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_2 ));
    InMux I__1374 (
            .O(N__8978),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_3 ));
    CascadeMux I__1373 (
            .O(N__8975),
            .I(N__8972));
    InMux I__1372 (
            .O(N__8972),
            .I(N__8969));
    LocalMux I__1371 (
            .O(N__8969),
            .I(N__8966));
    Span4Mux_s2_v I__1370 (
            .O(N__8966),
            .I(N__8962));
    InMux I__1369 (
            .O(N__8965),
            .I(N__8959));
    Odrv4 I__1368 (
            .O(N__8962),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIMJ1QZ0 ));
    LocalMux I__1367 (
            .O(N__8959),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIMJ1QZ0 ));
    InMux I__1366 (
            .O(N__8954),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_4 ));
    CascadeMux I__1365 (
            .O(N__8951),
            .I(N__8948));
    InMux I__1364 (
            .O(N__8948),
            .I(N__8945));
    LocalMux I__1363 (
            .O(N__8945),
            .I(N__8942));
    Span4Mux_h I__1362 (
            .O(N__8942),
            .I(N__8938));
    InMux I__1361 (
            .O(N__8941),
            .I(N__8935));
    Odrv4 I__1360 (
            .O(N__8938),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIOM2QZ0 ));
    LocalMux I__1359 (
            .O(N__8935),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIOM2QZ0 ));
    InMux I__1358 (
            .O(N__8930),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_5 ));
    CascadeMux I__1357 (
            .O(N__8927),
            .I(N__8924));
    InMux I__1356 (
            .O(N__8924),
            .I(N__8921));
    LocalMux I__1355 (
            .O(N__8921),
            .I(N__8918));
    Span4Mux_h I__1354 (
            .O(N__8918),
            .I(N__8914));
    InMux I__1353 (
            .O(N__8917),
            .I(N__8911));
    Odrv4 I__1352 (
            .O(N__8914),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIQP3QZ0 ));
    LocalMux I__1351 (
            .O(N__8911),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIQP3QZ0 ));
    InMux I__1350 (
            .O(N__8906),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_6 ));
    InMux I__1349 (
            .O(N__8903),
            .I(bfn_15_4_0_));
    CascadeMux I__1348 (
            .O(N__8900),
            .I(N__8897));
    InMux I__1347 (
            .O(N__8897),
            .I(N__8894));
    LocalMux I__1346 (
            .O(N__8894),
            .I(N__8891));
    Span4Mux_h I__1345 (
            .O(N__8891),
            .I(N__8887));
    InMux I__1344 (
            .O(N__8890),
            .I(N__8884));
    Odrv4 I__1343 (
            .O(N__8887),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIE7TPZ0 ));
    LocalMux I__1342 (
            .O(N__8884),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIE7TPZ0 ));
    CascadeMux I__1341 (
            .O(N__8879),
            .I(N__8876));
    InMux I__1340 (
            .O(N__8876),
            .I(N__8873));
    LocalMux I__1339 (
            .O(N__8873),
            .I(N__8870));
    Span4Mux_h I__1338 (
            .O(N__8870),
            .I(N__8866));
    InMux I__1337 (
            .O(N__8869),
            .I(N__8863));
    Odrv4 I__1336 (
            .O(N__8866),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNISS4QZ0 ));
    LocalMux I__1335 (
            .O(N__8863),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNISS4QZ0 ));
    InMux I__1334 (
            .O(N__8858),
            .I(N__8855));
    LocalMux I__1333 (
            .O(N__8855),
            .I(N__8852));
    Span4Mux_s1_v I__1332 (
            .O(N__8852),
            .I(N__8849));
    Odrv4 I__1331 (
            .O(N__8849),
            .I(\fifo_inst.tx_fifo_inst.ram512x8_inst.mem_0 ));
    IoInMux I__1330 (
            .O(N__8846),
            .I(N__8843));
    LocalMux I__1329 (
            .O(N__8843),
            .I(N__8840));
    Span4Mux_s0_v I__1328 (
            .O(N__8840),
            .I(N__8837));
    Odrv4 I__1327 (
            .O(N__8837),
            .I(wTxRdData_0));
    InMux I__1326 (
            .O(N__8834),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_0 ));
    InMux I__1325 (
            .O(N__8831),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_1 ));
    InMux I__1324 (
            .O(N__8828),
            .I(N__8825));
    LocalMux I__1323 (
            .O(N__8825),
            .I(\uart_inst0.uart_inst0.N_141_0 ));
    InMux I__1322 (
            .O(N__8822),
            .I(N__8819));
    LocalMux I__1321 (
            .O(N__8819),
            .I(\uart_inst0.uart_inst0.N_143_0 ));
    CascadeMux I__1320 (
            .O(N__8816),
            .I(\uart_inst0.uart_inst0.N_143_0_cascade_ ));
    CEMux I__1319 (
            .O(N__8813),
            .I(N__8810));
    LocalMux I__1318 (
            .O(N__8810),
            .I(N__8807));
    Span4Mux_v I__1317 (
            .O(N__8807),
            .I(N__8803));
    CEMux I__1316 (
            .O(N__8806),
            .I(N__8800));
    Odrv4 I__1315 (
            .O(N__8803),
            .I(\uart_inst0.uart_inst0.N_143_0_0 ));
    LocalMux I__1314 (
            .O(N__8800),
            .I(\uart_inst0.uart_inst0.N_143_0_0 ));
    CascadeMux I__1313 (
            .O(N__8795),
            .I(N__8792));
    InMux I__1312 (
            .O(N__8792),
            .I(N__8789));
    LocalMux I__1311 (
            .O(N__8789),
            .I(\uart_inst0.uart_inst0.un1_m3_0_a2_2_1 ));
    CascadeMux I__1310 (
            .O(N__8786),
            .I(\uart_inst0.uart_inst0.N_136_0_cascade_ ));
    InMux I__1309 (
            .O(N__8783),
            .I(N__8780));
    LocalMux I__1308 (
            .O(N__8780),
            .I(\uart_inst0.uart_inst0.un1_tx_bits_remaining_c1 ));
    InMux I__1307 (
            .O(N__8777),
            .I(N__8772));
    InMux I__1306 (
            .O(N__8776),
            .I(N__8767));
    InMux I__1305 (
            .O(N__8775),
            .I(N__8767));
    LocalMux I__1304 (
            .O(N__8772),
            .I(\uart_inst0.uart_inst0.N_136_0 ));
    LocalMux I__1303 (
            .O(N__8767),
            .I(\uart_inst0.uart_inst0.N_136_0 ));
    InMux I__1302 (
            .O(N__8762),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_3 ));
    InMux I__1301 (
            .O(N__8759),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_4 ));
    InMux I__1300 (
            .O(N__8756),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_5 ));
    InMux I__1299 (
            .O(N__8753),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_6 ));
    InMux I__1298 (
            .O(N__8750),
            .I(bfn_14_12_0_));
    CascadeMux I__1297 (
            .O(N__8747),
            .I(N__8744));
    InMux I__1296 (
            .O(N__8744),
            .I(N__8739));
    InMux I__1295 (
            .O(N__8743),
            .I(N__8736));
    InMux I__1294 (
            .O(N__8742),
            .I(N__8733));
    LocalMux I__1293 (
            .O(N__8739),
            .I(N__8730));
    LocalMux I__1292 (
            .O(N__8736),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_7 ));
    LocalMux I__1291 (
            .O(N__8733),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_7 ));
    Odrv12 I__1290 (
            .O(N__8730),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_7 ));
    CascadeMux I__1289 (
            .O(N__8723),
            .I(N__8720));
    InMux I__1288 (
            .O(N__8720),
            .I(N__8717));
    LocalMux I__1287 (
            .O(N__8717),
            .I(N__8714));
    Span4Mux_h I__1286 (
            .O(N__8714),
            .I(N__8709));
    InMux I__1285 (
            .O(N__8713),
            .I(N__8706));
    InMux I__1284 (
            .O(N__8712),
            .I(N__8703));
    Odrv4 I__1283 (
            .O(N__8709),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_5 ));
    LocalMux I__1282 (
            .O(N__8706),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_5 ));
    LocalMux I__1281 (
            .O(N__8703),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_5 ));
    CascadeMux I__1280 (
            .O(N__8696),
            .I(N__8693));
    InMux I__1279 (
            .O(N__8693),
            .I(N__8689));
    CascadeMux I__1278 (
            .O(N__8692),
            .I(N__8686));
    LocalMux I__1277 (
            .O(N__8689),
            .I(N__8682));
    InMux I__1276 (
            .O(N__8686),
            .I(N__8679));
    InMux I__1275 (
            .O(N__8685),
            .I(N__8676));
    Odrv12 I__1274 (
            .O(N__8682),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_6 ));
    LocalMux I__1273 (
            .O(N__8679),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_6 ));
    LocalMux I__1272 (
            .O(N__8676),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_6 ));
    CascadeMux I__1271 (
            .O(N__8669),
            .I(N__8666));
    InMux I__1270 (
            .O(N__8666),
            .I(N__8663));
    LocalMux I__1269 (
            .O(N__8663),
            .I(N__8658));
    InMux I__1268 (
            .O(N__8662),
            .I(N__8655));
    InMux I__1267 (
            .O(N__8661),
            .I(N__8652));
    Odrv12 I__1266 (
            .O(N__8658),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_4 ));
    LocalMux I__1265 (
            .O(N__8655),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_4 ));
    LocalMux I__1264 (
            .O(N__8652),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_4 ));
    CascadeMux I__1263 (
            .O(N__8645),
            .I(N__8641));
    CascadeMux I__1262 (
            .O(N__8644),
            .I(N__8638));
    InMux I__1261 (
            .O(N__8641),
            .I(N__8635));
    InMux I__1260 (
            .O(N__8638),
            .I(N__8632));
    LocalMux I__1259 (
            .O(N__8635),
            .I(N__8629));
    LocalMux I__1258 (
            .O(N__8632),
            .I(N__8626));
    Span4Mux_h I__1257 (
            .O(N__8629),
            .I(N__8623));
    Span4Mux_h I__1256 (
            .O(N__8626),
            .I(N__8620));
    Odrv4 I__1255 (
            .O(N__8623),
            .I(\uart_inst0.tx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_5 ));
    Odrv4 I__1254 (
            .O(N__8620),
            .I(\uart_inst0.tx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_5 ));
    IoInMux I__1253 (
            .O(N__8615),
            .I(N__8612));
    LocalMux I__1252 (
            .O(N__8612),
            .I(N__8609));
    IoSpan4Mux I__1251 (
            .O(N__8609),
            .I(N__8606));
    Span4Mux_s0_v I__1250 (
            .O(N__8606),
            .I(N__8603));
    Sp12to4 I__1249 (
            .O(N__8603),
            .I(N__8599));
    CascadeMux I__1248 (
            .O(N__8602),
            .I(N__8596));
    Span12Mux_v I__1247 (
            .O(N__8599),
            .I(N__8593));
    InMux I__1246 (
            .O(N__8596),
            .I(N__8590));
    Odrv12 I__1245 (
            .O(N__8593),
            .I(P1A7_c));
    LocalMux I__1244 (
            .O(N__8590),
            .I(P1A7_c));
    InMux I__1243 (
            .O(N__8585),
            .I(N__8576));
    InMux I__1242 (
            .O(N__8584),
            .I(N__8563));
    InMux I__1241 (
            .O(N__8583),
            .I(N__8563));
    InMux I__1240 (
            .O(N__8582),
            .I(N__8563));
    InMux I__1239 (
            .O(N__8581),
            .I(N__8563));
    InMux I__1238 (
            .O(N__8580),
            .I(N__8563));
    InMux I__1237 (
            .O(N__8579),
            .I(N__8559));
    LocalMux I__1236 (
            .O(N__8576),
            .I(N__8556));
    InMux I__1235 (
            .O(N__8575),
            .I(N__8551));
    InMux I__1234 (
            .O(N__8574),
            .I(N__8551));
    LocalMux I__1233 (
            .O(N__8563),
            .I(N__8548));
    InMux I__1232 (
            .O(N__8562),
            .I(N__8545));
    LocalMux I__1231 (
            .O(N__8559),
            .I(\uart_inst0.uart_inst0.tx_state_81_d ));
    Odrv4 I__1230 (
            .O(N__8556),
            .I(\uart_inst0.uart_inst0.tx_state_81_d ));
    LocalMux I__1229 (
            .O(N__8551),
            .I(\uart_inst0.uart_inst0.tx_state_81_d ));
    Odrv4 I__1228 (
            .O(N__8548),
            .I(\uart_inst0.uart_inst0.tx_state_81_d ));
    LocalMux I__1227 (
            .O(N__8545),
            .I(\uart_inst0.uart_inst0.tx_state_81_d ));
    InMux I__1226 (
            .O(N__8534),
            .I(N__8531));
    LocalMux I__1225 (
            .O(N__8531),
            .I(\uart_inst0.uart_inst0.rTxDataZ0Z_0 ));
    InMux I__1224 (
            .O(N__8528),
            .I(N__8525));
    LocalMux I__1223 (
            .O(N__8525),
            .I(\uart_inst0.uart_inst0.rTx_6_f1_0 ));
    InMux I__1222 (
            .O(N__8522),
            .I(N__8519));
    LocalMux I__1221 (
            .O(N__8519),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c2 ));
    CascadeMux I__1220 (
            .O(N__8516),
            .I(N__8511));
    InMux I__1219 (
            .O(N__8515),
            .I(N__8506));
    InMux I__1218 (
            .O(N__8514),
            .I(N__8502));
    InMux I__1217 (
            .O(N__8511),
            .I(N__8499));
    CEMux I__1216 (
            .O(N__8510),
            .I(N__8496));
    CascadeMux I__1215 (
            .O(N__8509),
            .I(N__8493));
    LocalMux I__1214 (
            .O(N__8506),
            .I(N__8488));
    InMux I__1213 (
            .O(N__8505),
            .I(N__8485));
    LocalMux I__1212 (
            .O(N__8502),
            .I(N__8480));
    LocalMux I__1211 (
            .O(N__8499),
            .I(N__8480));
    LocalMux I__1210 (
            .O(N__8496),
            .I(N__8477));
    InMux I__1209 (
            .O(N__8493),
            .I(N__8470));
    InMux I__1208 (
            .O(N__8492),
            .I(N__8470));
    InMux I__1207 (
            .O(N__8491),
            .I(N__8467));
    Span4Mux_v I__1206 (
            .O(N__8488),
            .I(N__8462));
    LocalMux I__1205 (
            .O(N__8485),
            .I(N__8462));
    Span4Mux_h I__1204 (
            .O(N__8480),
            .I(N__8457));
    Span4Mux_h I__1203 (
            .O(N__8477),
            .I(N__8457));
    InMux I__1202 (
            .O(N__8476),
            .I(N__8454));
    InMux I__1201 (
            .O(N__8475),
            .I(N__8451));
    LocalMux I__1200 (
            .O(N__8470),
            .I(N__8448));
    LocalMux I__1199 (
            .O(N__8467),
            .I(N__8445));
    Span4Mux_v I__1198 (
            .O(N__8462),
            .I(N__8440));
    Span4Mux_v I__1197 (
            .O(N__8457),
            .I(N__8440));
    LocalMux I__1196 (
            .O(N__8454),
            .I(\uart_inst0.tx_uart_fifo_inst.wRamWrEn_1 ));
    LocalMux I__1195 (
            .O(N__8451),
            .I(\uart_inst0.tx_uart_fifo_inst.wRamWrEn_1 ));
    Odrv4 I__1194 (
            .O(N__8448),
            .I(\uart_inst0.tx_uart_fifo_inst.wRamWrEn_1 ));
    Odrv12 I__1193 (
            .O(N__8445),
            .I(\uart_inst0.tx_uart_fifo_inst.wRamWrEn_1 ));
    Odrv4 I__1192 (
            .O(N__8440),
            .I(\uart_inst0.tx_uart_fifo_inst.wRamWrEn_1 ));
    CascadeMux I__1191 (
            .O(N__8429),
            .I(N__8426));
    InMux I__1190 (
            .O(N__8426),
            .I(N__8423));
    LocalMux I__1189 (
            .O(N__8423),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rDataCount_axbxc1_0 ));
    InMux I__1188 (
            .O(N__8420),
            .I(N__8414));
    InMux I__1187 (
            .O(N__8419),
            .I(N__8414));
    LocalMux I__1186 (
            .O(N__8414),
            .I(N__8411));
    Span4Mux_v I__1185 (
            .O(N__8411),
            .I(N__8404));
    InMux I__1184 (
            .O(N__8410),
            .I(N__8401));
    InMux I__1183 (
            .O(N__8409),
            .I(N__8394));
    InMux I__1182 (
            .O(N__8408),
            .I(N__8394));
    InMux I__1181 (
            .O(N__8407),
            .I(N__8394));
    Odrv4 I__1180 (
            .O(N__8404),
            .I(\uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_1 ));
    LocalMux I__1179 (
            .O(N__8401),
            .I(\uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_1 ));
    LocalMux I__1178 (
            .O(N__8394),
            .I(\uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_1 ));
    InMux I__1177 (
            .O(N__8387),
            .I(N__8383));
    CascadeMux I__1176 (
            .O(N__8386),
            .I(N__8378));
    LocalMux I__1175 (
            .O(N__8383),
            .I(N__8375));
    InMux I__1174 (
            .O(N__8382),
            .I(N__8370));
    InMux I__1173 (
            .O(N__8381),
            .I(N__8370));
    InMux I__1172 (
            .O(N__8378),
            .I(N__8367));
    Odrv12 I__1171 (
            .O(N__8375),
            .I(\uart_inst0.tx_uart_fifo_inst.rDataCountZ0Z_2 ));
    LocalMux I__1170 (
            .O(N__8370),
            .I(\uart_inst0.tx_uart_fifo_inst.rDataCountZ0Z_2 ));
    LocalMux I__1169 (
            .O(N__8367),
            .I(\uart_inst0.tx_uart_fifo_inst.rDataCountZ0Z_2 ));
    CascadeMux I__1168 (
            .O(N__8360),
            .I(N__8357));
    InMux I__1167 (
            .O(N__8357),
            .I(N__8352));
    InMux I__1166 (
            .O(N__8356),
            .I(N__8346));
    InMux I__1165 (
            .O(N__8355),
            .I(N__8343));
    LocalMux I__1164 (
            .O(N__8352),
            .I(N__8340));
    InMux I__1163 (
            .O(N__8351),
            .I(N__8337));
    InMux I__1162 (
            .O(N__8350),
            .I(N__8332));
    InMux I__1161 (
            .O(N__8349),
            .I(N__8332));
    LocalMux I__1160 (
            .O(N__8346),
            .I(\uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_0 ));
    LocalMux I__1159 (
            .O(N__8343),
            .I(\uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_0 ));
    Odrv12 I__1158 (
            .O(N__8340),
            .I(\uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_0 ));
    LocalMux I__1157 (
            .O(N__8337),
            .I(\uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_0 ));
    LocalMux I__1156 (
            .O(N__8332),
            .I(\uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_0 ));
    CascadeMux I__1155 (
            .O(N__8321),
            .I(\uart_inst0.tx_uart_fifo_inst.rDataCount_RNIJHQM1Z0Z_2_cascade_ ));
    InMux I__1154 (
            .O(N__8318),
            .I(N__8311));
    InMux I__1153 (
            .O(N__8317),
            .I(N__8308));
    InMux I__1152 (
            .O(N__8316),
            .I(N__8305));
    CascadeMux I__1151 (
            .O(N__8315),
            .I(N__8302));
    InMux I__1150 (
            .O(N__8314),
            .I(N__8297));
    LocalMux I__1149 (
            .O(N__8311),
            .I(N__8292));
    LocalMux I__1148 (
            .O(N__8308),
            .I(N__8292));
    LocalMux I__1147 (
            .O(N__8305),
            .I(N__8289));
    InMux I__1146 (
            .O(N__8302),
            .I(N__8286));
    InMux I__1145 (
            .O(N__8301),
            .I(N__8283));
    InMux I__1144 (
            .O(N__8300),
            .I(N__8280));
    LocalMux I__1143 (
            .O(N__8297),
            .I(\uart_inst0.tx_uart_fifo_inst.wUartTxFull ));
    Odrv4 I__1142 (
            .O(N__8292),
            .I(\uart_inst0.tx_uart_fifo_inst.wUartTxFull ));
    Odrv12 I__1141 (
            .O(N__8289),
            .I(\uart_inst0.tx_uart_fifo_inst.wUartTxFull ));
    LocalMux I__1140 (
            .O(N__8286),
            .I(\uart_inst0.tx_uart_fifo_inst.wUartTxFull ));
    LocalMux I__1139 (
            .O(N__8283),
            .I(\uart_inst0.tx_uart_fifo_inst.wUartTxFull ));
    LocalMux I__1138 (
            .O(N__8280),
            .I(\uart_inst0.tx_uart_fifo_inst.wUartTxFull ));
    InMux I__1137 (
            .O(N__8267),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_0 ));
    InMux I__1136 (
            .O(N__8264),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_1 ));
    InMux I__1135 (
            .O(N__8261),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_2 ));
    InMux I__1134 (
            .O(N__8258),
            .I(N__8253));
    InMux I__1133 (
            .O(N__8257),
            .I(N__8248));
    InMux I__1132 (
            .O(N__8256),
            .I(N__8248));
    LocalMux I__1131 (
            .O(N__8253),
            .I(N__8245));
    LocalMux I__1130 (
            .O(N__8248),
            .I(N__8240));
    Span4Mux_s2_v I__1129 (
            .O(N__8245),
            .I(N__8240));
    Odrv4 I__1128 (
            .O(N__8240),
            .I(fifo_inst_ft2232h_inst_rFifoState_3));
    InMux I__1127 (
            .O(N__8237),
            .I(N__8232));
    InMux I__1126 (
            .O(N__8236),
            .I(N__8227));
    InMux I__1125 (
            .O(N__8235),
            .I(N__8227));
    LocalMux I__1124 (
            .O(N__8232),
            .I(fifo_inst_rx_fifo_inst_un1_rDataCount15_2_0_0));
    LocalMux I__1123 (
            .O(N__8227),
            .I(fifo_inst_rx_fifo_inst_un1_rDataCount15_2_0_0));
    InMux I__1122 (
            .O(N__8222),
            .I(N__8217));
    InMux I__1121 (
            .O(N__8221),
            .I(N__8214));
    InMux I__1120 (
            .O(N__8220),
            .I(N__8211));
    LocalMux I__1119 (
            .O(N__8217),
            .I(fifo_inst_rx_fifo_inst_rDataCount_fast_0));
    LocalMux I__1118 (
            .O(N__8214),
            .I(fifo_inst_rx_fifo_inst_rDataCount_fast_0));
    LocalMux I__1117 (
            .O(N__8211),
            .I(fifo_inst_rx_fifo_inst_rDataCount_fast_0));
    InMux I__1116 (
            .O(N__8204),
            .I(N__8201));
    LocalMux I__1115 (
            .O(N__8201),
            .I(N__8196));
    InMux I__1114 (
            .O(N__8200),
            .I(N__8193));
    InMux I__1113 (
            .O(N__8199),
            .I(N__8190));
    Odrv4 I__1112 (
            .O(N__8196),
            .I(N_84_mux));
    LocalMux I__1111 (
            .O(N__8193),
            .I(N_84_mux));
    LocalMux I__1110 (
            .O(N__8190),
            .I(N_84_mux));
    CascadeMux I__1109 (
            .O(N__8183),
            .I(rUartTxEn_4_cascade_));
    CascadeMux I__1108 (
            .O(N__8180),
            .I(N__8176));
    InMux I__1107 (
            .O(N__8179),
            .I(N__8172));
    InMux I__1106 (
            .O(N__8176),
            .I(N__8167));
    InMux I__1105 (
            .O(N__8175),
            .I(N__8167));
    LocalMux I__1104 (
            .O(N__8172),
            .I(rFtdiRxStateZ0Z_0));
    LocalMux I__1103 (
            .O(N__8167),
            .I(rFtdiRxStateZ0Z_0));
    InMux I__1102 (
            .O(N__8162),
            .I(N__8159));
    LocalMux I__1101 (
            .O(N__8159),
            .I(N__8156));
    Span4Mux_s3_v I__1100 (
            .O(N__8156),
            .I(N__8153));
    Odrv4 I__1099 (
            .O(N__8153),
            .I(\fifo_inst.ft2232h_inst.rFifoStatesr_0 ));
    InMux I__1098 (
            .O(N__8150),
            .I(N__8147));
    LocalMux I__1097 (
            .O(N__8147),
            .I(N__8143));
    InMux I__1096 (
            .O(N__8146),
            .I(N__8140));
    Span4Mux_h I__1095 (
            .O(N__8143),
            .I(N__8137));
    LocalMux I__1094 (
            .O(N__8140),
            .I(N__8134));
    Span4Mux_v I__1093 (
            .O(N__8137),
            .I(N__8130));
    Span4Mux_h I__1092 (
            .O(N__8134),
            .I(N__8127));
    InMux I__1091 (
            .O(N__8133),
            .I(N__8124));
    Odrv4 I__1090 (
            .O(N__8130),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_2 ));
    Odrv4 I__1089 (
            .O(N__8127),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_2 ));
    LocalMux I__1088 (
            .O(N__8124),
            .I(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_2 ));
    InMux I__1087 (
            .O(N__8117),
            .I(N__8113));
    InMux I__1086 (
            .O(N__8116),
            .I(N__8110));
    LocalMux I__1085 (
            .O(N__8113),
            .I(N__8107));
    LocalMux I__1084 (
            .O(N__8110),
            .I(N__8104));
    Span4Mux_v I__1083 (
            .O(N__8107),
            .I(N__8098));
    Span4Mux_h I__1082 (
            .O(N__8104),
            .I(N__8098));
    InMux I__1081 (
            .O(N__8103),
            .I(N__8095));
    Span4Mux_v I__1080 (
            .O(N__8098),
            .I(N__8090));
    LocalMux I__1079 (
            .O(N__8095),
            .I(N__8090));
    Span4Mux_h I__1078 (
            .O(N__8090),
            .I(N__8087));
    Sp12to4 I__1077 (
            .O(N__8087),
            .I(N__8084));
    Span12Mux_v I__1076 (
            .O(N__8084),
            .I(N__8081));
    Odrv12 I__1075 (
            .O(N__8081),
            .I(iRxF_n_c));
    InMux I__1074 (
            .O(N__8078),
            .I(N__8074));
    InMux I__1073 (
            .O(N__8077),
            .I(N__8071));
    LocalMux I__1072 (
            .O(N__8074),
            .I(N__8068));
    LocalMux I__1071 (
            .O(N__8071),
            .I(N__8064));
    Span4Mux_h I__1070 (
            .O(N__8068),
            .I(N__8061));
    InMux I__1069 (
            .O(N__8067),
            .I(N__8058));
    Odrv12 I__1068 (
            .O(N__8064),
            .I(fifo_inst_ft2232h_inst_rFifoState_0));
    Odrv4 I__1067 (
            .O(N__8061),
            .I(fifo_inst_ft2232h_inst_rFifoState_0));
    LocalMux I__1066 (
            .O(N__8058),
            .I(fifo_inst_ft2232h_inst_rFifoState_0));
    CascadeMux I__1065 (
            .O(N__8051),
            .I(\fifo_inst.rx_fifo_inst.un1_rDataCount_axbxc3_1_1_cascade_ ));
    CascadeMux I__1064 (
            .O(N__8048),
            .I(\uart_inst0.tx_uart_fifo_inst.m15_xZ0Z0_cascade_ ));
    InMux I__1063 (
            .O(N__8045),
            .I(N__8042));
    LocalMux I__1062 (
            .O(N__8042),
            .I(\fifo_inst.rx_fifo_inst.un1_rDataCount_axbxc3_1_1 ));
    CascadeMux I__1061 (
            .O(N__8039),
            .I(N__8036));
    InMux I__1060 (
            .O(N__8036),
            .I(N__8031));
    InMux I__1059 (
            .O(N__8035),
            .I(N__8026));
    InMux I__1058 (
            .O(N__8034),
            .I(N__8026));
    LocalMux I__1057 (
            .O(N__8031),
            .I(fifo_inst_rx_fifo_inst_rDataCount_fast_3));
    LocalMux I__1056 (
            .O(N__8026),
            .I(fifo_inst_rx_fifo_inst_rDataCount_fast_3));
    IoInMux I__1055 (
            .O(N__8021),
            .I(N__8018));
    LocalMux I__1054 (
            .O(N__8018),
            .I(N__8015));
    IoSpan4Mux I__1053 (
            .O(N__8015),
            .I(N__8011));
    IoInMux I__1052 (
            .O(N__8014),
            .I(N__8008));
    Span4Mux_s0_v I__1051 (
            .O(N__8011),
            .I(N__8005));
    LocalMux I__1050 (
            .O(N__8008),
            .I(N__8002));
    Sp12to4 I__1049 (
            .O(N__8005),
            .I(N__7999));
    IoSpan4Mux I__1048 (
            .O(N__8002),
            .I(N__7996));
    Span12Mux_v I__1047 (
            .O(N__7999),
            .I(N__7993));
    Span4Mux_s3_v I__1046 (
            .O(N__7996),
            .I(N__7990));
    Span12Mux_v I__1045 (
            .O(N__7993),
            .I(N__7986));
    Span4Mux_h I__1044 (
            .O(N__7990),
            .I(N__7983));
    InMux I__1043 (
            .O(N__7989),
            .I(N__7980));
    Odrv12 I__1042 (
            .O(N__7986),
            .I(P1A4_c));
    Odrv4 I__1041 (
            .O(N__7983),
            .I(P1A4_c));
    LocalMux I__1040 (
            .O(N__7980),
            .I(P1A4_c));
    CascadeMux I__1039 (
            .O(N__7973),
            .I(\uart_inst0.tx_uart_fifo_inst.m8_xZ0Z0_cascade_ ));
    InMux I__1038 (
            .O(N__7970),
            .I(N__7967));
    LocalMux I__1037 (
            .O(N__7967),
            .I(N__7963));
    InMux I__1036 (
            .O(N__7966),
            .I(N__7960));
    Odrv4 I__1035 (
            .O(N__7963),
            .I(\fifo_inst.tx_fifo_inst.un1_rDataCount_axbxc3_2_tz ));
    LocalMux I__1034 (
            .O(N__7960),
            .I(\fifo_inst.tx_fifo_inst.un1_rDataCount_axbxc3_2_tz ));
    CascadeMux I__1033 (
            .O(N__7955),
            .I(N__7952));
    InMux I__1032 (
            .O(N__7952),
            .I(N__7948));
    CascadeMux I__1031 (
            .O(N__7951),
            .I(N__7945));
    LocalMux I__1030 (
            .O(N__7948),
            .I(N__7942));
    InMux I__1029 (
            .O(N__7945),
            .I(N__7939));
    Odrv4 I__1028 (
            .O(N__7942),
            .I(\fifo_inst.tx_fifo_inst.un1_rDataCount_axbxc3_a0_2 ));
    LocalMux I__1027 (
            .O(N__7939),
            .I(\fifo_inst.tx_fifo_inst.un1_rDataCount_axbxc3_a0_2 ));
    InMux I__1026 (
            .O(N__7934),
            .I(N__7931));
    LocalMux I__1025 (
            .O(N__7931),
            .I(\fifo_inst.tx_fifo_inst.un1_rDataCount_c2_0 ));
    CEMux I__1024 (
            .O(N__7928),
            .I(N__7924));
    InMux I__1023 (
            .O(N__7927),
            .I(N__7920));
    LocalMux I__1022 (
            .O(N__7924),
            .I(N__7915));
    CascadeMux I__1021 (
            .O(N__7923),
            .I(N__7912));
    LocalMux I__1020 (
            .O(N__7920),
            .I(N__7909));
    CascadeMux I__1019 (
            .O(N__7919),
            .I(N__7906));
    InMux I__1018 (
            .O(N__7918),
            .I(N__7903));
    Span4Mux_h I__1017 (
            .O(N__7915),
            .I(N__7900));
    InMux I__1016 (
            .O(N__7912),
            .I(N__7897));
    Span4Mux_v I__1015 (
            .O(N__7909),
            .I(N__7894));
    InMux I__1014 (
            .O(N__7906),
            .I(N__7891));
    LocalMux I__1013 (
            .O(N__7903),
            .I(N__7886));
    Span4Mux_h I__1012 (
            .O(N__7900),
            .I(N__7886));
    LocalMux I__1011 (
            .O(N__7897),
            .I(fifo_inst_tx_fifo_inst_wRamWrEn));
    Odrv4 I__1010 (
            .O(N__7894),
            .I(fifo_inst_tx_fifo_inst_wRamWrEn));
    LocalMux I__1009 (
            .O(N__7891),
            .I(fifo_inst_tx_fifo_inst_wRamWrEn));
    Odrv4 I__1008 (
            .O(N__7886),
            .I(fifo_inst_tx_fifo_inst_wRamWrEn));
    CascadeMux I__1007 (
            .O(N__7877),
            .I(N__7874));
    InMux I__1006 (
            .O(N__7874),
            .I(N__7870));
    InMux I__1005 (
            .O(N__7873),
            .I(N__7867));
    LocalMux I__1004 (
            .O(N__7870),
            .I(N__7863));
    LocalMux I__1003 (
            .O(N__7867),
            .I(N__7860));
    InMux I__1002 (
            .O(N__7866),
            .I(N__7857));
    Span4Mux_h I__1001 (
            .O(N__7863),
            .I(N__7854));
    Odrv4 I__1000 (
            .O(N__7860),
            .I(\fifo_inst.tx_fifo_inst.un1_rDataCount_ac0_1_a0_0 ));
    LocalMux I__999 (
            .O(N__7857),
            .I(\fifo_inst.tx_fifo_inst.un1_rDataCount_ac0_1_a0_0 ));
    Odrv4 I__998 (
            .O(N__7854),
            .I(\fifo_inst.tx_fifo_inst.un1_rDataCount_ac0_1_a0_0 ));
    CascadeMux I__997 (
            .O(N__7847),
            .I(\fifo_inst.tx_fifo_inst.un1_rDataCount_c2_1_cascade_ ));
    InMux I__996 (
            .O(N__7844),
            .I(N__7841));
    LocalMux I__995 (
            .O(N__7841),
            .I(\fifo_inst.tx_fifo_inst.un1_rDataCount_ac0_2 ));
    InMux I__994 (
            .O(N__7838),
            .I(N__7834));
    InMux I__993 (
            .O(N__7837),
            .I(N__7831));
    LocalMux I__992 (
            .O(N__7834),
            .I(fifo_inst_tx_fifo_inst_un1_rDataCount15_2_0_0));
    LocalMux I__991 (
            .O(N__7831),
            .I(fifo_inst_tx_fifo_inst_un1_rDataCount15_2_0_0));
    InMux I__990 (
            .O(N__7826),
            .I(N__7820));
    InMux I__989 (
            .O(N__7825),
            .I(N__7820));
    LocalMux I__988 (
            .O(N__7820),
            .I(N__7816));
    CascadeMux I__987 (
            .O(N__7819),
            .I(N__7810));
    Span4Mux_s3_v I__986 (
            .O(N__7816),
            .I(N__7807));
    InMux I__985 (
            .O(N__7815),
            .I(N__7804));
    InMux I__984 (
            .O(N__7814),
            .I(N__7799));
    InMux I__983 (
            .O(N__7813),
            .I(N__7799));
    InMux I__982 (
            .O(N__7810),
            .I(N__7796));
    Odrv4 I__981 (
            .O(N__7807),
            .I(fifo_inst_tx_fifo_inst_rDataCount_2));
    LocalMux I__980 (
            .O(N__7804),
            .I(fifo_inst_tx_fifo_inst_rDataCount_2));
    LocalMux I__979 (
            .O(N__7799),
            .I(fifo_inst_tx_fifo_inst_rDataCount_2));
    LocalMux I__978 (
            .O(N__7796),
            .I(fifo_inst_tx_fifo_inst_rDataCount_2));
    InMux I__977 (
            .O(N__7787),
            .I(N__7780));
    InMux I__976 (
            .O(N__7786),
            .I(N__7780));
    CascadeMux I__975 (
            .O(N__7785),
            .I(N__7777));
    LocalMux I__974 (
            .O(N__7780),
            .I(N__7774));
    InMux I__973 (
            .O(N__7777),
            .I(N__7766));
    Span4Mux_h I__972 (
            .O(N__7774),
            .I(N__7763));
    InMux I__971 (
            .O(N__7773),
            .I(N__7758));
    InMux I__970 (
            .O(N__7772),
            .I(N__7758));
    InMux I__969 (
            .O(N__7771),
            .I(N__7753));
    InMux I__968 (
            .O(N__7770),
            .I(N__7753));
    InMux I__967 (
            .O(N__7769),
            .I(N__7750));
    LocalMux I__966 (
            .O(N__7766),
            .I(fifo_inst_tx_fifo_inst_rDataCount_1));
    Odrv4 I__965 (
            .O(N__7763),
            .I(fifo_inst_tx_fifo_inst_rDataCount_1));
    LocalMux I__964 (
            .O(N__7758),
            .I(fifo_inst_tx_fifo_inst_rDataCount_1));
    LocalMux I__963 (
            .O(N__7753),
            .I(fifo_inst_tx_fifo_inst_rDataCount_1));
    LocalMux I__962 (
            .O(N__7750),
            .I(fifo_inst_tx_fifo_inst_rDataCount_1));
    CascadeMux I__961 (
            .O(N__7739),
            .I(N__7736));
    InMux I__960 (
            .O(N__7736),
            .I(N__7731));
    InMux I__959 (
            .O(N__7735),
            .I(N__7726));
    InMux I__958 (
            .O(N__7734),
            .I(N__7726));
    LocalMux I__957 (
            .O(N__7731),
            .I(fifo_inst_tx_fifo_inst_rDataCount_fast_3));
    LocalMux I__956 (
            .O(N__7726),
            .I(fifo_inst_tx_fifo_inst_rDataCount_fast_3));
    InMux I__955 (
            .O(N__7721),
            .I(N__7712));
    InMux I__954 (
            .O(N__7720),
            .I(N__7712));
    InMux I__953 (
            .O(N__7719),
            .I(N__7706));
    InMux I__952 (
            .O(N__7718),
            .I(N__7701));
    InMux I__951 (
            .O(N__7717),
            .I(N__7701));
    LocalMux I__950 (
            .O(N__7712),
            .I(N__7698));
    InMux I__949 (
            .O(N__7711),
            .I(N__7695));
    InMux I__948 (
            .O(N__7710),
            .I(N__7690));
    InMux I__947 (
            .O(N__7709),
            .I(N__7690));
    LocalMux I__946 (
            .O(N__7706),
            .I(fifo_inst_tx_fifo_inst_rDataCount_0));
    LocalMux I__945 (
            .O(N__7701),
            .I(fifo_inst_tx_fifo_inst_rDataCount_0));
    Odrv4 I__944 (
            .O(N__7698),
            .I(fifo_inst_tx_fifo_inst_rDataCount_0));
    LocalMux I__943 (
            .O(N__7695),
            .I(fifo_inst_tx_fifo_inst_rDataCount_0));
    LocalMux I__942 (
            .O(N__7690),
            .I(fifo_inst_tx_fifo_inst_rDataCount_0));
    InMux I__941 (
            .O(N__7679),
            .I(N__7676));
    LocalMux I__940 (
            .O(N__7676),
            .I(N__7673));
    Span4Mux_v I__939 (
            .O(N__7673),
            .I(N__7670));
    Odrv4 I__938 (
            .O(N__7670),
            .I(\uart_inst0.wTxRdData_4 ));
    InMux I__937 (
            .O(N__7667),
            .I(N__7664));
    LocalMux I__936 (
            .O(N__7664),
            .I(\uart_inst0.uart_inst0.rTxDataZ0Z_4 ));
    InMux I__935 (
            .O(N__7661),
            .I(N__7658));
    LocalMux I__934 (
            .O(N__7658),
            .I(\uart_inst0.uart_inst0.rTxDataZ0Z_3 ));
    InMux I__933 (
            .O(N__7655),
            .I(N__7652));
    LocalMux I__932 (
            .O(N__7652),
            .I(N__7649));
    Odrv12 I__931 (
            .O(N__7649),
            .I(\uart_inst0.wTxRdData_2 ));
    InMux I__930 (
            .O(N__7646),
            .I(N__7643));
    LocalMux I__929 (
            .O(N__7643),
            .I(\uart_inst0.uart_inst0.rTxDataZ0Z_2 ));
    InMux I__928 (
            .O(N__7640),
            .I(N__7637));
    LocalMux I__927 (
            .O(N__7637),
            .I(\uart_inst0.uart_inst0.rTxDataZ0Z_6 ));
    InMux I__926 (
            .O(N__7634),
            .I(N__7631));
    LocalMux I__925 (
            .O(N__7631),
            .I(N__7628));
    Odrv12 I__924 (
            .O(N__7628),
            .I(\uart_inst0.wTxRdData_5 ));
    InMux I__923 (
            .O(N__7625),
            .I(N__7622));
    LocalMux I__922 (
            .O(N__7622),
            .I(\uart_inst0.uart_inst0.rTxDataZ0Z_5 ));
    InMux I__921 (
            .O(N__7619),
            .I(N__7616));
    LocalMux I__920 (
            .O(N__7616),
            .I(N__7613));
    Odrv12 I__919 (
            .O(N__7613),
            .I(\uart_inst0.wTxRdData_7 ));
    CascadeMux I__918 (
            .O(N__7610),
            .I(N__7607));
    InMux I__917 (
            .O(N__7607),
            .I(N__7603));
    InMux I__916 (
            .O(N__7606),
            .I(N__7600));
    LocalMux I__915 (
            .O(N__7603),
            .I(\uart_inst0.uart_inst0.rTxDataZ0Z_7 ));
    LocalMux I__914 (
            .O(N__7600),
            .I(\uart_inst0.uart_inst0.rTxDataZ0Z_7 ));
    CascadeMux I__913 (
            .O(N__7595),
            .I(N_97_cascade_));
    InMux I__912 (
            .O(N__7592),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_3 ));
    InMux I__911 (
            .O(N__7589),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_4 ));
    InMux I__910 (
            .O(N__7586),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_5 ));
    InMux I__909 (
            .O(N__7583),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_6 ));
    InMux I__908 (
            .O(N__7580),
            .I(bfn_13_13_0_));
    CascadeMux I__907 (
            .O(N__7577),
            .I(N__7574));
    InMux I__906 (
            .O(N__7574),
            .I(N__7571));
    LocalMux I__905 (
            .O(N__7571),
            .I(N__7568));
    Span4Mux_v I__904 (
            .O(N__7568),
            .I(N__7564));
    InMux I__903 (
            .O(N__7567),
            .I(N__7560));
    Span4Mux_h I__902 (
            .O(N__7564),
            .I(N__7557));
    InMux I__901 (
            .O(N__7563),
            .I(N__7554));
    LocalMux I__900 (
            .O(N__7560),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_8 ));
    Odrv4 I__899 (
            .O(N__7557),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_8 ));
    LocalMux I__898 (
            .O(N__7554),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_8 ));
    InMux I__897 (
            .O(N__7547),
            .I(N__7544));
    LocalMux I__896 (
            .O(N__7544),
            .I(N__7541));
    Odrv12 I__895 (
            .O(N__7541),
            .I(\uart_inst0.wTxRdData_0 ));
    InMux I__894 (
            .O(N__7538),
            .I(N__7535));
    LocalMux I__893 (
            .O(N__7535),
            .I(N__7532));
    Odrv12 I__892 (
            .O(N__7532),
            .I(\uart_inst0.wTxRdData_1 ));
    InMux I__891 (
            .O(N__7529),
            .I(N__7526));
    LocalMux I__890 (
            .O(N__7526),
            .I(\uart_inst0.uart_inst0.rTxDataZ0Z_1 ));
    InMux I__889 (
            .O(N__7523),
            .I(N__7520));
    LocalMux I__888 (
            .O(N__7520),
            .I(N__7517));
    Odrv12 I__887 (
            .O(N__7517),
            .I(\uart_inst0.wTxRdData_6 ));
    InMux I__886 (
            .O(N__7514),
            .I(N__7511));
    LocalMux I__885 (
            .O(N__7511),
            .I(N__7508));
    Odrv12 I__884 (
            .O(N__7508),
            .I(\uart_inst0.wTxRdData_3 ));
    InMux I__883 (
            .O(N__7505),
            .I(N__7502));
    LocalMux I__882 (
            .O(N__7502),
            .I(N__7499));
    Span4Mux_v I__881 (
            .O(N__7499),
            .I(N__7496));
    Span4Mux_h I__880 (
            .O(N__7496),
            .I(N__7493));
    Odrv4 I__879 (
            .O(N__7493),
            .I(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_3 ));
    InMux I__878 (
            .O(N__7490),
            .I(N__7487));
    LocalMux I__877 (
            .O(N__7487),
            .I(N__7484));
    Span4Mux_h I__876 (
            .O(N__7484),
            .I(N__7481));
    Odrv4 I__875 (
            .O(N__7481),
            .I(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_4 ));
    InMux I__874 (
            .O(N__7478),
            .I(N__7475));
    LocalMux I__873 (
            .O(N__7475),
            .I(N__7472));
    Span4Mux_h I__872 (
            .O(N__7472),
            .I(N__7469));
    Odrv4 I__871 (
            .O(N__7469),
            .I(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_5 ));
    InMux I__870 (
            .O(N__7466),
            .I(N__7463));
    LocalMux I__869 (
            .O(N__7463),
            .I(N__7460));
    Odrv12 I__868 (
            .O(N__7460),
            .I(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_6 ));
    InMux I__867 (
            .O(N__7457),
            .I(N__7454));
    LocalMux I__866 (
            .O(N__7454),
            .I(N__7451));
    Span4Mux_h I__865 (
            .O(N__7451),
            .I(N__7448));
    Odrv4 I__864 (
            .O(N__7448),
            .I(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_7 ));
    CascadeMux I__863 (
            .O(N__7445),
            .I(N__7442));
    InMux I__862 (
            .O(N__7442),
            .I(N__7439));
    LocalMux I__861 (
            .O(N__7439),
            .I(N__7436));
    Span4Mux_h I__860 (
            .O(N__7436),
            .I(N__7432));
    InMux I__859 (
            .O(N__7435),
            .I(N__7428));
    Span4Mux_h I__858 (
            .O(N__7432),
            .I(N__7425));
    InMux I__857 (
            .O(N__7431),
            .I(N__7422));
    LocalMux I__856 (
            .O(N__7428),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ1Z_0 ));
    Odrv4 I__855 (
            .O(N__7425),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ1Z_0 ));
    LocalMux I__854 (
            .O(N__7422),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ1Z_0 ));
    InMux I__853 (
            .O(N__7415),
            .I(N__7412));
    LocalMux I__852 (
            .O(N__7412),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNO_0Z0Z_0 ));
    CascadeMux I__851 (
            .O(N__7409),
            .I(N__7406));
    InMux I__850 (
            .O(N__7406),
            .I(N__7402));
    InMux I__849 (
            .O(N__7405),
            .I(N__7398));
    LocalMux I__848 (
            .O(N__7402),
            .I(N__7395));
    InMux I__847 (
            .O(N__7401),
            .I(N__7392));
    LocalMux I__846 (
            .O(N__7398),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ1Z_1 ));
    Odrv12 I__845 (
            .O(N__7395),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ1Z_1 ));
    LocalMux I__844 (
            .O(N__7392),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ1Z_1 ));
    InMux I__843 (
            .O(N__7385),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_0 ));
    CascadeMux I__842 (
            .O(N__7382),
            .I(N__7379));
    InMux I__841 (
            .O(N__7379),
            .I(N__7376));
    LocalMux I__840 (
            .O(N__7376),
            .I(N__7372));
    InMux I__839 (
            .O(N__7375),
            .I(N__7368));
    Span4Mux_h I__838 (
            .O(N__7372),
            .I(N__7365));
    InMux I__837 (
            .O(N__7371),
            .I(N__7362));
    LocalMux I__836 (
            .O(N__7368),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ0Z_2 ));
    Odrv4 I__835 (
            .O(N__7365),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ0Z_2 ));
    LocalMux I__834 (
            .O(N__7362),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ0Z_2 ));
    InMux I__833 (
            .O(N__7355),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_1 ));
    CascadeMux I__832 (
            .O(N__7352),
            .I(N__7349));
    InMux I__831 (
            .O(N__7349),
            .I(N__7346));
    LocalMux I__830 (
            .O(N__7346),
            .I(N__7343));
    Span4Mux_h I__829 (
            .O(N__7343),
            .I(N__7340));
    Span4Mux_h I__828 (
            .O(N__7340),
            .I(N__7335));
    InMux I__827 (
            .O(N__7339),
            .I(N__7332));
    InMux I__826 (
            .O(N__7338),
            .I(N__7329));
    Odrv4 I__825 (
            .O(N__7335),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_3 ));
    LocalMux I__824 (
            .O(N__7332),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_3 ));
    LocalMux I__823 (
            .O(N__7329),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_3 ));
    InMux I__822 (
            .O(N__7322),
            .I(N__7319));
    LocalMux I__821 (
            .O(N__7319),
            .I(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNO_0Z0Z_3 ));
    InMux I__820 (
            .O(N__7316),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_2 ));
    InMux I__819 (
            .O(N__7313),
            .I(N__7310));
    LocalMux I__818 (
            .O(N__7310),
            .I(N__7306));
    InMux I__817 (
            .O(N__7309),
            .I(N__7303));
    Odrv4 I__816 (
            .O(N__7306),
            .I(rUartTxEnZ0));
    LocalMux I__815 (
            .O(N__7303),
            .I(rUartTxEnZ0));
    InMux I__814 (
            .O(N__7298),
            .I(N__7295));
    LocalMux I__813 (
            .O(N__7295),
            .I(N__7292));
    Span4Mux_v I__812 (
            .O(N__7292),
            .I(N__7289));
    Odrv4 I__811 (
            .O(N__7289),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c3_0_0 ));
    CascadeMux I__810 (
            .O(N__7286),
            .I(N__7283));
    InMux I__809 (
            .O(N__7283),
            .I(N__7280));
    LocalMux I__808 (
            .O(N__7280),
            .I(N__7277));
    Span4Mux_v I__807 (
            .O(N__7277),
            .I(N__7274));
    Odrv4 I__806 (
            .O(N__7274),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c2_d ));
    InMux I__805 (
            .O(N__7271),
            .I(N__7267));
    InMux I__804 (
            .O(N__7270),
            .I(N__7264));
    LocalMux I__803 (
            .O(N__7267),
            .I(N__7258));
    LocalMux I__802 (
            .O(N__7264),
            .I(N__7258));
    InMux I__801 (
            .O(N__7263),
            .I(N__7255));
    Odrv12 I__800 (
            .O(N__7258),
            .I(\uart_inst0.tx_uart_fifo_inst.rDataCount_0_sqmuxa ));
    LocalMux I__799 (
            .O(N__7255),
            .I(\uart_inst0.tx_uart_fifo_inst.rDataCount_0_sqmuxa ));
    CascadeMux I__798 (
            .O(N__7250),
            .I(\uart_inst0.wTxRdEmpty_cascade_ ));
    InMux I__797 (
            .O(N__7247),
            .I(N__7244));
    LocalMux I__796 (
            .O(N__7244),
            .I(N__7241));
    Span4Mux_h I__795 (
            .O(N__7241),
            .I(N__7238));
    Span4Mux_h I__794 (
            .O(N__7238),
            .I(N__7235));
    Odrv4 I__793 (
            .O(N__7235),
            .I(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_0 ));
    InMux I__792 (
            .O(N__7232),
            .I(N__7229));
    LocalMux I__791 (
            .O(N__7229),
            .I(N__7226));
    Span4Mux_h I__790 (
            .O(N__7226),
            .I(N__7223));
    Span4Mux_h I__789 (
            .O(N__7223),
            .I(N__7220));
    Odrv4 I__788 (
            .O(N__7220),
            .I(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_1 ));
    InMux I__787 (
            .O(N__7217),
            .I(N__7214));
    LocalMux I__786 (
            .O(N__7214),
            .I(N__7211));
    Span12Mux_h I__785 (
            .O(N__7211),
            .I(N__7208));
    Odrv12 I__784 (
            .O(N__7208),
            .I(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_2 ));
    CascadeMux I__783 (
            .O(N__7205),
            .I(\uart_inst0.tx_uart_fifo_inst.m65_bmZ0_cascade_ ));
    CascadeMux I__782 (
            .O(N__7202),
            .I(\fifo_inst.rx_fifo_inst.un1_rDataCount_c2_1_1_0_cascade_ ));
    InMux I__781 (
            .O(N__7199),
            .I(N__7196));
    LocalMux I__780 (
            .O(N__7196),
            .I(\uart_inst0.tx_uart_fifo_inst.m65_nsZ0Z_1 ));
    InMux I__779 (
            .O(N__7193),
            .I(N__7190));
    LocalMux I__778 (
            .O(N__7190),
            .I(\fifo_inst.rx_fifo_inst.un1_rDataCount_c2_1 ));
    CascadeMux I__777 (
            .O(N__7187),
            .I(N__7184));
    InMux I__776 (
            .O(N__7184),
            .I(N__7178));
    InMux I__775 (
            .O(N__7183),
            .I(N__7178));
    LocalMux I__774 (
            .O(N__7178),
            .I(fifo_inst_rx_fifo_inst_rDataCount_0_sqmuxa));
    CascadeMux I__773 (
            .O(N__7175),
            .I(N__7172));
    InMux I__772 (
            .O(N__7172),
            .I(N__7169));
    LocalMux I__771 (
            .O(N__7169),
            .I(\fifo_inst.rx_fifo_inst.un1_rDataCount_ac0_2 ));
    InMux I__770 (
            .O(N__7166),
            .I(N__7163));
    LocalMux I__769 (
            .O(N__7163),
            .I(\uart_inst0.tx_uart_fifo_inst.m78_bmZ0 ));
    CascadeMux I__768 (
            .O(N__7160),
            .I(\uart_inst0.tx_uart_fifo_inst.m78_nsZ0Z_1_cascade_ ));
    CEMux I__767 (
            .O(N__7157),
            .I(N__7154));
    LocalMux I__766 (
            .O(N__7154),
            .I(N__7151));
    Odrv4 I__765 (
            .O(N__7151),
            .I(\fifo_inst.ft2232h_inst.un1_rFifoState_12_0_i_0 ));
    CascadeMux I__764 (
            .O(N__7148),
            .I(\uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c2_d_cascade_ ));
    CascadeMux I__763 (
            .O(N__7145),
            .I(N_84_mux_cascade_));
    CascadeMux I__762 (
            .O(N__7142),
            .I(N__7139));
    InMux I__761 (
            .O(N__7139),
            .I(N__7136));
    LocalMux I__760 (
            .O(N__7136),
            .I(N__7132));
    InMux I__759 (
            .O(N__7135),
            .I(N__7128));
    Span4Mux_h I__758 (
            .O(N__7132),
            .I(N__7125));
    InMux I__757 (
            .O(N__7131),
            .I(N__7122));
    LocalMux I__756 (
            .O(N__7128),
            .I(N__7119));
    Odrv4 I__755 (
            .O(N__7125),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_5));
    LocalMux I__754 (
            .O(N__7122),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_5));
    Odrv4 I__753 (
            .O(N__7119),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_5));
    InMux I__752 (
            .O(N__7112),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_4 ));
    CascadeMux I__751 (
            .O(N__7109),
            .I(N__7106));
    InMux I__750 (
            .O(N__7106),
            .I(N__7103));
    LocalMux I__749 (
            .O(N__7103),
            .I(N__7098));
    InMux I__748 (
            .O(N__7102),
            .I(N__7095));
    InMux I__747 (
            .O(N__7101),
            .I(N__7092));
    Odrv12 I__746 (
            .O(N__7098),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_6));
    LocalMux I__745 (
            .O(N__7095),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_6));
    LocalMux I__744 (
            .O(N__7092),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_6));
    InMux I__743 (
            .O(N__7085),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_5 ));
    CascadeMux I__742 (
            .O(N__7082),
            .I(N__7079));
    InMux I__741 (
            .O(N__7079),
            .I(N__7075));
    InMux I__740 (
            .O(N__7078),
            .I(N__7071));
    LocalMux I__739 (
            .O(N__7075),
            .I(N__7068));
    InMux I__738 (
            .O(N__7074),
            .I(N__7065));
    LocalMux I__737 (
            .O(N__7071),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_7));
    Odrv12 I__736 (
            .O(N__7068),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_7));
    LocalMux I__735 (
            .O(N__7065),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_7));
    InMux I__734 (
            .O(N__7058),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_6 ));
    InMux I__733 (
            .O(N__7055),
            .I(bfn_13_3_0_));
    CascadeMux I__732 (
            .O(N__7052),
            .I(N__7049));
    InMux I__731 (
            .O(N__7049),
            .I(N__7046));
    LocalMux I__730 (
            .O(N__7046),
            .I(N__7042));
    CascadeMux I__729 (
            .O(N__7045),
            .I(N__7039));
    Span4Mux_s2_v I__728 (
            .O(N__7042),
            .I(N__7035));
    InMux I__727 (
            .O(N__7039),
            .I(N__7032));
    InMux I__726 (
            .O(N__7038),
            .I(N__7029));
    Span4Mux_h I__725 (
            .O(N__7035),
            .I(N__7026));
    LocalMux I__724 (
            .O(N__7032),
            .I(N__7023));
    LocalMux I__723 (
            .O(N__7029),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_8));
    Odrv4 I__722 (
            .O(N__7026),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_8));
    Odrv4 I__721 (
            .O(N__7023),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_8));
    CascadeMux I__720 (
            .O(N__7016),
            .I(fifo_inst_ft2232h_inst_un1_rFifoState_12_0_i_cascade_));
    CascadeMux I__719 (
            .O(N__7013),
            .I(N__7010));
    InMux I__718 (
            .O(N__7010),
            .I(N__7007));
    LocalMux I__717 (
            .O(N__7007),
            .I(\fifo_inst.tx_fifo_inst.un1_rDataCount_ac0_1_a1_1 ));
    CascadeMux I__716 (
            .O(N__7004),
            .I(\uart_inst0.tx_uart_fifo_inst.m68_eZ0Z_5_cascade_ ));
    InMux I__715 (
            .O(N__7001),
            .I(N__6998));
    LocalMux I__714 (
            .O(N__6998),
            .I(\uart_inst0.tx_uart_fifo_inst.m68_eZ0Z_6 ));
    InMux I__713 (
            .O(N__6995),
            .I(N__6991));
    InMux I__712 (
            .O(N__6994),
            .I(N__6988));
    LocalMux I__711 (
            .O(N__6991),
            .I(\uart_inst0.tx_uart_fifo_inst.N_92 ));
    LocalMux I__710 (
            .O(N__6988),
            .I(\uart_inst0.tx_uart_fifo_inst.N_92 ));
    CascadeMux I__709 (
            .O(N__6983),
            .I(N__6980));
    InMux I__708 (
            .O(N__6980),
            .I(N__6977));
    LocalMux I__707 (
            .O(N__6977),
            .I(N__6974));
    Span4Mux_v I__706 (
            .O(N__6974),
            .I(N__6971));
    Span4Mux_h I__705 (
            .O(N__6971),
            .I(N__6966));
    InMux I__704 (
            .O(N__6970),
            .I(N__6963));
    InMux I__703 (
            .O(N__6969),
            .I(N__6960));
    Odrv4 I__702 (
            .O(N__6966),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_0));
    LocalMux I__701 (
            .O(N__6963),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_0));
    LocalMux I__700 (
            .O(N__6960),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_0));
    InMux I__699 (
            .O(N__6953),
            .I(N__6950));
    LocalMux I__698 (
            .O(N__6950),
            .I(rRamWrAddr_RNI10581_0));
    CascadeMux I__697 (
            .O(N__6947),
            .I(N__6944));
    InMux I__696 (
            .O(N__6944),
            .I(N__6941));
    LocalMux I__695 (
            .O(N__6941),
            .I(N__6936));
    InMux I__694 (
            .O(N__6940),
            .I(N__6933));
    InMux I__693 (
            .O(N__6939),
            .I(N__6930));
    Odrv12 I__692 (
            .O(N__6936),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_1));
    LocalMux I__691 (
            .O(N__6933),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_1));
    LocalMux I__690 (
            .O(N__6930),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_1));
    InMux I__689 (
            .O(N__6923),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_0 ));
    CascadeMux I__688 (
            .O(N__6920),
            .I(N__6917));
    InMux I__687 (
            .O(N__6917),
            .I(N__6914));
    LocalMux I__686 (
            .O(N__6914),
            .I(N__6911));
    Span4Mux_h I__685 (
            .O(N__6911),
            .I(N__6906));
    InMux I__684 (
            .O(N__6910),
            .I(N__6903));
    InMux I__683 (
            .O(N__6909),
            .I(N__6900));
    Odrv4 I__682 (
            .O(N__6906),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_2));
    LocalMux I__681 (
            .O(N__6903),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_2));
    LocalMux I__680 (
            .O(N__6900),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_2));
    InMux I__679 (
            .O(N__6893),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_1 ));
    CascadeMux I__678 (
            .O(N__6890),
            .I(N__6887));
    InMux I__677 (
            .O(N__6887),
            .I(N__6884));
    LocalMux I__676 (
            .O(N__6884),
            .I(N__6881));
    Span12Mux_v I__675 (
            .O(N__6881),
            .I(N__6876));
    InMux I__674 (
            .O(N__6880),
            .I(N__6873));
    InMux I__673 (
            .O(N__6879),
            .I(N__6870));
    Odrv12 I__672 (
            .O(N__6876),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_3));
    LocalMux I__671 (
            .O(N__6873),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_3));
    LocalMux I__670 (
            .O(N__6870),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_3));
    InMux I__669 (
            .O(N__6863),
            .I(N__6860));
    LocalMux I__668 (
            .O(N__6860),
            .I(un1_rRamWrAddr_cry_2_c_RNISJKU));
    InMux I__667 (
            .O(N__6857),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_2 ));
    CascadeMux I__666 (
            .O(N__6854),
            .I(N__6851));
    InMux I__665 (
            .O(N__6851),
            .I(N__6847));
    CascadeMux I__664 (
            .O(N__6850),
            .I(N__6844));
    LocalMux I__663 (
            .O(N__6847),
            .I(N__6840));
    InMux I__662 (
            .O(N__6844),
            .I(N__6837));
    InMux I__661 (
            .O(N__6843),
            .I(N__6834));
    Span12Mux_s1_v I__660 (
            .O(N__6840),
            .I(N__6829));
    LocalMux I__659 (
            .O(N__6837),
            .I(N__6829));
    LocalMux I__658 (
            .O(N__6834),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_4));
    Odrv12 I__657 (
            .O(N__6829),
            .I(fifo_inst_tx_fifo_inst_rRamWrAddr_4));
    InMux I__656 (
            .O(N__6824),
            .I(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_3 ));
    IoInMux I__655 (
            .O(N__6821),
            .I(N__6817));
    IoInMux I__654 (
            .O(N__6820),
            .I(N__6814));
    LocalMux I__653 (
            .O(N__6817),
            .I(N__6811));
    LocalMux I__652 (
            .O(N__6814),
            .I(N__6808));
    Span4Mux_s3_v I__651 (
            .O(N__6811),
            .I(N__6805));
    Span4Mux_s1_v I__650 (
            .O(N__6808),
            .I(N__6802));
    Span4Mux_h I__649 (
            .O(N__6805),
            .I(N__6798));
    Span4Mux_h I__648 (
            .O(N__6802),
            .I(N__6795));
    InMux I__647 (
            .O(N__6801),
            .I(N__6792));
    Odrv4 I__646 (
            .O(N__6798),
            .I(P1A3_c));
    Odrv4 I__645 (
            .O(N__6795),
            .I(P1A3_c));
    LocalMux I__644 (
            .O(N__6792),
            .I(P1A3_c));
    InMux I__643 (
            .O(N__6785),
            .I(N__6782));
    LocalMux I__642 (
            .O(N__6782),
            .I(N_86_mux));
    CascadeMux I__641 (
            .O(N__6779),
            .I(\uart_inst0.tx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_0_cascade_ ));
    InMux I__640 (
            .O(N__6776),
            .I(N__6772));
    InMux I__639 (
            .O(N__6775),
            .I(N__6769));
    LocalMux I__638 (
            .O(N__6772),
            .I(\uart_inst0.tx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_6 ));
    LocalMux I__637 (
            .O(N__6769),
            .I(\uart_inst0.tx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_6 ));
    IoInMux I__636 (
            .O(N__6764),
            .I(N__6761));
    LocalMux I__635 (
            .O(N__6761),
            .I(GB_BUFFER_wPllLocked_i_g_THRU_CO));
    CascadeMux I__634 (
            .O(N__6758),
            .I(fifo_inst_tx_fifo_inst_wRamWrEn_cascade_));
    InMux I__633 (
            .O(N__6755),
            .I(N__6752));
    LocalMux I__632 (
            .O(N__6752),
            .I(\uart_inst0.uart_inst0.un1_rx_clk_divider_10 ));
    InMux I__631 (
            .O(N__6749),
            .I(N__6746));
    LocalMux I__630 (
            .O(N__6746),
            .I(\uart_inst0.uart_inst0.un1_rx_clk_divider_9 ));
    CascadeMux I__629 (
            .O(N__6743),
            .I(\uart_inst0.uart_inst0.un1_rx_clk_divider_7_cascade_ ));
    CascadeMux I__628 (
            .O(N__6740),
            .I(\uart_inst0.uart_inst0.un1_rx_clk_divider_0_cascade_ ));
    InMux I__627 (
            .O(N__6737),
            .I(N__6733));
    InMux I__626 (
            .O(N__6736),
            .I(N__6730));
    LocalMux I__625 (
            .O(N__6733),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_3 ));
    LocalMux I__624 (
            .O(N__6730),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_3 ));
    InMux I__623 (
            .O(N__6725),
            .I(N__6721));
    InMux I__622 (
            .O(N__6724),
            .I(N__6718));
    LocalMux I__621 (
            .O(N__6721),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_1 ));
    LocalMux I__620 (
            .O(N__6718),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_1 ));
    CascadeMux I__619 (
            .O(N__6713),
            .I(N__6709));
    InMux I__618 (
            .O(N__6712),
            .I(N__6706));
    InMux I__617 (
            .O(N__6709),
            .I(N__6703));
    LocalMux I__616 (
            .O(N__6706),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_4 ));
    LocalMux I__615 (
            .O(N__6703),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_4 ));
    InMux I__614 (
            .O(N__6698),
            .I(N__6694));
    InMux I__613 (
            .O(N__6697),
            .I(N__6691));
    LocalMux I__612 (
            .O(N__6694),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_2 ));
    LocalMux I__611 (
            .O(N__6691),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_2 ));
    InMux I__610 (
            .O(N__6686),
            .I(N__6683));
    LocalMux I__609 (
            .O(N__6683),
            .I(\uart_inst0.uart_inst0.un1_rx_clk_divider_8 ));
    InMux I__608 (
            .O(N__6680),
            .I(N__6675));
    InMux I__607 (
            .O(N__6679),
            .I(N__6672));
    InMux I__606 (
            .O(N__6678),
            .I(N__6669));
    LocalMux I__605 (
            .O(N__6675),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_0 ));
    LocalMux I__604 (
            .O(N__6672),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_0 ));
    LocalMux I__603 (
            .O(N__6669),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_0 ));
    SRMux I__602 (
            .O(N__6662),
            .I(N__6657));
    SRMux I__601 (
            .O(N__6661),
            .I(N__6654));
    SRMux I__600 (
            .O(N__6660),
            .I(N__6651));
    LocalMux I__599 (
            .O(N__6657),
            .I(\uart_inst0.uart_inst0.rx_clk_divider_1_sqmuxa_i ));
    LocalMux I__598 (
            .O(N__6654),
            .I(\uart_inst0.uart_inst0.rx_clk_divider_1_sqmuxa_i ));
    LocalMux I__597 (
            .O(N__6651),
            .I(\uart_inst0.uart_inst0.rx_clk_divider_1_sqmuxa_i ));
    InMux I__596 (
            .O(N__6644),
            .I(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_8 ));
    InMux I__595 (
            .O(N__6641),
            .I(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_9 ));
    InMux I__594 (
            .O(N__6638),
            .I(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_10 ));
    InMux I__593 (
            .O(N__6635),
            .I(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_11 ));
    InMux I__592 (
            .O(N__6632),
            .I(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_12 ));
    InMux I__591 (
            .O(N__6629),
            .I(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_13 ));
    InMux I__590 (
            .O(N__6626),
            .I(N__6622));
    InMux I__589 (
            .O(N__6625),
            .I(N__6619));
    LocalMux I__588 (
            .O(N__6622),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_8 ));
    LocalMux I__587 (
            .O(N__6619),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_8 ));
    InMux I__586 (
            .O(N__6614),
            .I(N__6610));
    InMux I__585 (
            .O(N__6613),
            .I(N__6607));
    LocalMux I__584 (
            .O(N__6610),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_7 ));
    LocalMux I__583 (
            .O(N__6607),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_7 ));
    CascadeMux I__582 (
            .O(N__6602),
            .I(N__6598));
    InMux I__581 (
            .O(N__6601),
            .I(N__6595));
    InMux I__580 (
            .O(N__6598),
            .I(N__6592));
    LocalMux I__579 (
            .O(N__6595),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_14 ));
    LocalMux I__578 (
            .O(N__6592),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_14 ));
    InMux I__577 (
            .O(N__6587),
            .I(N__6583));
    InMux I__576 (
            .O(N__6586),
            .I(N__6580));
    LocalMux I__575 (
            .O(N__6583),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_10 ));
    LocalMux I__574 (
            .O(N__6580),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_10 ));
    CascadeMux I__573 (
            .O(N__6575),
            .I(N__6572));
    InMux I__572 (
            .O(N__6572),
            .I(N__6568));
    InMux I__571 (
            .O(N__6571),
            .I(N__6565));
    LocalMux I__570 (
            .O(N__6568),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_11 ));
    LocalMux I__569 (
            .O(N__6565),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_11 ));
    CascadeMux I__568 (
            .O(N__6560),
            .I(N__6556));
    InMux I__567 (
            .O(N__6559),
            .I(N__6553));
    InMux I__566 (
            .O(N__6556),
            .I(N__6550));
    LocalMux I__565 (
            .O(N__6553),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_12 ));
    LocalMux I__564 (
            .O(N__6550),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_12 ));
    CascadeMux I__563 (
            .O(N__6545),
            .I(N__6542));
    InMux I__562 (
            .O(N__6542),
            .I(N__6538));
    InMux I__561 (
            .O(N__6541),
            .I(N__6535));
    LocalMux I__560 (
            .O(N__6538),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_9 ));
    LocalMux I__559 (
            .O(N__6535),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_9 ));
    CascadeMux I__558 (
            .O(N__6530),
            .I(N__6527));
    InMux I__557 (
            .O(N__6527),
            .I(N__6523));
    InMux I__556 (
            .O(N__6526),
            .I(N__6520));
    LocalMux I__555 (
            .O(N__6523),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_13 ));
    LocalMux I__554 (
            .O(N__6520),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_13 ));
    InMux I__553 (
            .O(N__6515),
            .I(N__6511));
    InMux I__552 (
            .O(N__6514),
            .I(N__6508));
    LocalMux I__551 (
            .O(N__6511),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_6 ));
    LocalMux I__550 (
            .O(N__6508),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_6 ));
    InMux I__549 (
            .O(N__6503),
            .I(N__6499));
    InMux I__548 (
            .O(N__6502),
            .I(N__6496));
    LocalMux I__547 (
            .O(N__6499),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_5 ));
    LocalMux I__546 (
            .O(N__6496),
            .I(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_5 ));
    InMux I__545 (
            .O(N__6491),
            .I(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_0 ));
    InMux I__544 (
            .O(N__6488),
            .I(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_1 ));
    InMux I__543 (
            .O(N__6485),
            .I(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_2 ));
    InMux I__542 (
            .O(N__6482),
            .I(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_3 ));
    InMux I__541 (
            .O(N__6479),
            .I(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_4 ));
    InMux I__540 (
            .O(N__6476),
            .I(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_5 ));
    InMux I__539 (
            .O(N__6473),
            .I(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_6 ));
    InMux I__538 (
            .O(N__6470),
            .I(bfn_9_15_0_));
    InMux I__537 (
            .O(N__6467),
            .I(N__6464));
    LocalMux I__536 (
            .O(N__6464),
            .I(\PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_CO ));
    IoInMux I__535 (
            .O(N__6461),
            .I(N__6458));
    LocalMux I__534 (
            .O(N__6458),
            .I(N__6455));
    Span12Mux_s9_v I__533 (
            .O(N__6455),
            .I(N__6452));
    Span12Mux_v I__532 (
            .O(N__6452),
            .I(N__6449));
    Odrv12 I__531 (
            .O(N__6449),
            .I(BTN_N_c));
    INV \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_0C  (
            .O(\INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net ),
            .I(N__16957));
    INV \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_5C  (
            .O(\INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_5C_net ),
            .I(N__16963));
    INV \INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7C  (
            .O(\INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7C_net ),
            .I(N__16980));
    INV \INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_4C  (
            .O(\INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_4C_net ),
            .I(N__16983));
    INV \INVfifo_inst.tx_fifo_inst.ram512x8_inst.RDATA_0C  (
            .O(\INVfifo_inst.tx_fifo_inst.ram512x8_inst.RDATA_0C_net ),
            .I(N__16977));
    INV \INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0C  (
            .O(\INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net ),
            .I(N__16924));
    INV \INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN  (
            .O(\INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net ),
            .I(N__16964));
    INV \INVfifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN  (
            .O(\INVfifo_inst.rx_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net ),
            .I(N__16986));
    INV \INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN  (
            .O(\INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net ),
            .I(N__16951));
    INV \INVfifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN  (
            .O(\INVfifo_inst.tx_fifo_inst.ram512x8_inst.mem_mem_0_0WCLKN_net ),
            .I(N__16991));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_7 ),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_16_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_15_0_));
    defparam IN_MUX_bfv_16_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_18_0_));
    defparam IN_MUX_bfv_16_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_19_0_ (
            .carryinitin(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_7_s1 ),
            .carryinitout(bfn_16_19_0_));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_13_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_13_0_ (
            .carryinitin(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_7 ),
            .carryinitout(bfn_13_13_0_));
    defparam IN_MUX_bfv_14_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_11_0_));
    defparam IN_MUX_bfv_14_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_12_0_ (
            .carryinitin(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_7 ),
            .carryinitout(bfn_14_12_0_));
    defparam IN_MUX_bfv_17_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_6_0_));
    defparam IN_MUX_bfv_17_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_7_0_ (
            .carryinitin(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_7 ),
            .carryinitout(bfn_17_7_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_7 ),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_13_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_2_0_));
    defparam IN_MUX_bfv_13_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_3_0_ (
            .carryinitin(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_7 ),
            .carryinitout(bfn_13_3_0_));
    defparam IN_MUX_bfv_15_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_3_0_));
    defparam IN_MUX_bfv_15_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_4_0_ (
            .carryinitin(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_7 ),
            .carryinitout(bfn_15_4_0_));
    defparam IN_MUX_bfv_17_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_2_0_));
    defparam IN_MUX_bfv_17_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_3_0_ (
            .carryinitin(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_7 ),
            .carryinitout(bfn_17_3_0_));
    defparam IN_MUX_bfv_15_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_5_0_));
    defparam IN_MUX_bfv_15_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_6_0_ (
            .carryinitin(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_7 ),
            .carryinitout(bfn_15_6_0_));
    ICE_GB N_292_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__6764),
            .GLOBALBUFFEROUTPUT(N_292_g));
    ICE_GB wPllLocked_i_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__14101),
            .GLOBALBUFFEROUTPUT(wPllLocked_i_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0 .C_ON=1'b0;
    defparam \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0 .SEQ_MODE=4'b0000;
    defparam \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PLL_BUFFER_top_pll_inst.top_pll_inst_LOCK_THRU_LUT4_0_LC_1_30_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6467),
            .lcout(wPllLocked),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.wPllLocked_i_LC_8_16_5 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.wPllLocked_i_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.wPllLocked_i_LC_8_16_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uart_inst0.uart_inst0.wPllLocked_i_LC_8_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13921),
            .lcout(wPllLocked_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_0_c_LC_9_14_0 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_0_c_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_0_c_LC_9_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \uart_inst0.uart_inst0.un2_rx_clk_divider_cry_0_c_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__6679),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_clk_divider_1_LC_9_14_1 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_1_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_1_LC_9_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_inst0.uart_inst0.rx_clk_divider_1_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(N__6725),
            .in2(N__12338),
            .in3(N__6491),
            .lcout(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_1 ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_0 ),
            .carryout(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_1 ),
            .clk(N__16923),
            .ce(),
            .sr(N__6661));
    defparam \uart_inst0.uart_inst0.rx_clk_divider_2_LC_9_14_2 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_2_LC_9_14_2 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_2_LC_9_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_inst0.uart_inst0.rx_clk_divider_2_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__6698),
            .in2(N__12342),
            .in3(N__6488),
            .lcout(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_2 ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_1 ),
            .carryout(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_2 ),
            .clk(N__16923),
            .ce(),
            .sr(N__6661));
    defparam \uart_inst0.uart_inst0.rx_clk_divider_3_LC_9_14_3 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_3_LC_9_14_3 .SEQ_MODE=4'b1001;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_3_LC_9_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_inst0.uart_inst0.rx_clk_divider_3_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__6737),
            .in2(N__12339),
            .in3(N__6485),
            .lcout(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_3 ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_2 ),
            .carryout(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_3 ),
            .clk(N__16923),
            .ce(),
            .sr(N__6661));
    defparam \uart_inst0.uart_inst0.rx_clk_divider_4_LC_9_14_4 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_4_LC_9_14_4 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_4_LC_9_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_inst0.uart_inst0.rx_clk_divider_4_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(N__6712),
            .in2(N__12343),
            .in3(N__6482),
            .lcout(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_4 ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_3 ),
            .carryout(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_4 ),
            .clk(N__16923),
            .ce(),
            .sr(N__6661));
    defparam \uart_inst0.uart_inst0.rx_clk_divider_5_LC_9_14_5 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_5_LC_9_14_5 .SEQ_MODE=4'b1001;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_5_LC_9_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_inst0.uart_inst0.rx_clk_divider_5_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(N__6503),
            .in2(N__12340),
            .in3(N__6479),
            .lcout(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_5 ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_4 ),
            .carryout(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_5 ),
            .clk(N__16923),
            .ce(),
            .sr(N__6661));
    defparam \uart_inst0.uart_inst0.rx_clk_divider_6_LC_9_14_6 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_6_LC_9_14_6 .SEQ_MODE=4'b1001;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_6_LC_9_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_inst0.uart_inst0.rx_clk_divider_6_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(N__6515),
            .in2(N__12344),
            .in3(N__6476),
            .lcout(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_6 ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_5 ),
            .carryout(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_6 ),
            .clk(N__16923),
            .ce(),
            .sr(N__6661));
    defparam \uart_inst0.uart_inst0.rx_clk_divider_7_LC_9_14_7 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_7_LC_9_14_7 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_7_LC_9_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_inst0.uart_inst0.rx_clk_divider_7_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(N__6614),
            .in2(N__12341),
            .in3(N__6473),
            .lcout(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_7 ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_6 ),
            .carryout(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_7 ),
            .clk(N__16923),
            .ce(),
            .sr(N__6661));
    defparam \uart_inst0.uart_inst0.rx_clk_divider_8_LC_9_15_0 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_8_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_8_LC_9_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_inst0.uart_inst0.rx_clk_divider_8_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__6626),
            .in2(N__12404),
            .in3(N__6470),
            .lcout(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_8 ),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_8 ),
            .clk(N__16917),
            .ce(),
            .sr(N__6662));
    defparam \uart_inst0.uart_inst0.rx_clk_divider_9_LC_9_15_1 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_9_LC_9_15_1 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_9_LC_9_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_inst0.uart_inst0.rx_clk_divider_9_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__12356),
            .in2(N__6545),
            .in3(N__6644),
            .lcout(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_9 ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_8 ),
            .carryout(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_9 ),
            .clk(N__16917),
            .ce(),
            .sr(N__6662));
    defparam \uart_inst0.uart_inst0.rx_clk_divider_10_LC_9_15_2 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_10_LC_9_15_2 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_10_LC_9_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_inst0.uart_inst0.rx_clk_divider_10_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__6587),
            .in2(N__12402),
            .in3(N__6641),
            .lcout(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_10 ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_9 ),
            .carryout(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_10 ),
            .clk(N__16917),
            .ce(),
            .sr(N__6662));
    defparam \uart_inst0.uart_inst0.rx_clk_divider_11_LC_9_15_3 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_11_LC_9_15_3 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_11_LC_9_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_inst0.uart_inst0.rx_clk_divider_11_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__12348),
            .in2(N__6575),
            .in3(N__6638),
            .lcout(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_11 ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_10 ),
            .carryout(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_11 ),
            .clk(N__16917),
            .ce(),
            .sr(N__6662));
    defparam \uart_inst0.uart_inst0.rx_clk_divider_12_LC_9_15_4 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_12_LC_9_15_4 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_12_LC_9_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_inst0.uart_inst0.rx_clk_divider_12_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__6559),
            .in2(N__12403),
            .in3(N__6635),
            .lcout(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_12 ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_11 ),
            .carryout(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_12 ),
            .clk(N__16917),
            .ce(),
            .sr(N__6662));
    defparam \uart_inst0.uart_inst0.rx_clk_divider_13_LC_9_15_5 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_13_LC_9_15_5 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_13_LC_9_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_inst0.uart_inst0.rx_clk_divider_13_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(N__12352),
            .in2(N__6530),
            .in3(N__6632),
            .lcout(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_13 ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_12 ),
            .carryout(\uart_inst0.uart_inst0.un2_rx_clk_divider_cry_13 ),
            .clk(N__16917),
            .ce(),
            .sr(N__6662));
    defparam \uart_inst0.uart_inst0.rx_clk_divider_14_LC_9_15_6 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_14_LC_9_15_6 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_14_LC_9_15_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \uart_inst0.uart_inst0.rx_clk_divider_14_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(N__6601),
            .in2(_gnd_net_),
            .in3(N__6629),
            .lcout(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16917),
            .ce(),
            .sr(N__6662));
    defparam \uart_inst0.uart_inst0.rx_clk_divider_RNI0H8H_14_LC_10_14_0 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_RNI0H8H_14_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_RNI0H8H_14_LC_10_14_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_inst0.uart_inst0.rx_clk_divider_RNI0H8H_14_LC_10_14_0  (
            .in0(N__6625),
            .in1(N__6613),
            .in2(N__6602),
            .in3(N__6678),
            .lcout(\uart_inst0.uart_inst0.un1_rx_clk_divider_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_clk_divider_RNIRKBC1_9_LC_10_14_2 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_RNIRKBC1_9_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_RNIRKBC1_9_LC_10_14_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_inst0.uart_inst0.rx_clk_divider_RNIRKBC1_9_LC_10_14_2  (
            .in0(N__6586),
            .in1(N__6571),
            .in2(N__6560),
            .in3(N__6541),
            .lcout(\uart_inst0.uart_inst0.un1_rx_clk_divider_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_clk_divider_RNISPAG_5_LC_10_14_3 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_RNISPAG_5_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_RNISPAG_5_LC_10_14_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart_inst0.uart_inst0.rx_clk_divider_RNISPAG_5_LC_10_14_3  (
            .in0(N__6526),
            .in1(N__6514),
            .in2(_gnd_net_),
            .in3(N__6502),
            .lcout(),
            .ltout(\uart_inst0.uart_inst0.un1_rx_clk_divider_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_clk_divider_RNITHLH2_1_LC_10_14_4 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_RNITHLH2_1_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_RNITHLH2_1_LC_10_14_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uart_inst0.uart_inst0.rx_clk_divider_RNITHLH2_1_LC_10_14_4  (
            .in0(N__6755),
            .in1(N__6749),
            .in2(N__6743),
            .in3(N__6686),
            .lcout(\uart_inst0.uart_inst0.un1_rx_clk_divider_0 ),
            .ltout(\uart_inst0.uart_inst0.un1_rx_clk_divider_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_state_RNIPLGK2_0_LC_10_14_5 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_state_RNIPLGK2_0_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_state_RNIPLGK2_0_LC_10_14_5 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \uart_inst0.uart_inst0.rx_state_RNIPLGK2_0_LC_10_14_5  (
            .in0(N__13894),
            .in1(_gnd_net_),
            .in2(N__6740),
            .in3(N__11155),
            .lcout(\uart_inst0.uart_inst0.rx_clk_divider_1_sqmuxa_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_clk_divider_RNI6IM3_1_LC_10_14_6 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_RNI6IM3_1_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_RNI6IM3_1_LC_10_14_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_inst0.uart_inst0.rx_clk_divider_RNI6IM3_1_LC_10_14_6  (
            .in0(N__6736),
            .in1(N__6724),
            .in2(N__6713),
            .in3(N__6697),
            .lcout(\uart_inst0.uart_inst0.un1_rx_clk_divider_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_clk_divider_0_LC_10_15_6 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_0_LC_10_15_6 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_clk_divider_0_LC_10_15_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uart_inst0.uart_inst0.rx_clk_divider_0_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6680),
            .lcout(\uart_inst0.uart_inst0.rx_clk_dividerZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16909),
            .ce(),
            .sr(N__6660));
    defparam \fifo_inst.tx_fifo_inst.rDataCount_3_LC_12_2_4 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_3_LC_12_2_4 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_3_LC_12_2_4 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rDataCount_3_LC_12_2_4  (
            .in0(N__7966),
            .in1(N__7866),
            .in2(N__7951),
            .in3(N__10161),
            .lcout(wTxFull),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16958),
            .ce(),
            .sr(N__16340));
    defparam rTxEn_LC_12_2_6.C_ON=1'b0;
    defparam rTxEn_LC_12_2_6.SEQ_MODE=4'b1000;
    defparam rTxEn_LC_12_2_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 rTxEn_LC_12_2_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10160),
            .lcout(rTxEnZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16958),
            .ce(),
            .sr(N__16340));
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNIA7U81_2_LC_12_3_1 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNIA7U81_2_LC_12_3_1 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNIA7U81_2_LC_12_3_1 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \fifo_inst.tx_fifo_inst.rDataCount_RNIA7U81_2_LC_12_3_1  (
            .in0(N__7825),
            .in1(N__7787),
            .in2(N__9259),
            .in3(N__7721),
            .lcout(\fifo_inst.tx_fifo_inst.un1_rDataCount_axbxc3_2_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNIEM211_2_LC_12_3_2 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNIEM211_2_LC_12_3_2 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNIEM211_2_LC_12_3_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rDataCount_RNIEM211_2_LC_12_3_2  (
            .in0(N__9303),
            .in1(N__9251),
            .in2(_gnd_net_),
            .in3(N__7826),
            .lcout(\fifo_inst.tx_fifo_inst.un1_rDataCount_axbxc3_a0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNIDPRL_0_LC_12_3_7 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNIDPRL_0_LC_12_3_7 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNIDPRL_0_LC_12_3_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rDataCount_RNIDPRL_0_LC_12_3_7  (
            .in0(_gnd_net_),
            .in1(N__7786),
            .in2(_gnd_net_),
            .in3(N__7720),
            .lcout(\fifo_inst.tx_fifo_inst.un1_rDataCount_ac0_1_a0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ft2232h_inst.rRx_n_LC_12_4_1 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rRx_n_LC_12_4_1 .SEQ_MODE=4'b1001;
    defparam \fifo_inst.ft2232h_inst.rRx_n_LC_12_4_1 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \fifo_inst.ft2232h_inst.rRx_n_LC_12_4_1  (
            .in0(N__6801),
            .in1(N__6785),
            .in2(_gnd_net_),
            .in3(N__8150),
            .lcout(P1A3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16946),
            .ce(),
            .sr(N__16350));
    defparam \uart_inst0.tx_uart_fifo_inst.m39_LC_12_5_0 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m39_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m39_LC_12_5_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m39_LC_12_5_0  (
            .in0(N__8116),
            .in1(N__8078),
            .in2(_gnd_net_),
            .in3(N__12764),
            .lcout(N_86_mux),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_3_LC_12_11_6 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_3_LC_12_11_6 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_3_LC_12_11_6 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_3_LC_12_11_6  (
            .in0(N__6776),
            .in1(N__7322),
            .in2(N__8645),
            .in3(N__8505),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16918),
            .ce(),
            .sr(N__13595));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNIVHG3_8_LC_12_12_0 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNIVHG3_8_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNIVHG3_8_LC_12_12_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNIVHG3_8_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__7563),
            .in2(_gnd_net_),
            .in3(N__7338),
            .lcout(),
            .ltout(\uart_inst0.tx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNI0VO8_0_LC_12_12_1 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNI0VO8_0_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNI0VO8_0_LC_12_12_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNI0VO8_0_LC_12_12_1  (
            .in0(N__7375),
            .in1(N__7405),
            .in2(N__6779),
            .in3(N__7435),
            .lcout(\uart_inst0.tx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ0Z_0_LC_12_13_2 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ0Z_0_LC_12_13_2 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ0Z_0_LC_12_13_2 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ0Z_0_LC_12_13_2  (
            .in0(N__6775),
            .in1(N__7415),
            .in2(N__8644),
            .in3(N__8515),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16908),
            .ce(),
            .sr(N__13593));
    defparam GB_BUFFER_wPllLocked_i_g_THRU_LUT4_0_LC_12_30_0.C_ON=1'b0;
    defparam GB_BUFFER_wPllLocked_i_g_THRU_LUT4_0_LC_12_30_0.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_wPllLocked_i_g_THRU_LUT4_0_LC_12_30_0.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_wPllLocked_i_g_THRU_LUT4_0_LC_12_30_0 (
            .in0(N__16696),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_wPllLocked_i_g_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNIQ7UO_3_LC_13_1_1 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNIQ7UO_3_LC_13_1_1 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNIQ7UO_3_LC_13_1_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rDataCount_RNIQ7UO_3_LC_13_1_1  (
            .in0(_gnd_net_),
            .in1(N__10143),
            .in2(_gnd_net_),
            .in3(N__9288),
            .lcout(fifo_inst_tx_fifo_inst_wRamWrEn),
            .ltout(fifo_inst_tx_fifo_inst_wRamWrEn_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_3_LC_13_1_2 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_3_LC_13_1_2 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_3_LC_13_1_2 .LUT_INIT=16'b0001101100000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamWrAddr_3_LC_13_1_2  (
            .in0(N__6995),
            .in1(N__16619),
            .in2(N__6758),
            .in3(N__6863),
            .lcout(fifo_inst_tx_fifo_inst_rRamWrAddr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16971),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_0_LC_13_1_4 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_0_LC_13_1_4 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_0_LC_13_1_4 .LUT_INIT=16'b0000100000101010;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamWrAddr_0_LC_13_1_4  (
            .in0(N__6953),
            .in1(N__6994),
            .in2(N__7923),
            .in3(N__16618),
            .lcout(fifo_inst_tx_fifo_inst_rRamWrAddr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16971),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m68_e_6_LC_13_1_5 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m68_e_6_LC_13_1_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m68_e_6_LC_13_1_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m68_e_6_LC_13_1_5  (
            .in0(N__6879),
            .in1(N__6939),
            .in2(N__7045),
            .in3(N__6969),
            .lcout(\uart_inst0.tx_uart_fifo_inst.m68_eZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m68_e_5_LC_13_1_6 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m68_e_5_LC_13_1_6 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m68_e_5_LC_13_1_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m68_e_5_LC_13_1_6  (
            .in0(N__7135),
            .in1(N__16620),
            .in2(N__6854),
            .in3(N__6909),
            .lcout(),
            .ltout(\uart_inst0.tx_uart_fifo_inst.m68_eZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m68_e_LC_13_1_7 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m68_e_LC_13_1_7 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m68_e_LC_13_1_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m68_e_LC_13_1_7  (
            .in0(N__7074),
            .in1(N__7101),
            .in2(N__7004),
            .in3(N__7001),
            .lcout(\uart_inst0.tx_uart_fifo_inst.N_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_RNI10581_0_LC_13_2_0 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_RNI10581_0_LC_13_2_0 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_RNI10581_0_LC_13_2_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamWrAddr_RNI10581_0_LC_13_2_0  (
            .in0(_gnd_net_),
            .in1(N__6970),
            .in2(N__7919),
            .in3(N__7918),
            .lcout(rRamWrAddr_RNI10581_0),
            .ltout(),
            .carryin(bfn_13_2_0_),
            .carryout(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_1_LC_13_2_1 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_1_LC_13_2_1 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_1_LC_13_2_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamWrAddr_1_LC_13_2_1  (
            .in0(N__16621),
            .in1(N__6940),
            .in2(_gnd_net_),
            .in3(N__6923),
            .lcout(fifo_inst_tx_fifo_inst_rRamWrAddr_1),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_0 ),
            .carryout(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_1 ),
            .clk(N__16966),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_2_LC_13_2_2 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_2_LC_13_2_2 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_2_LC_13_2_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamWrAddr_2_LC_13_2_2  (
            .in0(N__16624),
            .in1(N__6910),
            .in2(_gnd_net_),
            .in3(N__6893),
            .lcout(fifo_inst_tx_fifo_inst_rRamWrAddr_2),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_1 ),
            .carryout(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_2 ),
            .clk(N__16966),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_2_c_RNISJKU_LC_13_2_3 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_2_c_RNISJKU_LC_13_2_3 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_2_c_RNISJKU_LC_13_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_2_c_RNISJKU_LC_13_2_3  (
            .in0(_gnd_net_),
            .in1(N__6880),
            .in2(_gnd_net_),
            .in3(N__6857),
            .lcout(un1_rRamWrAddr_cry_2_c_RNISJKU),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_2 ),
            .carryout(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_4_LC_13_2_4 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_4_LC_13_2_4 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_4_LC_13_2_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamWrAddr_4_LC_13_2_4  (
            .in0(N__16625),
            .in1(N__6843),
            .in2(_gnd_net_),
            .in3(N__6824),
            .lcout(fifo_inst_tx_fifo_inst_rRamWrAddr_4),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_3 ),
            .carryout(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_4 ),
            .clk(N__16966),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_5_LC_13_2_5 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_5_LC_13_2_5 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_5_LC_13_2_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamWrAddr_5_LC_13_2_5  (
            .in0(N__16622),
            .in1(N__7131),
            .in2(_gnd_net_),
            .in3(N__7112),
            .lcout(fifo_inst_tx_fifo_inst_rRamWrAddr_5),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_4 ),
            .carryout(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_5 ),
            .clk(N__16966),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_6_LC_13_2_6 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_6_LC_13_2_6 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_6_LC_13_2_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamWrAddr_6_LC_13_2_6  (
            .in0(N__16626),
            .in1(N__7102),
            .in2(_gnd_net_),
            .in3(N__7085),
            .lcout(fifo_inst_tx_fifo_inst_rRamWrAddr_6),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_5 ),
            .carryout(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_6 ),
            .clk(N__16966),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_7_LC_13_2_7 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_7_LC_13_2_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_7_LC_13_2_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamWrAddr_7_LC_13_2_7  (
            .in0(N__16623),
            .in1(N__7078),
            .in2(_gnd_net_),
            .in3(N__7058),
            .lcout(fifo_inst_tx_fifo_inst_rRamWrAddr_7),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_6 ),
            .carryout(\fifo_inst.tx_fifo_inst.un1_rRamWrAddr_cry_7 ),
            .clk(N__16966),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_8_LC_13_3_0 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_8_LC_13_3_0 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rRamWrAddr_8_LC_13_3_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamWrAddr_8_LC_13_3_0  (
            .in0(N__16627),
            .in1(N__7038),
            .in2(_gnd_net_),
            .in3(N__7055),
            .lcout(fifo_inst_tx_fifo_inst_rRamWrAddr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16959),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNO_3_2_LC_13_3_1 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNO_3_2_LC_13_3_1 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNO_3_2_LC_13_3_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \fifo_inst.tx_fifo_inst.rDataCount_RNO_3_2_LC_13_3_1  (
            .in0(_gnd_net_),
            .in1(N__9239),
            .in2(_gnd_net_),
            .in3(N__7772),
            .lcout(\fifo_inst.tx_fifo_inst.un1_rDataCount_ac0_1_a1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rFifoState_12_0_i_LC_13_3_2 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rFifoState_12_0_i_LC_13_3_2 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rFifoState_12_0_i_LC_13_3_2 .LUT_INIT=16'b1100110011001110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.un1_rFifoState_12_0_i_LC_13_3_2  (
            .in0(N__10636),
            .in1(N__8258),
            .in2(N__10613),
            .in3(N__10499),
            .lcout(),
            .ltout(fifo_inst_ft2232h_inst_un1_rFifoState_12_0_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ft2232h_inst.rTxRdEn_esr_RNO_LC_13_3_3 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rTxRdEn_esr_RNO_LC_13_3_3 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ft2232h_inst.rTxRdEn_esr_RNO_LC_13_3_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \fifo_inst.ft2232h_inst.rTxRdEn_esr_RNO_LC_13_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__7016),
            .in3(N__14102),
            .lcout(\fifo_inst.ft2232h_inst.un1_rFifoState_12_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m78_bm_LC_13_3_5 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m78_bm_LC_13_3_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m78_bm_LC_13_3_5 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m78_bm_LC_13_3_5  (
            .in0(N__7815),
            .in1(N__7773),
            .in2(N__10162),
            .in3(N__7717),
            .lcout(\uart_inst0.tx_uart_fifo_inst.m78_bmZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNO_2_2_LC_13_3_7 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNO_2_2_LC_13_3_7 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNO_2_2_LC_13_3_7 .LUT_INIT=16'b1011000000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rDataCount_RNO_2_2_LC_13_3_7  (
            .in0(N__10147),
            .in1(N__9295),
            .in2(N__7013),
            .in3(N__7718),
            .lcout(\fifo_inst.tx_fifo_inst.un1_rDataCount_c2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m78_ns_1_LC_13_4_0 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m78_ns_1_LC_13_4_0 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m78_ns_1_LC_13_4_0 .LUT_INIT=16'b0011001101000100;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m78_ns_1_LC_13_4_0  (
            .in0(N__10163),
            .in1(N__9302),
            .in2(_gnd_net_),
            .in3(N__9257),
            .lcout(),
            .ltout(\uart_inst0.tx_uart_fifo_inst.m78_nsZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m78_ns_LC_13_4_1 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m78_ns_LC_13_4_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m78_ns_LC_13_4_1 .LUT_INIT=16'b1010110100001101;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m78_ns_LC_13_4_1  (
            .in0(N__9258),
            .in1(N__7166),
            .in2(N__7160),
            .in3(N__10523),
            .lcout(fifo_inst_tx_fifo_inst_un1_rDataCount15_2_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ft2232h_inst.rTxRdEn_esr_LC_13_4_3 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rTxRdEn_esr_LC_13_4_3 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rTxRdEn_esr_LC_13_4_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \fifo_inst.ft2232h_inst.rTxRdEn_esr_LC_13_4_3  (
            .in0(N__10608),
            .in1(N__10656),
            .in2(_gnd_net_),
            .in3(N__10524),
            .lcout(fifo_inst_wTxRdEn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16952),
            .ce(N__7157),
            .sr(N__16355));
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNI1JE32_0_LC_13_4_5 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNI1JE32_0_LC_13_4_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNI1JE32_0_LC_13_4_5 .LUT_INIT=16'b0101010010100000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rDataCount_RNI1JE32_0_LC_13_4_5  (
            .in0(N__8491),
            .in1(N__8419),
            .in2(N__8360),
            .in3(N__9509),
            .lcout(\uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c2_d ),
            .ltout(\uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c2_d_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNO_0_3_LC_13_4_6 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNO_0_3_LC_13_4_6 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNO_0_3_LC_13_4_6 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rDataCount_RNO_0_3_LC_13_4_6  (
            .in0(N__8420),
            .in1(N__7263),
            .in2(N__7148),
            .in3(N__8387),
            .lcout(\uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIO6DU2_3_LC_13_4_7 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIO6DU2_3_LC_13_4_7 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIO6DU2_3_LC_13_4_7 .LUT_INIT=16'b0000110100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIO6DU2_3_LC_13_4_7  (
            .in0(N__7313),
            .in1(N__8316),
            .in2(N__9850),
            .in3(N__9508),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rDataCount_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m14_LC_13_5_0 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m14_LC_13_5_0 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m14_LC_13_5_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m14_LC_13_5_0  (
            .in0(N__8221),
            .in1(N__12689),
            .in2(N__8039),
            .in3(N__12587),
            .lcout(N_84_mux),
            .ltout(N_84_mux_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m17_LC_13_5_1 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m17_LC_13_5_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m17_LC_13_5_1 .LUT_INIT=16'b1000101000000010;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m17_LC_13_5_1  (
            .in0(N__15364),
            .in1(N__9074),
            .in2(N__7145),
            .in3(N__12757),
            .lcout(fifo_inst_rx_fifo_inst_rDataCount_0_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m65_bm_LC_13_5_2 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m65_bm_LC_13_5_2 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m65_bm_LC_13_5_2 .LUT_INIT=16'b0101010101010100;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m65_bm_LC_13_5_2  (
            .in0(N__12755),
            .in1(N__12690),
            .in2(N__12650),
            .in3(N__12588),
            .lcout(),
            .ltout(\uart_inst0.tx_uart_fifo_inst.m65_bmZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m65_ns_LC_13_5_3 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m65_ns_LC_13_5_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m65_ns_LC_13_5_3 .LUT_INIT=16'b1011100100110001;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m65_ns_LC_13_5_3  (
            .in0(N__15365),
            .in1(N__7199),
            .in2(N__7205),
            .in3(N__8199),
            .lcout(fifo_inst_rx_fifo_inst_un1_rDataCount15_2_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rDataCount_RNO_2_2_LC_13_5_4 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.rDataCount_RNO_2_2_LC_13_5_4 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.rx_fifo_inst.rDataCount_RNO_2_2_LC_13_5_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \fifo_inst.rx_fifo_inst.rDataCount_RNO_2_2_LC_13_5_4  (
            .in0(N__12756),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9073),
            .lcout(),
            .ltout(\fifo_inst.rx_fifo_inst.un1_rDataCount_c2_1_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rDataCount_RNO_1_2_LC_13_5_5 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.rDataCount_RNO_1_2_LC_13_5_5 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.rx_fifo_inst.rDataCount_RNO_1_2_LC_13_5_5 .LUT_INIT=16'b0100001000000000;
    LogicCell40 \fifo_inst.rx_fifo_inst.rDataCount_RNO_1_2_LC_13_5_5  (
            .in0(N__15367),
            .in1(N__12592),
            .in2(N__7202),
            .in3(N__12637),
            .lcout(\fifo_inst.rx_fifo_inst.un1_rDataCount_c2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m65_ns_1_LC_13_5_6 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m65_ns_1_LC_13_5_6 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m65_ns_1_LC_13_5_6 .LUT_INIT=16'b0011001101000100;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m65_ns_1_LC_13_5_6  (
            .in0(N__12754),
            .in1(N__9072),
            .in2(_gnd_net_),
            .in3(N__15363),
            .lcout(\uart_inst0.tx_uart_fifo_inst.m65_nsZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rDataCount_RNO_0_2_LC_13_5_7 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.rDataCount_RNO_0_2_LC_13_5_7 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.rx_fifo_inst.rDataCount_RNO_0_2_LC_13_5_7 .LUT_INIT=16'b1000000010100000;
    LogicCell40 \fifo_inst.rx_fifo_inst.rDataCount_RNO_0_2_LC_13_5_7  (
            .in0(N__15366),
            .in1(N__12758),
            .in2(N__12598),
            .in3(N__9075),
            .lcout(\fifo_inst.rx_fifo_inst.un1_rDataCount_ac0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rDataCount_1_LC_13_6_3 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.rDataCount_1_LC_13_6_3 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rDataCount_1_LC_13_6_3 .LUT_INIT=16'b0100101110110100;
    LogicCell40 \fifo_inst.rx_fifo_inst.rDataCount_1_LC_13_6_3  (
            .in0(N__8237),
            .in1(N__12646),
            .in2(N__7187),
            .in3(N__12594),
            .lcout(fifo_inst_rx_fifo_inst_rDataCount_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16941),
            .ce(),
            .sr(N__16366));
    defparam \fifo_inst.rx_fifo_inst.rDataCount_2_LC_13_6_6 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.rDataCount_2_LC_13_6_6 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rDataCount_2_LC_13_6_6 .LUT_INIT=16'b1100100100110110;
    LogicCell40 \fifo_inst.rx_fifo_inst.rDataCount_2_LC_13_6_6  (
            .in0(N__7193),
            .in1(N__7183),
            .in2(N__7175),
            .in3(N__12691),
            .lcout(fifo_inst_rx_fifo_inst_rDataCount_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16941),
            .ce(),
            .sr(N__16366));
    defparam rUartTxEn_LC_13_7_4.C_ON=1'b0;
    defparam rUartTxEn_LC_13_7_4.SEQ_MODE=4'b1000;
    defparam rUartTxEn_LC_13_7_4.LUT_INIT=16'b0000000011101110;
    LogicCell40 rUartTxEn_LC_13_7_4 (
            .in0(N__11217),
            .in1(N__15376),
            .in2(_gnd_net_),
            .in3(N__8318),
            .lcout(rUartTxEnZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16938),
            .ce(),
            .sr(N__16384));
    defparam rUartRxFlag_LC_13_7_6.C_ON=1'b0;
    defparam rUartRxFlag_LC_13_7_6.SEQ_MODE=4'b1000;
    defparam rUartRxFlag_LC_13_7_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 rUartRxFlag_LC_13_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13049),
            .lcout(rUartRxFlagZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16938),
            .ce(),
            .sr(N__16384));
    defparam CONSTANT_ONE_LUT4_LC_13_8_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_13_8_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_13_8_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_13_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIPA3Q_3_LC_13_8_1 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIPA3Q_3_LC_13_8_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIPA3Q_3_LC_13_8_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIPA3Q_3_LC_13_8_1  (
            .in0(_gnd_net_),
            .in1(N__7309),
            .in2(_gnd_net_),
            .in3(N__8301),
            .lcout(\uart_inst0.tx_uart_fifo_inst.wRamWrEn_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCountZ0Z_0_LC_13_9_0 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCountZ0Z_0_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCountZ0Z_0_LC_13_9_0 .LUT_INIT=16'b0101100110100110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rDataCountZ0Z_0_LC_13_9_0  (
            .in0(N__8475),
            .in1(N__9499),
            .in2(N__9848),
            .in3(N__8356),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16930),
            .ce(),
            .sr(N__16413));
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_3_LC_13_9_6 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_3_LC_13_9_6 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_3_LC_13_9_6 .LUT_INIT=16'b1011100101000110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rDataCount_3_LC_13_9_6  (
            .in0(N__7270),
            .in1(N__7298),
            .in2(N__7286),
            .in3(N__8314),
            .lcout(\uart_inst0.tx_uart_fifo_inst.wUartTxFull ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16930),
            .ce(),
            .sr(N__16413));
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_2_LC_13_10_0 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_2_LC_13_10_0 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_2_LC_13_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rDataCount_2_LC_13_10_0  (
            .in0(N__8522),
            .in1(N__7271),
            .in2(_gnd_net_),
            .in3(N__8382),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rDataCountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16926),
            .ce(),
            .sr(N__16415));
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIA3TL1_2_LC_13_10_5 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIA3TL1_2_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIA3TL1_2_LC_13_10_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIA3TL1_2_LC_13_10_5  (
            .in0(N__8381),
            .in1(N__8351),
            .in2(N__8315),
            .in3(N__8410),
            .lcout(\uart_inst0.wTxRdEmpty ),
            .ltout(\uart_inst0.wTxRdEmpty_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rTxRdEn_LC_13_10_6 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rTxRdEn_LC_13_10_6 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rTxRdEn_LC_13_10_6 .LUT_INIT=16'b1011101100000001;
    LogicCell40 \uart_inst0.uart_inst0.rTxRdEn_LC_13_10_6  (
            .in0(N__11591),
            .in1(N__11669),
            .in2(N__7250),
            .in3(N__9500),
            .lcout(\uart_inst0.wTxRdEn_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16926),
            .ce(),
            .sr(N__16415));
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0_LC_13_11_0 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0_LC_13_11_0 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0_LC_13_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7247),
            .lcout(\uart_inst0.wTxRdData_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net ),
            .ce(N__9593),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_1_LC_13_11_1 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_1_LC_13_11_1 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_1_LC_13_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_1_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7232),
            .lcout(\uart_inst0.wTxRdData_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net ),
            .ce(N__9593),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_2_LC_13_11_2 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_2_LC_13_11_2 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_2_LC_13_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_2_LC_13_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7217),
            .lcout(\uart_inst0.wTxRdData_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net ),
            .ce(N__9593),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_3_LC_13_11_3 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_3_LC_13_11_3 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_3_LC_13_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_3_LC_13_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7505),
            .lcout(\uart_inst0.wTxRdData_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net ),
            .ce(N__9593),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_4_LC_13_11_4 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_4_LC_13_11_4 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_4_LC_13_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_4_LC_13_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7490),
            .lcout(\uart_inst0.wTxRdData_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net ),
            .ce(N__9593),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_5_LC_13_11_5 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_5_LC_13_11_5 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_5_LC_13_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_5_LC_13_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7478),
            .lcout(\uart_inst0.wTxRdData_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net ),
            .ce(N__9593),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_6_LC_13_11_6 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_6_LC_13_11_6 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_6_LC_13_11_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_6_LC_13_11_6  (
            .in0(N__7466),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart_inst0.wTxRdData_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net ),
            .ce(N__9593),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_7_LC_13_11_7 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_7_LC_13_11_7 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_7_LC_13_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_7_LC_13_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7457),
            .lcout(\uart_inst0.wTxRdData_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuart_inst0.tx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net ),
            .ce(N__9593),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNO_0_0_LC_13_12_0 .C_ON=1'b1;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNO_0_0_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNO_0_0_LC_13_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNO_0_0_LC_13_12_0  (
            .in0(_gnd_net_),
            .in1(N__7431),
            .in2(N__8516),
            .in3(N__8514),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ0Z_1_LC_13_12_1 .C_ON=1'b1;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ0Z_1_LC_13_12_1 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ0Z_1_LC_13_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ0Z_1_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__7401),
            .in2(_gnd_net_),
            .in3(N__7385),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ1Z_1 ),
            .ltout(),
            .carryin(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_0 ),
            .carryout(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_1 ),
            .clk(N__16919),
            .ce(),
            .sr(N__13596));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_2_LC_13_12_2 .C_ON=1'b1;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_2_LC_13_12_2 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_2_LC_13_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_2_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(N__7371),
            .in2(_gnd_net_),
            .in3(N__7355),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rRamWrAddrZ0Z_2 ),
            .ltout(),
            .carryin(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_1 ),
            .carryout(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_2 ),
            .clk(N__16919),
            .ce(),
            .sr(N__13596));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNO_0_3_LC_13_12_3 .C_ON=1'b1;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNO_0_3_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNO_0_3_LC_13_12_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNO_0_3_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(N__7339),
            .in2(_gnd_net_),
            .in3(N__7316),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_2 ),
            .carryout(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_4_LC_13_12_4 .C_ON=1'b1;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_4_LC_13_12_4 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_4_LC_13_12_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_4_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(N__8661),
            .in2(_gnd_net_),
            .in3(N__7592),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_4 ),
            .ltout(),
            .carryin(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_3 ),
            .carryout(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_4 ),
            .clk(N__16919),
            .ce(),
            .sr(N__13596));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_5_LC_13_12_5 .C_ON=1'b1;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_5_LC_13_12_5 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_5_LC_13_12_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_5_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(N__8712),
            .in2(_gnd_net_),
            .in3(N__7589),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_5 ),
            .ltout(),
            .carryin(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_4 ),
            .carryout(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_5 ),
            .clk(N__16919),
            .ce(),
            .sr(N__13596));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_6_LC_13_12_6 .C_ON=1'b1;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_6_LC_13_12_6 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_6_LC_13_12_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_6_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(N__8685),
            .in2(_gnd_net_),
            .in3(N__7586),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_6 ),
            .ltout(),
            .carryin(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_5 ),
            .carryout(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_6 ),
            .clk(N__16919),
            .ce(),
            .sr(N__13596));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_7_LC_13_12_7 .C_ON=1'b1;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_7_LC_13_12_7 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_7_LC_13_12_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_7_LC_13_12_7  (
            .in0(_gnd_net_),
            .in1(N__8742),
            .in2(_gnd_net_),
            .in3(N__7583),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_7 ),
            .ltout(),
            .carryin(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_6 ),
            .carryout(\uart_inst0.tx_uart_fifo_inst.un1_rRamWrAddr_cry_7 ),
            .clk(N__16919),
            .ce(),
            .sr(N__13596));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_8_LC_13_13_0 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_8_LC_13_13_0 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_8_LC_13_13_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_8_LC_13_13_0  (
            .in0(_gnd_net_),
            .in1(N__7567),
            .in2(_gnd_net_),
            .in3(N__7580),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rRamWrAddr_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16913),
            .ce(),
            .sr(N__13594));
    defparam \uart_inst0.uart_inst0.rTxData_esr_0_LC_13_14_0 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rTxData_esr_0_LC_13_14_0 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rTxData_esr_0_LC_13_14_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uart_inst0.uart_inst0.rTxData_esr_0_LC_13_14_0  (
            .in0(N__7529),
            .in1(N__8574),
            .in2(_gnd_net_),
            .in3(N__7547),
            .lcout(\uart_inst0.uart_inst0.rTxDataZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16910),
            .ce(N__8813),
            .sr(N__16436));
    defparam \uart_inst0.uart_inst0.rTxData_esr_1_LC_13_14_6 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rTxData_esr_1_LC_13_14_6 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rTxData_esr_1_LC_13_14_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uart_inst0.uart_inst0.rTxData_esr_1_LC_13_14_6  (
            .in0(N__7646),
            .in1(N__8575),
            .in2(_gnd_net_),
            .in3(N__7538),
            .lcout(\uart_inst0.uart_inst0.rTxDataZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16910),
            .ce(N__8813),
            .sr(N__16436));
    defparam \uart_inst0.uart_inst0.rTxData_esr_6_LC_13_15_1 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rTxData_esr_6_LC_13_15_1 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rTxData_esr_6_LC_13_15_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uart_inst0.uart_inst0.rTxData_esr_6_LC_13_15_1  (
            .in0(N__7523),
            .in1(N__7606),
            .in2(_gnd_net_),
            .in3(N__8584),
            .lcout(\uart_inst0.uart_inst0.rTxDataZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16904),
            .ce(N__8806),
            .sr(N__16437));
    defparam \uart_inst0.uart_inst0.rTxData_esr_3_LC_13_15_3 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rTxData_esr_3_LC_13_15_3 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rTxData_esr_3_LC_13_15_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uart_inst0.uart_inst0.rTxData_esr_3_LC_13_15_3  (
            .in0(N__7667),
            .in1(N__8581),
            .in2(_gnd_net_),
            .in3(N__7514),
            .lcout(\uart_inst0.uart_inst0.rTxDataZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16904),
            .ce(N__8806),
            .sr(N__16437));
    defparam \uart_inst0.uart_inst0.rTxData_esr_4_LC_13_15_4 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rTxData_esr_4_LC_13_15_4 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rTxData_esr_4_LC_13_15_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uart_inst0.uart_inst0.rTxData_esr_4_LC_13_15_4  (
            .in0(N__8582),
            .in1(N__7625),
            .in2(_gnd_net_),
            .in3(N__7679),
            .lcout(\uart_inst0.uart_inst0.rTxDataZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16904),
            .ce(N__8806),
            .sr(N__16437));
    defparam \uart_inst0.uart_inst0.rTxData_esr_2_LC_13_15_5 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rTxData_esr_2_LC_13_15_5 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rTxData_esr_2_LC_13_15_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uart_inst0.uart_inst0.rTxData_esr_2_LC_13_15_5  (
            .in0(N__7661),
            .in1(N__8580),
            .in2(_gnd_net_),
            .in3(N__7655),
            .lcout(\uart_inst0.uart_inst0.rTxDataZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16904),
            .ce(N__8806),
            .sr(N__16437));
    defparam \uart_inst0.uart_inst0.rTxData_esr_5_LC_13_15_6 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rTxData_esr_5_LC_13_15_6 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rTxData_esr_5_LC_13_15_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \uart_inst0.uart_inst0.rTxData_esr_5_LC_13_15_6  (
            .in0(N__8583),
            .in1(N__7640),
            .in2(_gnd_net_),
            .in3(N__7634),
            .lcout(\uart_inst0.uart_inst0.rTxDataZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16904),
            .ce(N__8806),
            .sr(N__16437));
    defparam \uart_inst0.uart_inst0.rTxData_7_LC_13_16_2 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rTxData_7_LC_13_16_2 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rTxData_7_LC_13_16_2 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \uart_inst0.uart_inst0.rTxData_7_LC_13_16_2  (
            .in0(N__8562),
            .in1(N__7619),
            .in2(N__7610),
            .in3(N__8822),
            .lcout(\uart_inst0.uart_inst0.rTxDataZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16900),
            .ce(),
            .sr(N__16448));
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_3_LC_13_17_1 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_3_LC_13_17_1 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_3_LC_13_17_1 .LUT_INIT=16'b1011111111101010;
    LogicCell40 \uart_inst0.uart_inst0.tx_bits_remaining_3_LC_13_17_1  (
            .in0(N__8585),
            .in1(N__8777),
            .in2(N__8795),
            .in3(N__9766),
            .lcout(\uart_inst0.uart_inst0.tx_bits_remainingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16897),
            .ce(),
            .sr(N__16453));
    defparam \fifo_inst.ft2232h_inst.rFifoState_RNIM35O_0_LC_14_2_1 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rFifoState_RNIM35O_0_LC_14_2_1 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ft2232h_inst.rFifoState_RNIM35O_0_LC_14_2_1 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \fifo_inst.ft2232h_inst.rFifoState_RNIM35O_0_LC_14_2_1  (
            .in0(N__8117),
            .in1(N__8067),
            .in2(_gnd_net_),
            .in3(N__12750),
            .lcout(N_97),
            .ltout(N_97_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ft2232h_inst.rFifoState_0_LC_14_2_2 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rFifoState_0_LC_14_2_2 .SEQ_MODE=4'b1001;
    defparam \fifo_inst.ft2232h_inst.rFifoState_0_LC_14_2_2 .LUT_INIT=16'b1111001110110011;
    LogicCell40 \fifo_inst.ft2232h_inst.rFifoState_0_LC_14_2_2  (
            .in0(N__10609),
            .in1(N__8162),
            .in2(N__7595),
            .in3(N__10525),
            .lcout(fifo_inst_ft2232h_inst_rFifoState_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16972),
            .ce(),
            .sr(N__16351));
    defparam \uart_inst0.tx_uart_fifo_inst.m8_x0_LC_14_3_4 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m8_x0_LC_14_3_4 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m8_x0_LC_14_3_4 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m8_x0_LC_14_3_4  (
            .in0(N__7769),
            .in1(N__7709),
            .in2(N__7819),
            .in3(N__9237),
            .lcout(),
            .ltout(\uart_inst0.tx_uart_fifo_inst.m8_xZ0Z0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m8_ns_LC_14_3_5 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m8_ns_LC_14_3_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m8_ns_LC_14_3_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m8_ns_LC_14_3_5  (
            .in0(N__9238),
            .in1(_gnd_net_),
            .in2(N__7973),
            .in3(N__7734),
            .lcout(fifo_inst_tx_fifo_inst_wRamRdEn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rDataCount_fast_3_LC_14_3_6 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_fast_3_LC_14_3_6 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_fast_3_LC_14_3_6 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rDataCount_fast_3_LC_14_3_6  (
            .in0(N__7735),
            .in1(N__7970),
            .in2(N__7955),
            .in3(N__7873),
            .lcout(fifo_inst_tx_fifo_inst_rDataCount_fast_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16967),
            .ce(),
            .sr(N__16356));
    defparam \fifo_inst.tx_fifo_inst.rDataCount_0_LC_14_3_7 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_0_LC_14_3_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_0_LC_14_3_7 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \fifo_inst.tx_fifo_inst.rDataCount_0_LC_14_3_7  (
            .in0(N__7710),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7837),
            .lcout(fifo_inst_tx_fifo_inst_rDataCount_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16967),
            .ce(),
            .sr(N__16356));
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNO_1_2_LC_14_4_0 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNO_1_2_LC_14_4_0 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNO_1_2_LC_14_4_0 .LUT_INIT=16'b1010101011101010;
    LogicCell40 \fifo_inst.tx_fifo_inst.rDataCount_RNO_1_2_LC_14_4_0  (
            .in0(N__7934),
            .in1(N__7927),
            .in2(N__7877),
            .in3(N__9253),
            .lcout(),
            .ltout(\fifo_inst.tx_fifo_inst.un1_rDataCount_c2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rDataCount_2_LC_14_4_1 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_2_LC_14_4_1 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_2_LC_14_4_1 .LUT_INIT=16'b1010100101010110;
    LogicCell40 \fifo_inst.tx_fifo_inst.rDataCount_2_LC_14_4_1  (
            .in0(N__7814),
            .in1(N__7844),
            .in2(N__7847),
            .in3(N__9202),
            .lcout(fifo_inst_tx_fifo_inst_rDataCount_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16960),
            .ce(),
            .sr(N__16358));
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNO_0_2_LC_14_4_4 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNO_0_2_LC_14_4_4 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_RNO_0_2_LC_14_4_4 .LUT_INIT=16'b1010001000000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rDataCount_RNO_0_2_LC_14_4_4  (
            .in0(N__7771),
            .in1(N__9311),
            .in2(N__10178),
            .in3(N__9252),
            .lcout(\fifo_inst.tx_fifo_inst.un1_rDataCount_ac0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rDataCount_1_LC_14_4_5 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_1_LC_14_4_5 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rDataCount_1_LC_14_4_5 .LUT_INIT=16'b0011110010010110;
    LogicCell40 \fifo_inst.tx_fifo_inst.rDataCount_1_LC_14_4_5  (
            .in0(N__7719),
            .in1(N__9203),
            .in2(N__7785),
            .in3(N__7838),
            .lcout(fifo_inst_tx_fifo_inst_rDataCount_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16960),
            .ce(),
            .sr(N__16358));
    defparam \uart_inst0.tx_uart_fifo_inst.m7_LC_14_4_7 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m7_LC_14_4_7 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m7_LC_14_4_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m7_LC_14_4_7  (
            .in0(N__7813),
            .in1(N__7770),
            .in2(N__7739),
            .in3(N__7711),
            .lcout(N_8_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rDataCount_RNILHIG_0_LC_14_5_0 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.rDataCount_RNILHIG_0_LC_14_5_0 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.rx_fifo_inst.rDataCount_RNILHIG_0_LC_14_5_0 .LUT_INIT=16'b0100000000001010;
    LogicCell40 \fifo_inst.rx_fifo_inst.rDataCount_RNILHIG_0_LC_14_5_0  (
            .in0(N__15362),
            .in1(N__9076),
            .in2(N__12651),
            .in3(N__12593),
            .lcout(\fifo_inst.rx_fifo_inst.un1_rDataCount_axbxc3_1_1 ),
            .ltout(\fifo_inst.rx_fifo_inst.un1_rDataCount_axbxc3_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rDataCount_3_LC_14_5_1 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.rDataCount_3_LC_14_5_1 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rDataCount_3_LC_14_5_1 .LUT_INIT=16'b1110111110000000;
    LogicCell40 \fifo_inst.rx_fifo_inst.rDataCount_3_LC_14_5_1  (
            .in0(N__12687),
            .in1(N__12641),
            .in2(N__8051),
            .in3(N__12749),
            .lcout(fifo_inst_wRxWrFull),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16953),
            .ce(),
            .sr(N__16367));
    defparam \fifo_inst.ft2232h_inst.rRxWrEn_LC_14_5_3 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rRxWrEn_LC_14_5_3 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rRxWrEn_LC_14_5_3 .LUT_INIT=16'b1100110011101110;
    LogicCell40 \fifo_inst.ft2232h_inst.rRxWrEn_LC_14_5_3  (
            .in0(N__9077),
            .in1(N__17028),
            .in2(_gnd_net_),
            .in3(N__8146),
            .lcout(fifo_inst_wRxWrEn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16953),
            .ce(),
            .sr(N__16367));
    defparam \uart_inst0.tx_uart_fifo_inst.m15_x0_LC_14_5_4 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m15_x0_LC_14_5_4 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m15_x0_LC_14_5_4 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m15_x0_LC_14_5_4  (
            .in0(N__12586),
            .in1(N__12686),
            .in2(N__15377),
            .in3(N__8220),
            .lcout(),
            .ltout(\uart_inst0.tx_uart_fifo_inst.m15_xZ0Z0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m15_ns_LC_14_5_5 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m15_ns_LC_14_5_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m15_ns_LC_14_5_5 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m15_ns_LC_14_5_5  (
            .in0(_gnd_net_),
            .in1(N__8034),
            .in2(N__8048),
            .in3(N__15361),
            .lcout(fifo_inst_rx_fifo_inst_wRamRdEn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rDataCount_fast_3_LC_14_5_6 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.rDataCount_fast_3_LC_14_5_6 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rDataCount_fast_3_LC_14_5_6 .LUT_INIT=16'b1110101010100010;
    LogicCell40 \fifo_inst.rx_fifo_inst.rDataCount_fast_3_LC_14_5_6  (
            .in0(N__8035),
            .in1(N__8045),
            .in2(N__12652),
            .in3(N__12688),
            .lcout(fifo_inst_rx_fifo_inst_rDataCount_fast_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16953),
            .ce(),
            .sr(N__16367));
    defparam \fifo_inst.ft2232h_inst.rFifoState_4_LC_14_6_0 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rFifoState_4_LC_14_6_0 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rFifoState_4_LC_14_6_0 .LUT_INIT=16'b1111111100001010;
    LogicCell40 \fifo_inst.ft2232h_inst.rFifoState_4_LC_14_6_0  (
            .in0(N__9160),
            .in1(_gnd_net_),
            .in2(N__9188),
            .in3(N__8256),
            .lcout(fifo_inst_ft2232h_inst_rFifoState_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16947),
            .ce(),
            .sr(N__16385));
    defparam rRxEn_LC_14_6_1.C_ON=1'b0;
    defparam rRxEn_LC_14_6_1.SEQ_MODE=4'b1000;
    defparam rRxEn_LC_14_6_1.LUT_INIT=16'b0001000100010001;
    LogicCell40 rRxEn_LC_14_6_1 (
            .in0(N__8200),
            .in1(N__8179),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(P1A2_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16947),
            .ce(),
            .sr(N__16385));
    defparam \fifo_inst.ft2232h_inst.rWrDelay_LC_14_6_3 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rWrDelay_LC_14_6_3 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rWrDelay_LC_14_6_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \fifo_inst.ft2232h_inst.rWrDelay_LC_14_6_3  (
            .in0(_gnd_net_),
            .in1(N__9183),
            .in2(_gnd_net_),
            .in3(N__9159),
            .lcout(fifo_inst_ft2232h_inst_rWrDelay),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16947),
            .ce(),
            .sr(N__16385));
    defparam \fifo_inst.ft2232h_inst.rTx_n_LC_14_6_4 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rTx_n_LC_14_6_4 .SEQ_MODE=4'b1001;
    defparam \fifo_inst.ft2232h_inst.rTx_n_LC_14_6_4 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \fifo_inst.ft2232h_inst.rTx_n_LC_14_6_4  (
            .in0(N__7989),
            .in1(N__8257),
            .in2(_gnd_net_),
            .in3(N__10672),
            .lcout(P1A4_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16947),
            .ce(),
            .sr(N__16385));
    defparam \fifo_inst.rx_fifo_inst.rDataCount_0_LC_14_6_5 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.rDataCount_0_LC_14_6_5 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rDataCount_0_LC_14_6_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \fifo_inst.rx_fifo_inst.rDataCount_0_LC_14_6_5  (
            .in0(_gnd_net_),
            .in1(N__8235),
            .in2(_gnd_net_),
            .in3(N__12645),
            .lcout(fifo_inst_rx_fifo_inst_rDataCount_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16947),
            .ce(),
            .sr(N__16385));
    defparam \fifo_inst.ft2232h_inst.rFifoState_3_LC_14_6_6 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rFifoState_3_LC_14_6_6 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rFifoState_3_LC_14_6_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \fifo_inst.ft2232h_inst.rFifoState_3_LC_14_6_6  (
            .in0(N__10600),
            .in1(N__10658),
            .in2(_gnd_net_),
            .in3(N__10530),
            .lcout(fifo_inst_ft2232h_inst_rFifoState_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16947),
            .ce(),
            .sr(N__16385));
    defparam \fifo_inst.rx_fifo_inst.rDataCount_fast_0_LC_14_6_7 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.rDataCount_fast_0_LC_14_6_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rDataCount_fast_0_LC_14_6_7 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \fifo_inst.rx_fifo_inst.rDataCount_fast_0_LC_14_6_7  (
            .in0(_gnd_net_),
            .in1(N__8236),
            .in2(_gnd_net_),
            .in3(N__8222),
            .lcout(fifo_inst_rx_fifo_inst_rDataCount_fast_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16947),
            .ce(),
            .sr(N__16385));
    defparam rFtdiRxState_0_LC_14_7_0.C_ON=1'b0;
    defparam rFtdiRxState_0_LC_14_7_0.SEQ_MODE=4'b1000;
    defparam rFtdiRxState_0_LC_14_7_0.LUT_INIT=16'b0000010100000000;
    LogicCell40 rFtdiRxState_0_LC_14_7_0 (
            .in0(N__8204),
            .in1(_gnd_net_),
            .in2(N__8180),
            .in3(N__14015),
            .lcout(rFtdiRxStateZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16942),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNID3RQ_3_LC_14_7_2 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNID3RQ_3_LC_14_7_2 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNID3RQ_3_LC_14_7_2 .LUT_INIT=16'b0000000011101110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rDataCount_RNID3RQ_3_LC_14_7_2  (
            .in0(N__11216),
            .in1(N__15368),
            .in2(_gnd_net_),
            .in3(N__8317),
            .lcout(),
            .ltout(rUartTxEn_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNI9H5T_3_LC_14_7_3 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNI9H5T_3_LC_14_7_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNI9H5T_3_LC_14_7_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rDataCount_RNI9H5T_3_LC_14_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8183),
            .in3(N__16674),
            .lcout(rUartTxEn_4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m27_e_LC_14_7_5 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m27_e_LC_14_7_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m27_e_LC_14_7_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m27_e_LC_14_7_5  (
            .in0(N__14016),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8175),
            .lcout(N_27_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ft2232h_inst.rFifoState_RNO_0_0_LC_14_8_4 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rFifoState_RNO_0_0_LC_14_8_4 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ft2232h_inst.rFifoState_RNO_0_0_LC_14_8_4 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \fifo_inst.ft2232h_inst.rFifoState_RNO_0_0_LC_14_8_4  (
            .in0(N__8133),
            .in1(N__9187),
            .in2(_gnd_net_),
            .in3(N__9161),
            .lcout(\fifo_inst.ft2232h_inst.rFifoStatesr_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ft2232h_inst.rFifoState_2_LC_14_9_3 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rFifoState_2_LC_14_9_3 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rFifoState_2_LC_14_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.ft2232h_inst.rFifoState_2_LC_14_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17027),
            .lcout(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16933),
            .ce(),
            .sr(N__16416));
    defparam \fifo_inst.ft2232h_inst.rFifoState_1_LC_14_9_4 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rFifoState_1_LC_14_9_4 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rFifoState_1_LC_14_9_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \fifo_inst.ft2232h_inst.rFifoState_1_LC_14_9_4  (
            .in0(N__8103),
            .in1(N__8077),
            .in2(_gnd_net_),
            .in3(N__12762),
            .lcout(\fifo_inst.ft2232h_inst.rFifoStateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16933),
            .ce(),
            .sr(N__16416));
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCountZ0Z_1_LC_14_9_7 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCountZ0Z_1_LC_14_9_7 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCountZ0Z_1_LC_14_9_7 .LUT_INIT=16'b1011010001111000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rDataCountZ0Z_1_LC_14_9_7  (
            .in0(N__8476),
            .in1(N__8355),
            .in2(N__8429),
            .in3(N__9591),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rDataCountZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16933),
            .ce(),
            .sr(N__16416));
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNO_0_2_LC_14_10_0 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNO_0_2_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNO_0_2_LC_14_10_0 .LUT_INIT=16'b0100101000001000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rDataCount_RNO_0_2_LC_14_10_0  (
            .in0(N__9489),
            .in1(N__8408),
            .in2(N__8509),
            .in3(N__8350),
            .lcout(\uart_inst0.tx_uart_fifo_inst.un1_rDataCount_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNO_0_1_LC_14_10_3 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNO_0_1_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNO_0_1_LC_14_10_3 .LUT_INIT=16'b1010101010011010;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rDataCount_RNO_0_1_LC_14_10_3  (
            .in0(N__8409),
            .in1(N__9832),
            .in2(N__9506),
            .in3(N__8492),
            .lcout(\uart_inst0.tx_uart_fifo_inst.un1_rDataCount_axbxc1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIJHQM1_2_LC_14_10_6 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIJHQM1_2_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIJHQM1_2_LC_14_10_6 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIJHQM1_2_LC_14_10_6  (
            .in0(N__9487),
            .in1(N__8407),
            .in2(N__8386),
            .in3(N__8349),
            .lcout(),
            .ltout(\uart_inst0.tx_uart_fifo_inst.rDataCount_RNIJHQM1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIKKMI2_3_LC_14_10_7 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIKKMI2_3_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIKKMI2_3_LC_14_10_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rDataCount_RNIKKMI2_3_LC_14_10_7  (
            .in0(_gnd_net_),
            .in1(N__9488),
            .in2(N__8321),
            .in3(N__8300),
            .lcout(\uart_inst0.tx_uart_fifo_inst.wRamRdEn_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIBDOK2_0_LC_14_11_0 .C_ON=1'b1;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIBDOK2_0_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIBDOK2_0_LC_14_11_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIBDOK2_0_LC_14_11_0  (
            .in0(_gnd_net_),
            .in1(N__9415),
            .in2(N__9592),
            .in3(N__9587),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIBDOK2Z0Z_0 ),
            .ltout(),
            .carryin(bfn_14_11_0_),
            .carryout(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIOA54_LC_14_11_1 .C_ON=1'b1;
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIOA54_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIOA54_LC_14_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIOA54_LC_14_11_1  (
            .in0(_gnd_net_),
            .in1(N__11315),
            .in2(_gnd_net_),
            .in3(N__8267),
            .lcout(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIOAZ0Z54 ),
            .ltout(),
            .carryin(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_0 ),
            .carryout(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIQD64_LC_14_11_2 .C_ON=1'b1;
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIQD64_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIQD64_LC_14_11_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIQD64_LC_14_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11300),
            .in3(N__8264),
            .lcout(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIQDZ0Z64 ),
            .ltout(),
            .carryin(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_1 ),
            .carryout(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNISG74_LC_14_11_3 .C_ON=1'b1;
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNISG74_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNISG74_LC_14_11_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNISG74_LC_14_11_3  (
            .in0(_gnd_net_),
            .in1(N__9403),
            .in2(_gnd_net_),
            .in3(N__8261),
            .lcout(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNISGZ0Z74 ),
            .ltout(),
            .carryin(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_2 ),
            .carryout(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIUJ84_LC_14_11_4 .C_ON=1'b1;
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIUJ84_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIUJ84_LC_14_11_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIUJ84_LC_14_11_4  (
            .in0(_gnd_net_),
            .in1(N__9709),
            .in2(_gnd_net_),
            .in3(N__8762),
            .lcout(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIUJZ0Z84 ),
            .ltout(),
            .carryin(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_3 ),
            .carryout(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNI0N94_LC_14_11_5 .C_ON=1'b1;
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNI0N94_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNI0N94_LC_14_11_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNI0N94_LC_14_11_5  (
            .in0(_gnd_net_),
            .in1(N__9694),
            .in2(_gnd_net_),
            .in3(N__8759),
            .lcout(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNI0NZ0Z94 ),
            .ltout(),
            .carryin(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_4 ),
            .carryout(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNI2QA4_LC_14_11_6 .C_ON=1'b1;
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNI2QA4_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNI2QA4_LC_14_11_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNI2QA4_LC_14_11_6  (
            .in0(_gnd_net_),
            .in1(N__9667),
            .in2(_gnd_net_),
            .in3(N__8756),
            .lcout(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNI2QAZ0Z4 ),
            .ltout(),
            .carryin(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_5 ),
            .carryout(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI4TB4_LC_14_11_7 .C_ON=1'b1;
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI4TB4_LC_14_11_7 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI4TB4_LC_14_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI4TB4_LC_14_11_7  (
            .in0(_gnd_net_),
            .in1(N__9634),
            .in2(_gnd_net_),
            .in3(N__8753),
            .lcout(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI4TBZ0Z4 ),
            .ltout(),
            .carryin(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_6 ),
            .carryout(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI60D4_LC_14_12_0 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI60D4_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI60D4_LC_14_12_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI60D4_LC_14_12_0  (
            .in0(_gnd_net_),
            .in1(N__9611),
            .in2(_gnd_net_),
            .in3(N__8750),
            .lcout(\uart_inst0.tx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI60DZ0Z4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNIU317_4_LC_14_12_6 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNIU317_4_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNIU317_4_LC_14_12_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamWrAddr_RNIU317_4_LC_14_12_6  (
            .in0(N__8743),
            .in1(N__8713),
            .in2(N__8692),
            .in3(N__8662),
            .lcout(\uart_inst0.tx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rTx_LC_14_14_5 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rTx_LC_14_14_5 .SEQ_MODE=4'b1001;
    defparam \uart_inst0.uart_inst0.rTx_LC_14_14_5 .LUT_INIT=16'b0011000001110100;
    LogicCell40 \uart_inst0.uart_inst0.rTx_LC_14_14_5  (
            .in0(N__8579),
            .in1(N__8828),
            .in2(N__8602),
            .in3(N__8528),
            .lcout(P1A7_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16914),
            .ce(),
            .sr(N__16438));
    defparam \uart_inst0.uart_inst0.tx_state_RNI5LM6_0_LC_14_15_4 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_state_RNI5LM6_0_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_state_RNI5LM6_0_LC_14_15_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uart_inst0.uart_inst0.tx_state_RNI5LM6_0_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(N__11565),
            .in2(_gnd_net_),
            .in3(N__11660),
            .lcout(\uart_inst0.uart_inst0.tx_state_81_d ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rTx_RNO_1_LC_14_15_6 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rTx_RNO_1_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rTx_RNO_1_LC_14_15_6 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \uart_inst0.uart_inst0.rTx_RNO_1_LC_14_15_6  (
            .in0(N__11861),
            .in1(N__8534),
            .in2(_gnd_net_),
            .in3(N__9988),
            .lcout(\uart_inst0.uart_inst0.rTx_6_f1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rTx_RNO_0_LC_14_15_7 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rTx_RNO_0_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rTx_RNO_0_LC_14_15_7 .LUT_INIT=16'b0101101000001010;
    LogicCell40 \uart_inst0.uart_inst0.rTx_RNO_0_LC_14_15_7  (
            .in0(N__11661),
            .in1(_gnd_net_),
            .in2(N__11582),
            .in3(N__11860),
            .lcout(\uart_inst0.uart_inst0.N_141_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_state_RNI9VFM2_0_LC_14_16_1 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_state_RNI9VFM2_0_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_state_RNI9VFM2_0_LC_14_16_1 .LUT_INIT=16'b0001101000001010;
    LogicCell40 \uart_inst0.uart_inst0.tx_state_RNI9VFM2_0_LC_14_16_1  (
            .in0(N__11648),
            .in1(N__9748),
            .in2(N__11579),
            .in3(N__11853),
            .lcout(\uart_inst0.uart_inst0.N_143_0 ),
            .ltout(\uart_inst0.uart_inst0.N_143_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_state_RNI5DQO2_0_LC_14_16_2 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_state_RNI5DQO2_0_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_state_RNI5DQO2_0_LC_14_16_2 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \uart_inst0.uart_inst0.tx_state_RNI5DQO2_0_LC_14_16_2  (
            .in0(N__14068),
            .in1(_gnd_net_),
            .in2(N__8816),
            .in3(_gnd_net_),
            .lcout(\uart_inst0.uart_inst0.N_143_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_RNO_0_3_LC_14_16_4 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_RNO_0_3_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_RNO_0_3_LC_14_16_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart_inst0.uart_inst0.tx_bits_remaining_RNO_0_3_LC_14_16_4  (
            .in0(N__9928),
            .in1(N__9792),
            .in2(_gnd_net_),
            .in3(N__9956),
            .lcout(\uart_inst0.uart_inst0.un1_m3_0_a2_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_RNO_0_1_LC_14_16_5 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_RNO_0_1_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_RNO_0_1_LC_14_16_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uart_inst0.uart_inst0.tx_bits_remaining_RNO_0_1_LC_14_16_5  (
            .in0(N__11650),
            .in1(N__11855),
            .in2(N__11580),
            .in3(N__9927),
            .lcout(\uart_inst0.uart_inst0.un1_tx_bits_remaining_c1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_state_RNI9VFM2_0_0_LC_14_16_6 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_state_RNI9VFM2_0_0_LC_14_16_6 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_state_RNI9VFM2_0_0_LC_14_16_6 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \uart_inst0.uart_inst0.tx_state_RNI9VFM2_0_0_LC_14_16_6  (
            .in0(N__11854),
            .in1(N__11556),
            .in2(N__9752),
            .in3(N__11649),
            .lcout(\uart_inst0.uart_inst0.N_136_0 ),
            .ltout(\uart_inst0.uart_inst0.N_136_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_0_LC_14_16_7 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_0_LC_14_16_7 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_0_LC_14_16_7 .LUT_INIT=16'b0000001100110000;
    LogicCell40 \uart_inst0.uart_inst0.tx_bits_remaining_0_LC_14_16_7  (
            .in0(_gnd_net_),
            .in1(N__9970),
            .in2(N__8786),
            .in3(N__9929),
            .lcout(\uart_inst0.uart_inst0.tx_bits_remainingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16905),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_1_LC_14_17_0 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_1_LC_14_17_0 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_1_LC_14_17_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.uart_inst0.tx_bits_remaining_1_LC_14_17_0  (
            .in0(N__8783),
            .in1(N__8775),
            .in2(_gnd_net_),
            .in3(N__9957),
            .lcout(\uart_inst0.uart_inst0.tx_bits_remainingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16901),
            .ce(),
            .sr(N__9977));
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_2_LC_14_17_6 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_2_LC_14_17_6 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_2_LC_14_17_6 .LUT_INIT=16'b1110000101011010;
    LogicCell40 \uart_inst0.uart_inst0.tx_bits_remaining_2_LC_14_17_6  (
            .in0(N__9902),
            .in1(N__9958),
            .in2(N__9797),
            .in3(N__8776),
            .lcout(\uart_inst0.uart_inst0.tx_bits_remainingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16901),
            .ce(),
            .sr(N__9977));
    defparam \uart_inst0.uart_inst0.tx_countdown_0_LC_14_18_1 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_countdown_0_LC_14_18_1 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.tx_countdown_0_LC_14_18_1 .LUT_INIT=16'b1001100110101010;
    LogicCell40 \uart_inst0.uart_inst0.tx_countdown_0_LC_14_18_1  (
            .in0(N__14548),
            .in1(N__11875),
            .in2(_gnd_net_),
            .in3(N__10198),
            .lcout(\uart_inst0.uart_inst0.tx_countdownZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16898),
            .ce(),
            .sr(N__13591));
    defparam \uart_inst0.uart_inst0.tx_countdown_1_LC_14_18_6 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_countdown_1_LC_14_18_6 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.tx_countdown_1_LC_14_18_6 .LUT_INIT=16'b1100110011000110;
    LogicCell40 \uart_inst0.uart_inst0.tx_countdown_1_LC_14_18_6  (
            .in0(N__10199),
            .in1(N__14591),
            .in2(N__11879),
            .in3(N__14549),
            .lcout(\uart_inst0.uart_inst0.tx_countdownZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16898),
            .ce(),
            .sr(N__13591));
    defparam \fifo_inst.tx_fifo_inst.ram512x8_inst.RDATA_0_LC_15_1_4 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.ram512x8_inst.RDATA_0_LC_15_1_4 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.ram512x8_inst.RDATA_0_LC_15_1_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.ram512x8_inst.RDATA_0_LC_15_1_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8858),
            .lcout(wTxRdData_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVfifo_inst.tx_fifo_inst.ram512x8_inst.RDATA_0C_net ),
            .ce(N__10276),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_6_LC_15_2_2 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_6_LC_15_2_2 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_6_LC_15_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_6_LC_15_2_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8941),
            .lcout(fifo_inst_tx_fifo_inst_rRamRdAddr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16975),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_5_LC_15_2_6 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_5_LC_15_2_6 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_5_LC_15_2_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_5_LC_15_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8965),
            .lcout(fifo_inst_tx_fifo_inst_rRamRdAddr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16975),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_7_LC_15_2_7 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_7_LC_15_2_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_7_LC_15_2_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_7_LC_15_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8917),
            .lcout(fifo_inst_tx_fifo_inst_rRamRdAddr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16975),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNI9KL42_0_LC_15_3_0 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNI9KL42_0_LC_15_3_0 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_RNI9KL42_0_LC_15_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_RNI9KL42_0_LC_15_3_0  (
            .in0(_gnd_net_),
            .in1(N__10214),
            .in2(N__10275),
            .in3(N__10265),
            .lcout(rRamRdAddr_RNI9KL42_0),
            .ltout(),
            .carryin(bfn_15_3_0_),
            .carryout(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIE7TP_LC_15_3_1 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIE7TP_LC_15_3_1 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIE7TP_LC_15_3_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIE7TP_LC_15_3_1  (
            .in0(N__16628),
            .in1(N__10349),
            .in2(_gnd_net_),
            .in3(N__8834),
            .lcout(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIE7TPZ0 ),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_0 ),
            .carryout(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIGAUP_LC_15_3_2 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIGAUP_LC_15_3_2 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIGAUP_LC_15_3_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIGAUP_LC_15_3_2  (
            .in0(N__16631),
            .in1(N__12779),
            .in2(_gnd_net_),
            .in3(N__8831),
            .lcout(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIGAUPZ0 ),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_1 ),
            .carryout(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_2_c_RNIMVKN_LC_15_3_3 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_2_c_RNIMVKN_LC_15_3_3 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_2_c_RNIMVKN_LC_15_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_2_c_RNIMVKN_LC_15_3_3  (
            .in0(_gnd_net_),
            .in1(N__10361),
            .in2(_gnd_net_),
            .in3(N__8981),
            .lcout(un1_rRamRdAddr_cry_2_c_RNIMVKN),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_2 ),
            .carryout(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIKG0Q_LC_15_3_4 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIKG0Q_LC_15_3_4 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIKG0Q_LC_15_3_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIKG0Q_LC_15_3_4  (
            .in0(N__16632),
            .in1(N__10292),
            .in2(_gnd_net_),
            .in3(N__8978),
            .lcout(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIKG0QZ0 ),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_3 ),
            .carryout(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIMJ1Q_LC_15_3_5 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIMJ1Q_LC_15_3_5 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIMJ1Q_LC_15_3_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIMJ1Q_LC_15_3_5  (
            .in0(N__16629),
            .in1(N__10418),
            .in2(_gnd_net_),
            .in3(N__8954),
            .lcout(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIMJ1QZ0 ),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_4 ),
            .carryout(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIOM2Q_LC_15_3_6 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIOM2Q_LC_15_3_6 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIOM2Q_LC_15_3_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIOM2Q_LC_15_3_6  (
            .in0(N__16633),
            .in1(N__10393),
            .in2(_gnd_net_),
            .in3(N__8930),
            .lcout(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIOM2QZ0 ),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_5 ),
            .carryout(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIQP3Q_LC_15_3_7 .C_ON=1'b1;
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIQP3Q_LC_15_3_7 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIQP3Q_LC_15_3_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIQP3Q_LC_15_3_7  (
            .in0(N__16630),
            .in1(N__10406),
            .in2(_gnd_net_),
            .in3(N__8906),
            .lcout(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIQP3QZ0 ),
            .ltout(),
            .carryin(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_6 ),
            .carryout(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNISS4Q_LC_15_4_0 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNISS4Q_LC_15_4_0 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNISS4Q_LC_15_4_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNISS4Q_LC_15_4_0  (
            .in0(N__16649),
            .in1(N__10333),
            .in2(_gnd_net_),
            .in3(N__8903),
            .lcout(\fifo_inst.tx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNISS4QZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_1_LC_15_4_1 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_1_LC_15_4_1 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_1_LC_15_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_1_LC_15_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8890),
            .lcout(fifo_inst_tx_fifo_inst_rRamRdAddr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16968),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_2_LC_15_4_2 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_2_LC_15_4_2 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_2_LC_15_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.rx_fifo_inst.rRamRdAddr_2_LC_15_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9031),
            .lcout(fifo_inst_rx_fifo_inst_rRamRdAddr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16968),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_8_LC_15_4_3 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_8_LC_15_4_3 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_8_LC_15_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_8_LC_15_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8869),
            .lcout(fifo_inst_tx_fifo_inst_rRamRdAddr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16968),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_6_LC_15_4_5 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_6_LC_15_4_5 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_6_LC_15_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.rx_fifo_inst.rRamRdAddr_6_LC_15_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8995),
            .lcout(fifo_inst_rx_fifo_inst_rRamRdAddr_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16968),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m12_LC_15_4_7 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m12_LC_15_4_7 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m12_LC_15_4_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m12_LC_15_4_7  (
            .in0(_gnd_net_),
            .in1(N__12725),
            .in2(_gnd_net_),
            .in3(N__9071),
            .lcout(fifo_inst_rx_fifo_inst_wRamWrEn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_RNI0S8U_0_LC_15_5_0 .C_ON=1'b1;
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_RNI0S8U_0_LC_15_5_0 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_RNI0S8U_0_LC_15_5_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \fifo_inst.rx_fifo_inst.rRamRdAddr_RNI0S8U_0_LC_15_5_0  (
            .in0(_gnd_net_),
            .in1(N__10913),
            .in2(N__10954),
            .in3(N__10942),
            .lcout(rRamRdAddr_RNI0S8U_0),
            .ltout(),
            .carryin(bfn_15_5_0_),
            .carryout(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIAHVB_LC_15_5_1 .C_ON=1'b1;
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIAHVB_LC_15_5_1 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIAHVB_LC_15_5_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIAHVB_LC_15_5_1  (
            .in0(N__16660),
            .in1(N__10700),
            .in2(_gnd_net_),
            .in3(N__9044),
            .lcout(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIAHVBZ0 ),
            .ltout(),
            .carryin(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_0 ),
            .carryout(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNICK0C_LC_15_5_2 .C_ON=1'b1;
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNICK0C_LC_15_5_2 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNICK0C_LC_15_5_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNICK0C_LC_15_5_2  (
            .in0(N__16663),
            .in1(N__11044),
            .in2(_gnd_net_),
            .in3(N__9020),
            .lcout(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_1_c_RNICK0CZ0 ),
            .ltout(),
            .carryin(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_1 ),
            .carryout(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_2_c_RNII9N9_LC_15_5_3 .C_ON=1'b1;
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_2_c_RNII9N9_LC_15_5_3 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_2_c_RNII9N9_LC_15_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_2_c_RNII9N9_LC_15_5_3  (
            .in0(_gnd_net_),
            .in1(N__10712),
            .in2(_gnd_net_),
            .in3(N__9017),
            .lcout(un1_rRamRdAddr_cry_2_c_RNII9N9),
            .ltout(),
            .carryin(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_2 ),
            .carryout(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIGQ2C_LC_15_5_4 .C_ON=1'b1;
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIGQ2C_LC_15_5_4 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIGQ2C_LC_15_5_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIGQ2C_LC_15_5_4  (
            .in0(N__16664),
            .in1(N__11063),
            .in2(_gnd_net_),
            .in3(N__9014),
            .lcout(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIGQ2CZ0 ),
            .ltout(),
            .carryin(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_3 ),
            .carryout(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIIT3C_LC_15_5_5 .C_ON=1'b1;
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIIT3C_LC_15_5_5 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIIT3C_LC_15_5_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIIT3C_LC_15_5_5  (
            .in0(N__16661),
            .in1(N__11077),
            .in2(_gnd_net_),
            .in3(N__9011),
            .lcout(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_4_c_RNIIT3CZ0 ),
            .ltout(),
            .carryin(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_4 ),
            .carryout(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIK05C_LC_15_5_6 .C_ON=1'b1;
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIK05C_LC_15_5_6 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIK05C_LC_15_5_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIK05C_LC_15_5_6  (
            .in0(N__16665),
            .in1(N__11018),
            .in2(_gnd_net_),
            .in3(N__8984),
            .lcout(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIK05CZ0 ),
            .ltout(),
            .carryin(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_5 ),
            .carryout(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIM36C_LC_15_5_7 .C_ON=1'b1;
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIM36C_LC_15_5_7 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIM36C_LC_15_5_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIM36C_LC_15_5_7  (
            .in0(N__16662),
            .in1(N__11032),
            .in2(_gnd_net_),
            .in3(N__9338),
            .lcout(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_6_c_RNIM36CZ0 ),
            .ltout(),
            .carryin(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_6 ),
            .carryout(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNIO67C_LC_15_6_0 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNIO67C_LC_15_6_0 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNIO67C_LC_15_6_0 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNIO67C_LC_15_6_0  (
            .in0(N__10687),
            .in1(N__16670),
            .in2(_gnd_net_),
            .in3(N__9335),
            .lcout(\fifo_inst.rx_fifo_inst.un1_rRamRdAddr_cry_7_c_RNIO67CZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_5_LC_15_6_1 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_5_LC_15_6_1 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_5_LC_15_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.rx_fifo_inst.rRamRdAddr_5_LC_15_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9322),
            .lcout(fifo_inst_rx_fifo_inst_rRamRdAddr_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16954),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m10_LC_15_6_3 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m10_LC_15_6_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m10_LC_15_6_3 .LUT_INIT=16'b1000000010110000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m10_LC_15_6_3  (
            .in0(N__10174),
            .in1(N__9310),
            .in2(N__9263),
            .in3(N__10526),
            .lcout(fifo_inst_tx_fifo_inst_rDataCount_0_sqmuxa),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m23_LC_15_6_6 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m23_LC_15_6_6 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m23_LC_15_6_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m23_LC_15_6_6  (
            .in0(_gnd_net_),
            .in1(N__9179),
            .in2(_gnd_net_),
            .in3(N__9155),
            .lcout(N_101),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_8_LC_15_6_7 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_8_LC_15_6_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_8_LC_15_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.rx_fifo_inst.rRamRdAddr_8_LC_15_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9127),
            .lcout(fifo_inst_rx_fifo_inst_rRamRdAddr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16954),
            .ce(),
            .sr(_gnd_net_));
    defparam rUartTxData_ess_6_LC_15_7_0.C_ON=1'b0;
    defparam rUartTxData_ess_6_LC_15_7_0.SEQ_MODE=4'b1001;
    defparam rUartTxData_ess_6_LC_15_7_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 rUartTxData_ess_6_LC_15_7_0 (
            .in0(N__9380),
            .in1(N__12548),
            .in2(_gnd_net_),
            .in3(N__11230),
            .lcout(rUartTxDataZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16948),
            .ce(N__11179),
            .sr(N__16414));
    defparam rUartTxData_esr_5_LC_15_7_1.C_ON=1'b0;
    defparam rUartTxData_esr_5_LC_15_7_1.SEQ_MODE=4'b1000;
    defparam rUartTxData_esr_5_LC_15_7_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 rUartTxData_esr_5_LC_15_7_1 (
            .in0(N__11229),
            .in1(N__9386),
            .in2(_gnd_net_),
            .in3(N__12872),
            .lcout(rUartTxDataZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16948),
            .ce(N__11179),
            .sr(N__16414));
    defparam rUartTxData_esr_1_LC_15_7_4.C_ON=1'b0;
    defparam rUartTxData_esr_1_LC_15_7_4.SEQ_MODE=4'b1000;
    defparam rUartTxData_esr_1_LC_15_7_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 rUartTxData_esr_1_LC_15_7_4 (
            .in0(N__9374),
            .in1(N__12536),
            .in2(_gnd_net_),
            .in3(N__11228),
            .lcout(rUartTxDataZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16948),
            .ce(N__11179),
            .sr(N__16414));
    defparam rUartRxData_esr_5_LC_15_8_0.C_ON=1'b0;
    defparam rUartRxData_esr_5_LC_15_8_0.SEQ_MODE=4'b1000;
    defparam rUartRxData_esr_5_LC_15_8_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 rUartRxData_esr_5_LC_15_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15008),
            .lcout(rUartRxDataZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16943),
            .ce(N__11167),
            .sr(N__16417));
    defparam rUartRxData_esr_7_LC_15_8_5.C_ON=1'b0;
    defparam rUartRxData_esr_7_LC_15_8_5.SEQ_MODE=4'b1000;
    defparam rUartRxData_esr_7_LC_15_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 rUartRxData_esr_7_LC_15_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14894),
            .lcout(rUartRxDataZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16943),
            .ce(N__11167),
            .sr(N__16417));
    defparam rUartRxData_esr_6_LC_15_8_6.C_ON=1'b0;
    defparam rUartRxData_esr_6_LC_15_8_6.SEQ_MODE=4'b1000;
    defparam rUartRxData_esr_6_LC_15_8_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 rUartRxData_esr_6_LC_15_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14984),
            .lcout(rUartRxDataZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16943),
            .ce(N__11167),
            .sr(N__16417));
    defparam rUartRxData_esr_2_LC_15_9_0.C_ON=1'b0;
    defparam rUartRxData_esr_2_LC_15_9_0.SEQ_MODE=4'b1000;
    defparam rUartRxData_esr_2_LC_15_9_0.LUT_INIT=16'b1100110011001100;
    LogicCell40 rUartRxData_esr_2_LC_15_9_0 (
            .in0(_gnd_net_),
            .in1(N__15551),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(rUartRxDataZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16939),
            .ce(N__11168),
            .sr(N__16420));
    defparam rUartRxData_esr_0_LC_15_9_2.C_ON=1'b0;
    defparam rUartRxData_esr_0_LC_15_9_2.SEQ_MODE=4'b1000;
    defparam rUartRxData_esr_0_LC_15_9_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 rUartRxData_esr_0_LC_15_9_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14864),
            .lcout(rUartRxDataZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16939),
            .ce(N__11168),
            .sr(N__16420));
    defparam rUartRxData_esr_3_LC_15_9_3.C_ON=1'b0;
    defparam rUartRxData_esr_3_LC_15_9_3.SEQ_MODE=4'b1000;
    defparam rUartRxData_esr_3_LC_15_9_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 rUartRxData_esr_3_LC_15_9_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15536),
            .lcout(rUartRxDataZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16939),
            .ce(N__11168),
            .sr(N__16420));
    defparam rUartRxData_esr_4_LC_15_9_4.C_ON=1'b0;
    defparam rUartRxData_esr_4_LC_15_9_4.SEQ_MODE=4'b1000;
    defparam rUartRxData_esr_4_LC_15_9_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 rUartRxData_esr_4_LC_15_9_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15521),
            .lcout(rUartRxDataZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16939),
            .ce(N__11168),
            .sr(N__16420));
    defparam rUartRxData_esr_1_LC_15_9_5.C_ON=1'b0;
    defparam rUartRxData_esr_1_LC_15_9_5.SEQ_MODE=4'b1000;
    defparam rUartRxData_esr_1_LC_15_9_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 rUartRxData_esr_1_LC_15_9_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15566),
            .lcout(rUartRxDataZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16939),
            .ce(N__11168),
            .sr(N__16420));
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_2_LC_15_10_1 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_2_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_2_LC_15_10_1 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_2_LC_15_10_1  (
            .in0(N__16676),
            .in1(N__9522),
            .in2(N__9350),
            .in3(N__9589),
            .lcout(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_3_LC_15_10_2 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_3_LC_15_10_2 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_3_LC_15_10_2 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_3_LC_15_10_2  (
            .in0(N__9590),
            .in1(N__9349),
            .in2(_gnd_net_),
            .in3(N__9526),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16934),
            .ce(),
            .sr(N__13600));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIIP78_4_LC_15_10_3 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIIP78_4_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIIP78_4_LC_15_10_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIIP78_4_LC_15_10_3  (
            .in0(N__9671),
            .in1(N__9698),
            .in2(N__9644),
            .in3(N__9713),
            .lcout(),
            .ltout(\uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIJ3HI_1_LC_15_10_4 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIJ3HI_1_LC_15_10_4 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIJ3HI_1_LC_15_10_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIJ3HI_1_LC_15_10_4  (
            .in0(N__9392),
            .in1(N__11296),
            .in2(N__9599),
            .in3(N__11314),
            .lcout(\uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7 ),
            .ltout(\uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_LC_15_10_5 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_LC_15_10_5 .LUT_INIT=16'b0000010001000100;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_LC_15_10_5  (
            .in0(N__16677),
            .in1(N__9535),
            .in2(N__9596),
            .in3(N__9588),
            .lcout(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ0Z_0_LC_15_10_6 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ0Z_0_LC_15_10_6 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ0Z_0_LC_15_10_6 .LUT_INIT=16'b1000101010101010;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ0Z_0_LC_15_10_6  (
            .in0(N__9536),
            .in1(N__9849),
            .in2(N__9527),
            .in3(N__9507),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16934),
            .ce(),
            .sr(N__13600));
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_5_LC_15_11_1 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_5_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_5_LC_15_11_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_5_LC_15_11_1  (
            .in0(_gnd_net_),
            .in1(N__16680),
            .in2(_gnd_net_),
            .in3(N__9682),
            .lcout(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_6_LC_15_11_2 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_6_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_6_LC_15_11_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_6_LC_15_11_2  (
            .in0(N__16681),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9655),
            .lcout(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_7_LC_15_11_3 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_7_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_7_LC_15_11_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_7_LC_15_11_3  (
            .in0(_gnd_net_),
            .in1(N__16682),
            .in2(_gnd_net_),
            .in3(N__9622),
            .lcout(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIGL56_8_LC_15_11_5 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIGL56_8_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIGL56_8_LC_15_11_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_RNIGL56_8_LC_15_11_5  (
            .in0(N__9416),
            .in1(N__9610),
            .in2(_gnd_net_),
            .in3(N__9404),
            .lcout(\uart_inst0.tx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_3_LC_15_11_6 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_3_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_3_LC_15_11_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_3_LC_15_11_6  (
            .in0(N__16679),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9724),
            .lcout(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_4_LC_15_12_0 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_4_LC_15_12_0 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_4_LC_15_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_4_LC_15_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9725),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16927),
            .ce(),
            .sr(N__13598));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_5_LC_15_12_1 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_5_LC_15_12_1 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_5_LC_15_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_5_LC_15_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15595),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16927),
            .ce(),
            .sr(N__13598));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_6_LC_15_12_2 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_6_LC_15_12_2 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_6_LC_15_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_6_LC_15_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9683),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16927),
            .ce(),
            .sr(N__13598));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_7_LC_15_12_3 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_7_LC_15_12_3 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_7_LC_15_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_7_LC_15_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9656),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16927),
            .ce(),
            .sr(N__13598));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_8_LC_15_12_5 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_8_LC_15_12_5 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_8_LC_15_12_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_8_LC_15_12_5  (
            .in0(_gnd_net_),
            .in1(N__9623),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rRamRdAddr_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16927),
            .ce(),
            .sr(N__13598));
    defparam \uart_inst0.uart_inst0.rx_countdown_4_LC_15_14_1 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_countdown_4_LC_15_14_1 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_countdown_4_LC_15_14_1 .LUT_INIT=16'b0010001000010001;
    LogicCell40 \uart_inst0.uart_inst0.rx_countdown_4_LC_15_14_1  (
            .in0(N__11333),
            .in1(N__11752),
            .in2(_gnd_net_),
            .in3(N__11762),
            .lcout(\uart_inst0.uart_inst0.rx_countdownZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16920),
            .ce(N__11710),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_countdown_2_LC_15_14_2 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_countdown_2_LC_15_14_2 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_countdown_2_LC_15_14_2 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \uart_inst0.uart_inst0.rx_countdown_2_LC_15_14_2  (
            .in0(N__11749),
            .in1(N__11363),
            .in2(N__14013),
            .in3(N__11693),
            .lcout(\uart_inst0.uart_inst0.rx_countdownZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16920),
            .ce(N__11710),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_countdown_3_LC_15_14_3 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_countdown_3_LC_15_14_3 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_countdown_3_LC_15_14_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \uart_inst0.uart_inst0.rx_countdown_3_LC_15_14_3  (
            .in0(N__11342),
            .in1(N__11275),
            .in2(N__14012),
            .in3(N__11750),
            .lcout(\uart_inst0.uart_inst0.rx_countdownZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16920),
            .ce(N__11710),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_countdown_1_LC_15_14_5 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_countdown_1_LC_15_14_5 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_countdown_1_LC_15_14_5 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \uart_inst0.uart_inst0.rx_countdown_1_LC_15_14_5  (
            .in0(N__11384),
            .in1(N__11151),
            .in2(N__14011),
            .in3(N__11748),
            .lcout(\uart_inst0.uart_inst0.rx_countdownZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16920),
            .ce(N__11710),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_countdown_0_LC_15_14_6 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_countdown_0_LC_15_14_6 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_countdown_0_LC_15_14_6 .LUT_INIT=16'b0100010000010001;
    LogicCell40 \uart_inst0.uart_inst0.rx_countdown_0_LC_15_14_6  (
            .in0(N__11751),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11432),
            .lcout(\uart_inst0.uart_inst0.rx_countdownZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16920),
            .ce(N__11710),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_state_RNO_2_0_LC_15_15_1 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_state_RNO_2_0_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_state_RNO_2_0_LC_15_15_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_inst0.uart_inst0.rx_state_RNO_2_0_LC_15_15_1  (
            .in0(N__11274),
            .in1(N__13780),
            .in2(N__13263),
            .in3(N__16034),
            .lcout(\uart_inst0.uart_inst0.rx_state_srsts_0_a5_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_state_RNI1VB3_5_LC_15_15_2 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_state_RNI1VB3_5_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_state_RNI1VB3_5_LC_15_15_2 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \uart_inst0.uart_inst0.rx_state_RNI1VB3_5_LC_15_15_2  (
            .in0(N__14014),
            .in1(N__11273),
            .in2(_gnd_net_),
            .in3(N__11128),
            .lcout(\uart_inst0.uart_inst0.rx_countdown_2_sqmuxa_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_countdown_RNIEE7V1_5_LC_15_15_3 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_countdown_RNIEE7V1_5_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_countdown_RNIEE7V1_5_LC_15_15_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_inst0.uart_inst0.rx_countdown_RNIEE7V1_5_LC_15_15_3  (
            .in0(N__11331),
            .in1(N__11353),
            .in2(N__11726),
            .in3(N__11374),
            .lcout(\uart_inst0.uart_inst0.rx_state_srsts_0_o2_3_3 ),
            .ltout(\uart_inst0.uart_inst0.rx_state_srsts_0_o2_3_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_countdown_RNIFVQU2_0_LC_15_15_4 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_countdown_RNIFVQU2_0_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_countdown_RNIFVQU2_0_LC_15_15_4 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \uart_inst0.uart_inst0.rx_countdown_RNIFVQU2_0_LC_15_15_4  (
            .in0(N__11430),
            .in1(_gnd_net_),
            .in2(N__9803),
            .in3(N__11404),
            .lcout(\uart_inst0.uart_inst0.N_257_0 ),
            .ltout(\uart_inst0.uart_inst0.N_257_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_state_RNIJD833_1_LC_15_15_5 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_state_RNIJD833_1_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_state_RNIJD833_1_LC_15_15_5 .LUT_INIT=16'b1110000011111111;
    LogicCell40 \uart_inst0.uart_inst0.rx_state_RNIJD833_1_LC_15_15_5  (
            .in0(N__13250),
            .in1(N__16033),
            .in2(N__9800),
            .in3(N__11455),
            .lcout(\uart_inst0.uart_inst0.N_252_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_RNIMJMP_3_LC_15_15_6 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_RNIMJMP_3_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_RNIMJMP_3_LC_15_15_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_inst0.uart_inst0.tx_bits_remaining_RNIMJMP_3_LC_15_15_6  (
            .in0(N__9796),
            .in1(N__9959),
            .in2(N__9773),
            .in3(N__9925),
            .lcout(\uart_inst0.uart_inst0.N_157 ),
            .ltout(\uart_inst0.uart_inst0.N_157_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_state_RNIR8D01_0_LC_15_15_7 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_state_RNIR8D01_0_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_state_RNIR8D01_0_LC_15_15_7 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \uart_inst0.uart_inst0.tx_state_RNIR8D01_0_LC_15_15_7  (
            .in0(_gnd_net_),
            .in1(N__11552),
            .in2(N__9740),
            .in3(N__11659),
            .lcout(\uart_inst0.uart_inst0.tx_state_1_sqmuxa_1_0_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_countdown_RNIEM2M1_0_2_LC_15_16_0 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_countdown_RNIEM2M1_0_2_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_countdown_RNIEM2M1_0_2_LC_15_16_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_inst0.uart_inst0.tx_countdown_RNIEM2M1_0_2_LC_15_16_0  (
            .in0(N__13630),
            .in1(N__14592),
            .in2(N__13684),
            .in3(N__14550),
            .lcout(\uart_inst0.uart_inst0.N_147_0 ),
            .ltout(\uart_inst0.uart_inst0.N_147_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_state_1_LC_15_16_1 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_state_1_LC_15_16_1 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.tx_state_1_LC_15_16_1 .LUT_INIT=16'b0010101010001000;
    LogicCell40 \uart_inst0.uart_inst0.tx_state_1_LC_15_16_1  (
            .in0(N__14004),
            .in1(N__11575),
            .in2(N__9890),
            .in3(N__11658),
            .lcout(\uart_inst0.uart_inst0.tx_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16911),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_state_RNO_0_1_LC_15_16_2 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_state_RNO_0_1_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_state_RNO_0_1_LC_15_16_2 .LUT_INIT=16'b0010001000110011;
    LogicCell40 \uart_inst0.uart_inst0.rx_state_RNO_0_1_LC_15_16_2  (
            .in0(N__13317),
            .in1(N__13254),
            .in2(_gnd_net_),
            .in3(N__11129),
            .lcout(),
            .ltout(\uart_inst0.uart_inst0.N_277_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_state_1_LC_15_16_3 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_state_1_LC_15_16_3 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_state_1_LC_15_16_3 .LUT_INIT=16'b0000100000001100;
    LogicCell40 \uart_inst0.uart_inst0.rx_state_1_LC_15_16_3  (
            .in0(N__11130),
            .in1(N__14023),
            .in2(N__9887),
            .in3(N__13823),
            .lcout(\uart_inst0.uart_inst0.rx_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16911),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_state_4_LC_15_16_4 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_state_4_LC_15_16_4 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_state_4_LC_15_16_4 .LUT_INIT=16'b1100010011000000;
    LogicCell40 \uart_inst0.uart_inst0.rx_state_4_LC_15_16_4  (
            .in0(N__13824),
            .in1(N__14003),
            .in2(N__11282),
            .in3(N__9875),
            .lcout(\uart_inst0.uart_inst0.rx_stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16911),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_state_RNO_1_0_LC_15_16_5 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_state_RNO_1_0_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_state_RNO_1_0_LC_15_16_5 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \uart_inst0.uart_inst0.rx_state_RNO_1_0_LC_15_16_5  (
            .in0(N__11691),
            .in1(N__9874),
            .in2(N__13787),
            .in3(N__13822),
            .lcout(),
            .ltout(\uart_inst0.uart_inst0.N_280_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_state_0_LC_15_16_6 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_state_0_LC_15_16_6 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_state_0_LC_15_16_6 .LUT_INIT=16'b1111010111111101;
    LogicCell40 \uart_inst0.uart_inst0.rx_state_0_LC_15_16_6  (
            .in0(N__14022),
            .in1(N__9884),
            .in2(N__9878),
            .in3(N__9860),
            .lcout(\uart_inst0.uart_inst0.rx_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16911),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_state_RNO_0_0_LC_15_16_7 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_state_RNO_0_0_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_state_RNO_0_0_LC_15_16_7 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \uart_inst0.uart_inst0.rx_state_RNO_0_0_LC_15_16_7  (
            .in0(N__11482),
            .in1(N__13316),
            .in2(_gnd_net_),
            .in3(N__9873),
            .lcout(\uart_inst0.uart_inst0.N_261_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_countdown_RNIEM2M1_2_LC_15_17_0 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_countdown_RNIEM2M1_2_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_countdown_RNIEM2M1_2_LC_15_17_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart_inst0.uart_inst0.tx_countdown_RNIEM2M1_2_LC_15_17_0  (
            .in0(N__13634),
            .in1(N__14590),
            .in2(N__13679),
            .in3(N__14543),
            .lcout(\uart_inst0.uart_inst0.N_147_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_state_RNO_0_0_LC_15_17_1 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_state_RNO_0_0_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_state_RNO_0_0_LC_15_17_1 .LUT_INIT=16'b1101111111011010;
    LogicCell40 \uart_inst0.uart_inst0.tx_state_RNO_0_0_LC_15_17_1  (
            .in0(N__11654),
            .in1(N__11858),
            .in2(N__11581),
            .in3(N__9854),
            .lcout(),
            .ltout(\uart_inst0.uart_inst0.tx_state_ns_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_state_0_LC_15_17_2 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_state_0_LC_15_17_2 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.tx_state_0_LC_15_17_2 .LUT_INIT=16'b1000110000001100;
    LogicCell40 \uart_inst0.uart_inst0.tx_state_0_LC_15_17_2  (
            .in0(N__11859),
            .in1(N__13999),
            .in2(N__9995),
            .in3(N__9992),
            .lcout(\uart_inst0.uart_inst0.tx_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16906),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_state_RNI1319_0_LC_15_17_3 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_state_RNI1319_0_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_state_RNI1319_0_LC_15_17_3 .LUT_INIT=16'b0101111100001111;
    LogicCell40 \uart_inst0.uart_inst0.tx_state_RNI1319_0_LC_15_17_3  (
            .in0(N__11560),
            .in1(_gnd_net_),
            .in2(N__14021),
            .in3(N__11651),
            .lcout(\uart_inst0.uart_inst0.tx_state_RNI1319Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_RNO_1_2_LC_15_17_4 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_RNO_1_2_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_RNO_1_2_LC_15_17_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uart_inst0.uart_inst0.tx_bits_remaining_RNO_1_2_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(N__9955),
            .in2(_gnd_net_),
            .in3(N__9926),
            .lcout(),
            .ltout(\uart_inst0.uart_inst0.un1_tx_bits_remaining_ac0_1_a0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_RNO_0_2_LC_15_17_5 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_RNO_0_2_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_bits_remaining_RNO_0_2_LC_15_17_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \uart_inst0.uart_inst0.tx_bits_remaining_RNO_0_2_LC_15_17_5  (
            .in0(N__11561),
            .in1(N__11857),
            .in2(N__9905),
            .in3(N__11652),
            .lcout(\uart_inst0.uart_inst0.un1_tx_bits_remaining_ac0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_countdown_RNIEGNA5_2_LC_15_17_6 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_countdown_RNIEGNA5_2_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_countdown_RNIEGNA5_2_LC_15_17_6 .LUT_INIT=16'b0111011100110011;
    LogicCell40 \uart_inst0.uart_inst0.tx_countdown_RNIEGNA5_2_LC_15_17_6  (
            .in0(N__11856),
            .in1(N__13998),
            .in2(_gnd_net_),
            .in3(N__10196),
            .lcout(\uart_inst0.uart_inst0.un1_rx_state49_i ),
            .ltout(\uart_inst0.uart_inst0.un1_rx_state49_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_clk_divider_esr_RNO_0_14_LC_15_17_7 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_esr_RNO_0_14_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_esr_RNO_0_14_LC_15_17_7 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \uart_inst0.uart_inst0.tx_clk_divider_esr_RNO_0_14_LC_15_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9896),
            .in3(N__13510),
            .lcout(\uart_inst0.uart_inst0.N_147_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_countdown_RNO_0_3_LC_15_18_0 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_countdown_RNO_0_3_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_countdown_RNO_0_3_LC_15_18_0 .LUT_INIT=16'b1011000011110000;
    LogicCell40 \uart_inst0.uart_inst0.tx_countdown_RNO_0_3_LC_15_18_0  (
            .in0(N__14547),
            .in1(N__11501),
            .in2(N__13680),
            .in3(N__10197),
            .lcout(),
            .ltout(\uart_inst0.uart_inst0.tx_countdown_RNO_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_countdown_3_LC_15_18_1 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_countdown_3_LC_15_18_1 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.tx_countdown_3_LC_15_18_1 .LUT_INIT=16'b1101100001110000;
    LogicCell40 \uart_inst0.uart_inst0.tx_countdown_3_LC_15_18_1  (
            .in0(N__11873),
            .in1(N__11587),
            .in2(N__9893),
            .in3(N__11665),
            .lcout(\uart_inst0.uart_inst0.tx_countdownZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16902),
            .ce(),
            .sr(N__13592));
    defparam \uart_inst0.uart_inst0.tx_clk_divider_esr_RNIIIJI_14_LC_15_18_2 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_esr_RNIIIJI_14_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_esr_RNIIIJI_14_LC_15_18_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \uart_inst0.uart_inst0.tx_clk_divider_esr_RNIIIJI_14_LC_15_18_2  (
            .in0(N__11955),
            .in1(N__11988),
            .in2(_gnd_net_),
            .in3(N__12115),
            .lcout(\uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_11_3 ),
            .ltout(\uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_11_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_clk_divider_esr_RNI4CAI3_14_LC_15_18_3 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_esr_RNI4CAI3_14_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_esr_RNI4CAI3_14_LC_15_18_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uart_inst0.uart_inst0.tx_clk_divider_esr_RNI4CAI3_14_LC_15_18_3  (
            .in0(N__14381),
            .in1(N__14470),
            .in2(N__10202),
            .in3(N__14500),
            .lcout(\uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_clk_divider_RNIQUQ11_4_LC_15_18_4 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_RNIQUQ11_4_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_RNIQUQ11_4_LC_15_18_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_inst0.uart_inst0.tx_clk_divider_RNIQUQ11_4_LC_15_18_4  (
            .in0(N__12045),
            .in1(N__12018),
            .in2(N__12077),
            .in3(N__11787),
            .lcout(\uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_clk_divider_RNIEC1S_10_LC_15_19_0 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_RNIEC1S_10_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_RNIEC1S_10_LC_15_19_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_inst0.uart_inst0.tx_clk_divider_RNIEC1S_10_LC_15_19_0  (
            .in0(N__12502),
            .in1(N__11901),
            .in2(N__12148),
            .in3(N__11925),
            .lcout(\uart_inst0.uart_inst0.tx_countdown_0_sqmuxa_1_13_11_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_clk_divider_10_LC_15_19_1 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_10_LC_15_19_1 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_10_LC_15_19_1 .LUT_INIT=16'b1010101001100110;
    LogicCell40 \uart_inst0.uart_inst0.tx_clk_divider_10_LC_15_19_1  (
            .in0(N__11926),
            .in1(N__13549),
            .in2(_gnd_net_),
            .in3(N__11912),
            .lcout(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16899),
            .ce(),
            .sr(N__14636));
    defparam \uart_inst0.uart_inst0.tx_clk_divider_11_LC_15_19_2 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_11_LC_15_19_2 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_11_LC_15_19_2 .LUT_INIT=16'b1101110100100010;
    LogicCell40 \uart_inst0.uart_inst0.tx_clk_divider_11_LC_15_19_2  (
            .in0(N__13550),
            .in1(N__11888),
            .in2(_gnd_net_),
            .in3(N__11902),
            .lcout(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16899),
            .ce(),
            .sr(N__14636));
    defparam \uart_inst0.uart_inst0.tx_clk_divider_13_LC_15_19_4 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_13_LC_15_19_4 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_13_LC_15_19_4 .LUT_INIT=16'b1010101001011010;
    LogicCell40 \uart_inst0.uart_inst0.tx_clk_divider_13_LC_15_19_4  (
            .in0(N__12144),
            .in1(_gnd_net_),
            .in2(N__13556),
            .in3(N__12128),
            .lcout(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16899),
            .ce(),
            .sr(N__14636));
    defparam \uart_inst0.uart_inst0.tx_clk_divider_5_LC_15_19_6 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_5_LC_15_19_6 .SEQ_MODE=4'b1001;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_5_LC_15_19_6 .LUT_INIT=16'b1101110100100010;
    LogicCell40 \uart_inst0.uart_inst0.tx_clk_divider_5_LC_15_19_6  (
            .in0(N__13554),
            .in1(N__12056),
            .in2(_gnd_net_),
            .in3(N__12076),
            .lcout(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16899),
            .ce(),
            .sr(N__14636));
    defparam \uart_inst0.uart_inst0.tx_clk_divider_6_LC_15_19_7 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_6_LC_15_19_7 .SEQ_MODE=4'b1001;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_6_LC_15_19_7 .LUT_INIT=16'b1101110100100010;
    LogicCell40 \uart_inst0.uart_inst0.tx_clk_divider_6_LC_15_19_7  (
            .in0(N__13555),
            .in1(N__12029),
            .in2(_gnd_net_),
            .in3(N__12047),
            .lcout(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16899),
            .ce(),
            .sr(N__14636));
    defparam rTxData_0_LC_16_1_5.C_ON=1'b0;
    defparam rTxData_0_LC_16_1_5.SEQ_MODE=4'b1000;
    defparam rTxData_0_LC_16_1_5.LUT_INIT=16'b1100110011101110;
    LogicCell40 rTxData_0_LC_16_1_5 (
            .in0(N__14020),
            .in1(N__10102),
            .in2(_gnd_net_),
            .in3(N__10173),
            .lcout(rTxDataZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16981),
            .ce(),
            .sr(N__16357));
    defparam \fifo_inst.ft2232h_inst.rTxBusReady_esr_LC_16_2_7 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rTxBusReady_esr_LC_16_2_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rTxBusReady_esr_LC_16_2_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \fifo_inst.ft2232h_inst.rTxBusReady_esr_LC_16_2_7  (
            .in0(N__10607),
            .in1(N__10652),
            .in2(_gnd_net_),
            .in3(N__10532),
            .lcout(rTxBusReady),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16978),
            .ce(N__10469),
            .sr(N__16359));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_3_LC_16_3_0 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_3_LC_16_3_0 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_3_LC_16_3_0 .LUT_INIT=16'b0001000010110000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_3_LC_16_3_0  (
            .in0(N__10226),
            .in1(N__16645),
            .in2(N__10445),
            .in3(N__10280),
            .lcout(fifo_inst_tx_fifo_inst_rRamRdAddr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16976),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m74_LC_16_3_1 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m74_LC_16_3_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m74_LC_16_3_1 .LUT_INIT=16'b0100011100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m74_LC_16_3_1  (
            .in0(N__10278),
            .in1(N__10224),
            .in2(N__16698),
            .in3(N__10441),
            .lcout(m74),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m72_e_5_LC_16_3_2 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m72_e_5_LC_16_3_2 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m72_e_5_LC_16_3_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m72_e_5_LC_16_3_2  (
            .in0(N__10417),
            .in1(N__10291),
            .in2(N__16697),
            .in3(N__12775),
            .lcout(),
            .ltout(\uart_inst0.tx_uart_fifo_inst.m72_eZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m72_e_LC_16_3_3 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m72_e_LC_16_3_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m72_e_LC_16_3_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m72_e_LC_16_3_3  (
            .in0(N__10405),
            .in1(N__10394),
            .in2(N__10382),
            .in3(N__10319),
            .lcout(\uart_inst0.tx_uart_fifo_inst.N_100 ),
            .ltout(\uart_inst0.tx_uart_fifo_inst.N_100_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m73_LC_16_3_4 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m73_LC_16_3_4 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m73_LC_16_3_4 .LUT_INIT=16'b0000010011000100;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m73_LC_16_3_4  (
            .in0(N__16644),
            .in1(N__10234),
            .in2(N__10379),
            .in3(N__10277),
            .lcout(m73),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m72_e_6_LC_16_3_5 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m72_e_6_LC_16_3_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m72_e_6_LC_16_3_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m72_e_6_LC_16_3_5  (
            .in0(N__10360),
            .in1(N__10348),
            .in2(N__10337),
            .in3(N__10213),
            .lcout(\uart_inst0.tx_uart_fifo_inst.m72_eZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_4_LC_16_3_6 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_4_LC_16_3_6 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_4_LC_16_3_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_4_LC_16_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10303),
            .lcout(fifo_inst_tx_fifo_inst_rRamRdAddr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16976),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_0_LC_16_3_7 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_0_LC_16_3_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_0_LC_16_3_7 .LUT_INIT=16'b0101000000110000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_0_LC_16_3_7  (
            .in0(N__10279),
            .in1(N__16640),
            .in2(N__10238),
            .in3(N__10225),
            .lcout(fifo_inst_tx_fifo_inst_rRamRdAddr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16976),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_7_LC_16_4_0 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_7_LC_16_4_0 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_7_LC_16_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.rx_fifo_inst.rRamRdAddr_7_LC_16_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10792),
            .lcout(fifo_inst_rx_fifo_inst_rRamRdAddr_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16973),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_3_LC_16_4_2 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_3_LC_16_4_2 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_3_LC_16_4_2 .LUT_INIT=16'b0000010010001100;
    LogicCell40 \fifo_inst.rx_fifo_inst.rRamRdAddr_3_LC_16_4_2  (
            .in0(N__10994),
            .in1(N__10757),
            .in2(N__16699),
            .in3(N__10966),
            .lcout(fifo_inst_rx_fifo_inst_rRamRdAddr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16973),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_1_LC_16_4_3 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_1_LC_16_4_3 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_1_LC_16_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.rx_fifo_inst.rRamRdAddr_1_LC_16_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10768),
            .lcout(fifo_inst_rx_fifo_inst_rRamRdAddr_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16973),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m60_LC_16_4_4 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m60_LC_16_4_4 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m60_LC_16_4_4 .LUT_INIT=16'b0001110100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m60_LC_16_4_4  (
            .in0(N__16653),
            .in1(N__10993),
            .in2(N__10967),
            .in3(N__10756),
            .lcout(m60),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_4_LC_16_5_0 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_4_LC_16_5_0 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_4_LC_16_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.rx_fifo_inst.rRamRdAddr_4_LC_16_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10723),
            .lcout(fifo_inst_rx_fifo_inst_rRamRdAddr_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16969),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m58_e_6_LC_16_5_1 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m58_e_6_LC_16_5_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m58_e_6_LC_16_5_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m58_e_6_LC_16_5_1  (
            .in0(N__10711),
            .in1(N__10699),
            .in2(N__10688),
            .in3(N__10912),
            .lcout(\uart_inst0.tx_uart_fifo_inst.m58_eZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rFifoState_1_sqmuxa_0_i_LC_16_5_2 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rFifoState_1_sqmuxa_0_i_LC_16_5_2 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.un1_rFifoState_1_sqmuxa_0_i_LC_16_5_2 .LUT_INIT=16'b1010101010101110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.un1_rFifoState_1_sqmuxa_0_i_LC_16_5_2  (
            .in0(N__10673),
            .in1(N__10657),
            .in2(N__10593),
            .in3(N__10531),
            .lcout(),
            .ltout(fifo_inst_ft2232h_inst_un1_rFifoState_1_sqmuxa_0_i_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ft2232h_inst.rTxBusReady_esr_RNO_LC_16_5_3 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rTxBusReady_esr_RNO_LC_16_5_3 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.ft2232h_inst.rTxBusReady_esr_RNO_LC_16_5_3 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \fifo_inst.ft2232h_inst.rTxBusReady_esr_RNO_LC_16_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10472),
            .in3(N__14100),
            .lcout(\fifo_inst.ft2232h_inst.un1_rFifoState_1_sqmuxa_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m59_LC_16_5_4 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m59_LC_16_5_4 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m59_LC_16_5_4 .LUT_INIT=16'b0000010010001100;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m59_LC_16_5_4  (
            .in0(N__10992),
            .in1(N__10975),
            .in2(N__16701),
            .in3(N__10961),
            .lcout(m59),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m58_e_5_LC_16_5_5 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m58_e_5_LC_16_5_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m58_e_5_LC_16_5_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m58_e_5_LC_16_5_5  (
            .in0(N__11078),
            .in1(N__11062),
            .in2(N__16702),
            .in3(N__11051),
            .lcout(),
            .ltout(\uart_inst0.tx_uart_fifo_inst.m58_eZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m58_e_LC_16_5_6 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m58_e_LC_16_5_6 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m58_e_LC_16_5_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m58_e_LC_16_5_6  (
            .in0(N__11033),
            .in1(N__11017),
            .in2(N__11003),
            .in3(N__11000),
            .lcout(\uart_inst0.tx_uart_fifo_inst.N_99 ),
            .ltout(\uart_inst0.tx_uart_fifo_inst.N_99_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_0_LC_16_5_7 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_0_LC_16_5_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rRamRdAddr_0_LC_16_5_7 .LUT_INIT=16'b0010000000101010;
    LogicCell40 \fifo_inst.rx_fifo_inst.rRamRdAddr_0_LC_16_5_7  (
            .in0(N__10976),
            .in1(N__10962),
            .in2(N__10916),
            .in3(N__16666),
            .lcout(fifo_inst_rx_fifo_inst_rRamRdAddr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16969),
            .ce(),
            .sr(_gnd_net_));
    defparam rRxData_4_LC_16_6_0.C_ON=1'b0;
    defparam rRxData_4_LC_16_6_0.SEQ_MODE=4'b1000;
    defparam rRxData_4_LC_16_6_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 rRxData_4_LC_16_6_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14774),
            .lcout(rRxDataZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16961),
            .ce(N__12850),
            .sr(_gnd_net_));
    defparam rUartTxData_esr_3_LC_16_7_3.C_ON=1'b0;
    defparam rUartTxData_esr_3_LC_16_7_3.SEQ_MODE=4'b1000;
    defparam rUartTxData_esr_3_LC_16_7_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 rUartTxData_esr_3_LC_16_7_3 (
            .in0(N__10901),
            .in1(N__12512),
            .in2(_gnd_net_),
            .in3(N__11244),
            .lcout(rUartTxDataZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16955),
            .ce(N__11183),
            .sr(N__16418));
    defparam rUartTxData_esr_4_LC_16_7_4.C_ON=1'b0;
    defparam rUartTxData_esr_4_LC_16_7_4.SEQ_MODE=4'b1000;
    defparam rUartTxData_esr_4_LC_16_7_4.LUT_INIT=16'b1111010110100000;
    LogicCell40 rUartTxData_esr_4_LC_16_7_4 (
            .in0(N__11245),
            .in1(_gnd_net_),
            .in2(N__10877),
            .in3(N__10865),
            .lcout(rUartTxDataZ0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16955),
            .ce(N__11183),
            .sr(N__16418));
    defparam rUartTxData_esr_7_LC_16_7_5.C_ON=1'b0;
    defparam rUartTxData_esr_7_LC_16_7_5.SEQ_MODE=4'b1000;
    defparam rUartTxData_esr_7_LC_16_7_5.LUT_INIT=16'b1111000010101010;
    LogicCell40 rUartTxData_esr_7_LC_16_7_5 (
            .in0(N__12860),
            .in1(_gnd_net_),
            .in2(N__10847),
            .in3(N__11246),
            .lcout(rUartTxDataZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16955),
            .ce(N__11183),
            .sr(N__16418));
    defparam rUartTxData_esr_2_LC_16_7_6.C_ON=1'b0;
    defparam rUartTxData_esr_2_LC_16_7_6.SEQ_MODE=4'b1000;
    defparam rUartTxData_esr_2_LC_16_7_6.LUT_INIT=16'b1111101001010000;
    LogicCell40 rUartTxData_esr_2_LC_16_7_6 (
            .in0(N__11243),
            .in1(_gnd_net_),
            .in2(N__12524),
            .in3(N__10826),
            .lcout(rUartTxDataZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16955),
            .ce(N__11183),
            .sr(N__16418));
    defparam rUartTxData_esr_0_LC_16_7_7.C_ON=1'b0;
    defparam rUartTxData_esr_0_LC_16_7_7.SEQ_MODE=4'b1000;
    defparam rUartTxData_esr_0_LC_16_7_7.LUT_INIT=16'b1100110010101010;
    LogicCell40 rUartTxData_esr_0_LC_16_7_7 (
            .in0(N__12881),
            .in1(N__11255),
            .in2(_gnd_net_),
            .in3(N__11242),
            .lcout(rUartTxDataZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16955),
            .ce(N__11183),
            .sr(N__16418));
    defparam rUartRxState_RNITBQ5_0_LC_16_8_3.C_ON=1'b0;
    defparam rUartRxState_RNITBQ5_0_LC_16_8_3.SEQ_MODE=4'b0000;
    defparam rUartRxState_RNITBQ5_0_LC_16_8_3.LUT_INIT=16'b1111111111001100;
    LogicCell40 rUartRxState_RNITBQ5_0_LC_16_8_3 (
            .in0(_gnd_net_),
            .in1(N__16675),
            .in2(_gnd_net_),
            .in3(N__13040),
            .lcout(rUartRxState_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNO_0_1_LC_16_8_6 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNO_0_1_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNO_0_1_LC_16_8_6 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rDataCount_RNO_0_1_LC_16_8_6  (
            .in0(N__13140),
            .in1(N__13093),
            .in2(_gnd_net_),
            .in3(N__14949),
            .lcout(\uart_inst0.rx_uart_fifo_inst.un1_rDataCount15_2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNIG8UP_3_LC_16_9_2 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNIG8UP_3_LC_16_9_2 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNIG8UP_3_LC_16_9_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rDataCount_RNIG8UP_3_LC_16_9_2  (
            .in0(_gnd_net_),
            .in1(N__11103),
            .in2(_gnd_net_),
            .in3(N__12929),
            .lcout(\uart_inst0.rx_uart_fifo_inst.wRamWrEn ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rRxWrEn_LC_16_9_3 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rRxWrEn_LC_16_9_3 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rRxWrEn_LC_16_9_3 .LUT_INIT=16'b1100010011110100;
    LogicCell40 \uart_inst0.uart_inst0.rRxWrEn_LC_16_9_3  (
            .in0(N__12930),
            .in1(N__11483),
            .in2(N__11108),
            .in3(N__11156),
            .lcout(\uart_inst0.wRxWrEn_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16944),
            .ce(),
            .sr(N__16425));
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNO_0_3_LC_16_9_4 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNO_0_3_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNO_0_3_LC_16_9_4 .LUT_INIT=16'b0001011100011111;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rDataCount_RNO_0_3_LC_16_9_4  (
            .in0(N__13002),
            .in1(N__13094),
            .in2(N__14962),
            .in3(N__11104),
            .lcout(\uart_inst0.rx_uart_fifo_inst.un1_rDataCount_axbxc3_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_0_LC_16_10_7 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_0_LC_16_10_7 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_0_LC_16_10_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_0_LC_16_10_7  (
            .in0(_gnd_net_),
            .in1(N__16678),
            .in2(_gnd_net_),
            .in3(N__13216),
            .lcout(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_1_LC_16_11_0 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_1_LC_16_11_0 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_1_LC_16_11_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_1_LC_16_11_0  (
            .in0(_gnd_net_),
            .in1(N__13217),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16935),
            .ce(),
            .sr(N__13601));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_2_LC_16_11_1 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_2_LC_16_11_1 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_2_LC_16_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_2_LC_16_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15710),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16935),
            .ce(),
            .sr(N__13601));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_4_LC_16_11_2 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_4_LC_16_11_2 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_4_LC_16_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_4_LC_16_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15491),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16935),
            .ce(),
            .sr(N__13601));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_5_LC_16_11_3 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_5_LC_16_11_3 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_5_LC_16_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_5_LC_16_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15446),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16935),
            .ce(),
            .sr(N__13601));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_6_LC_16_11_4 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_6_LC_16_11_4 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_6_LC_16_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_6_LC_16_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15512),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16935),
            .ce(),
            .sr(N__13601));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_7_LC_16_11_5 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_7_LC_16_11_5 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_7_LC_16_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_7_LC_16_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15731),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16935),
            .ce(),
            .sr(N__13601));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ0Z_1_LC_16_11_6 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ0Z_1_LC_16_11_6 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ0Z_1_LC_16_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ0Z_1_LC_16_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13484),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16935),
            .ce(),
            .sr(N__13601));
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_2_LC_16_11_7 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_2_LC_16_11_7 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_2_LC_16_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.rRamRdAddr_2_LC_16_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15623),
            .lcout(\uart_inst0.tx_uart_fifo_inst.rRamRdAddrZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16935),
            .ce(),
            .sr(N__13601));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_8_LC_16_12_1 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_8_LC_16_12_1 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_8_LC_16_12_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_8_LC_16_12_1  (
            .in0(_gnd_net_),
            .in1(N__15689),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16931),
            .ce(),
            .sr(N__13599));
    defparam \uart_inst0.uart_inst0.rRxData_7_LC_16_13_1 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rRxData_7_LC_16_13_1 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rRxData_7_LC_16_13_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uart_inst0.uart_inst0.rRxData_7_LC_16_13_1  (
            .in0(N__13290),
            .in1(N__16137),
            .in2(_gnd_net_),
            .in3(N__14036),
            .lcout(\uart_inst0.wRxWrData_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16928),
            .ce(),
            .sr(N__16449));
    defparam \uart_inst0.uart_inst0.rx_state_5_LC_16_14_0 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_state_5_LC_16_14_0 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_state_5_LC_16_14_0 .LUT_INIT=16'b1100101000000000;
    LogicCell40 \uart_inst0.uart_inst0.rx_state_5_LC_16_14_0  (
            .in0(N__13779),
            .in1(N__13259),
            .in2(N__13319),
            .in3(N__15937),
            .lcout(\uart_inst0.uart_inst0.rx_stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16925),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_countdown_RNIBD513_0_LC_16_14_3 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_countdown_RNIBD513_0_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_countdown_RNIBD513_0_LC_16_14_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \uart_inst0.uart_inst0.rx_countdown_RNIBD513_0_LC_16_14_3  (
            .in0(N__11402),
            .in1(N__11428),
            .in2(N__13986),
            .in3(N__11464),
            .lcout(\uart_inst0.uart_inst0.N_283 ),
            .ltout(\uart_inst0.uart_inst0.N_283_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_state_6_LC_16_14_4 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_state_6_LC_16_14_4 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_state_6_LC_16_14_4 .LUT_INIT=16'b1000000010000000;
    LogicCell40 \uart_inst0.uart_inst0.rx_state_6_LC_16_14_4  (
            .in0(N__13315),
            .in1(N__13778),
            .in2(N__11486),
            .in3(_gnd_net_),
            .lcout(\uart_inst0.uart_inst0.rx_stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16925),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_countdown_RNIHNBV2_0_LC_16_14_5 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_countdown_RNIHNBV2_0_LC_16_14_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_countdown_RNIHNBV2_0_LC_16_14_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \uart_inst0.uart_inst0.rx_countdown_RNIHNBV2_0_LC_16_14_5  (
            .in0(N__11403),
            .in1(N__11429),
            .in2(N__16044),
            .in3(N__11465),
            .lcout(\uart_inst0.uart_inst0.rRxData_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_state_RNI3F11_1_LC_16_14_6 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_state_RNI3F11_1_LC_16_14_6 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_state_RNI3F11_1_LC_16_14_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uart_inst0.uart_inst0.rx_state_RNI3F11_1_LC_16_14_6  (
            .in0(_gnd_net_),
            .in1(N__16032),
            .in2(_gnd_net_),
            .in3(N__13258),
            .lcout(\uart_inst0.uart_inst0.N_258_0 ),
            .ltout(\uart_inst0.uart_inst0.N_258_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_state_RNIGVTK5_5_LC_16_14_7 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_state_RNIGVTK5_5_LC_16_14_7 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_state_RNIGVTK5_5_LC_16_14_7 .LUT_INIT=16'b1101111111011101;
    LogicCell40 \uart_inst0.uart_inst0.rx_state_RNIGVTK5_5_LC_16_14_7  (
            .in0(N__11456),
            .in1(N__11444),
            .in2(N__11435),
            .in3(N__13825),
            .lcout(\uart_inst0.uart_inst0.rx_countdowne_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_countdown_cry_c_0_LC_16_15_0 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.rx_countdown_cry_c_0_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_countdown_cry_c_0_LC_16_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \uart_inst0.uart_inst0.rx_countdown_cry_c_0_LC_16_15_0  (
            .in0(_gnd_net_),
            .in1(N__11431),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_16_15_0_),
            .carryout(\uart_inst0.uart_inst0.rx_countdown_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_countdown_RNO_0_1_LC_16_15_1 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.rx_countdown_RNO_0_1_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_countdown_RNO_0_1_LC_16_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_inst0.uart_inst0.rx_countdown_RNO_0_1_LC_16_15_1  (
            .in0(_gnd_net_),
            .in1(N__11405),
            .in2(N__12405),
            .in3(N__11378),
            .lcout(\uart_inst0.uart_inst0.rx_countdown_s_1 ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.rx_countdown_cry_0 ),
            .carryout(\uart_inst0.uart_inst0.rx_countdown_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_countdown_RNO_0_2_LC_16_15_2 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.rx_countdown_RNO_0_2_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_countdown_RNO_0_2_LC_16_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_inst0.uart_inst0.rx_countdown_RNO_0_2_LC_16_15_2  (
            .in0(_gnd_net_),
            .in1(N__11375),
            .in2(N__12407),
            .in3(N__11357),
            .lcout(\uart_inst0.uart_inst0.rx_countdown_s_2 ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.rx_countdown_cry_1 ),
            .carryout(\uart_inst0.uart_inst0.rx_countdown_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_countdown_RNO_0_3_LC_16_15_3 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.rx_countdown_RNO_0_3_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_countdown_RNO_0_3_LC_16_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uart_inst0.uart_inst0.rx_countdown_RNO_0_3_LC_16_15_3  (
            .in0(_gnd_net_),
            .in1(N__11354),
            .in2(N__12406),
            .in3(N__11336),
            .lcout(\uart_inst0.uart_inst0.rx_countdown_s_3 ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.rx_countdown_cry_2 ),
            .carryout(\uart_inst0.uart_inst0.rx_countdown_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_countdown_cry_3_THRU_LUT4_0_LC_16_15_4 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.rx_countdown_cry_3_THRU_LUT4_0_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_countdown_cry_3_THRU_LUT4_0_LC_16_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.uart_inst0.rx_countdown_cry_3_THRU_LUT4_0_LC_16_15_4  (
            .in0(_gnd_net_),
            .in1(N__11332),
            .in2(N__12408),
            .in3(N__11756),
            .lcout(\uart_inst0.uart_inst0.rx_countdown_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.rx_countdown_cry_3 ),
            .carryout(\uart_inst0.uart_inst0.rx_countdown_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_countdown_5_LC_16_15_5 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_countdown_5_LC_16_15_5 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_countdown_5_LC_16_15_5 .LUT_INIT=16'b0100010000010001;
    LogicCell40 \uart_inst0.uart_inst0.rx_countdown_5_LC_16_15_5  (
            .in0(N__11753),
            .in1(N__11725),
            .in2(_gnd_net_),
            .in3(N__11729),
            .lcout(\uart_inst0.uart_inst0.rx_countdownZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16921),
            .ce(N__11711),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_state_RNO_1_2_LC_16_16_1 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_state_RNO_1_2_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_state_RNO_1_2_LC_16_16_1 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \uart_inst0.uart_inst0.rx_state_RNO_1_2_LC_16_16_1  (
            .in0(N__13724),
            .in1(N__13739),
            .in2(N__13264),
            .in3(N__13818),
            .lcout(),
            .ltout(\uart_inst0.uart_inst0.N_276_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_state_2_LC_16_16_2 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_state_2_LC_16_16_2 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_state_2_LC_16_16_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uart_inst0.uart_inst0.rx_state_2_LC_16_16_2  (
            .in0(N__14005),
            .in1(N__11692),
            .in2(N__11672),
            .in3(N__11492),
            .lcout(\uart_inst0.uart_inst0.rx_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16915),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_countdown_RNO_0_2_LC_16_16_4 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_countdown_RNO_0_2_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_countdown_RNO_0_2_LC_16_16_4 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \uart_inst0.uart_inst0.tx_countdown_RNO_0_2_LC_16_16_4  (
            .in0(N__14600),
            .in1(N__11653),
            .in2(N__11583),
            .in3(N__14555),
            .lcout(\uart_inst0.uart_inst0.tx_N_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_countdown_RNO_1_3_LC_16_16_5 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_countdown_RNO_1_3_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_countdown_RNO_1_3_LC_16_16_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \uart_inst0.uart_inst0.tx_countdown_RNO_1_3_LC_16_16_5  (
            .in0(N__13628),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14599),
            .lcout(\uart_inst0.uart_inst0.un1_m3_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_state_RNO_0_2_LC_16_16_7 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_state_RNO_0_2_LC_16_16_7 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_state_RNO_0_2_LC_16_16_7 .LUT_INIT=16'b0010001000110011;
    LogicCell40 \uart_inst0.uart_inst0.rx_state_RNO_0_2_LC_16_16_7  (
            .in0(N__13318),
            .in1(N__16022),
            .in2(_gnd_net_),
            .in3(N__13817),
            .lcout(\uart_inst0.uart_inst0.N_275 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_clk_divider_7_LC_16_17_0 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_7_LC_16_17_0 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_7_LC_16_17_0 .LUT_INIT=16'b1001100110101010;
    LogicCell40 \uart_inst0.uart_inst0.tx_clk_divider_7_LC_16_17_0  (
            .in0(N__12020),
            .in1(N__12002),
            .in2(_gnd_net_),
            .in3(N__13545),
            .lcout(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16912),
            .ce(),
            .sr(N__14635));
    defparam \uart_inst0.uart_inst0.tx_clk_divider_8_LC_16_17_1 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_8_LC_16_17_1 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_8_LC_16_17_1 .LUT_INIT=16'b1101110100100010;
    LogicCell40 \uart_inst0.uart_inst0.tx_clk_divider_8_LC_16_17_1  (
            .in0(N__13546),
            .in1(N__11972),
            .in2(_gnd_net_),
            .in3(N__11992),
            .lcout(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16912),
            .ce(),
            .sr(N__14635));
    defparam \uart_inst0.uart_inst0.tx_clk_divider_9_LC_16_17_2 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_9_LC_16_17_2 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_9_LC_16_17_2 .LUT_INIT=16'b1001100110101010;
    LogicCell40 \uart_inst0.uart_inst0.tx_clk_divider_9_LC_16_17_2  (
            .in0(N__11959),
            .in1(N__11939),
            .in2(_gnd_net_),
            .in3(N__13547),
            .lcout(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16912),
            .ce(),
            .sr(N__14635));
    defparam \uart_inst0.uart_inst0.tx_clk_divider_12_LC_16_17_3 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_12_LC_16_17_3 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_12_LC_16_17_3 .LUT_INIT=16'b1101110100100010;
    LogicCell40 \uart_inst0.uart_inst0.tx_clk_divider_12_LC_16_17_3  (
            .in0(N__13541),
            .in1(N__12482),
            .in2(_gnd_net_),
            .in3(N__12501),
            .lcout(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16912),
            .ce(),
            .sr(N__14635));
    defparam \uart_inst0.uart_inst0.tx_clk_divider_4_LC_16_17_4 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_4_LC_16_17_4 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_4_LC_16_17_4 .LUT_INIT=16'b1011101101000100;
    LogicCell40 \uart_inst0.uart_inst0.tx_clk_divider_4_LC_16_17_4  (
            .in0(N__11771),
            .in1(N__13544),
            .in2(_gnd_net_),
            .in3(N__11789),
            .lcout(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16912),
            .ce(),
            .sr(N__14635));
    defparam \uart_inst0.uart_inst0.tx_clk_divider_1_LC_16_17_5 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_1_LC_16_17_5 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_1_LC_16_17_5 .LUT_INIT=16'b1111010100001010;
    LogicCell40 \uart_inst0.uart_inst0.tx_clk_divider_1_LC_16_17_5  (
            .in0(N__13542),
            .in1(_gnd_net_),
            .in2(N__11813),
            .in3(N__14399),
            .lcout(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16912),
            .ce(),
            .sr(N__14635));
    defparam \uart_inst0.uart_inst0.tx_clk_divider_2_LC_16_17_7 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_2_LC_16_17_7 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_2_LC_16_17_7 .LUT_INIT=16'b1101110100100010;
    LogicCell40 \uart_inst0.uart_inst0.tx_clk_divider_2_LC_16_17_7  (
            .in0(N__13543),
            .in1(N__11801),
            .in2(_gnd_net_),
            .in3(N__14450),
            .lcout(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16912),
            .ce(),
            .sr(N__14635));
    defparam \uart_inst0.uart_inst0.tx_clk_divider_0_LC_16_18_0 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_0_LC_16_18_0 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_0_LC_16_18_0 .LUT_INIT=16'b1001100110011001;
    LogicCell40 \uart_inst0.uart_inst0.tx_clk_divider_0_LC_16_18_0  (
            .in0(N__11874),
            .in1(N__14432),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_0 ),
            .ltout(),
            .carryin(bfn_16_18_0_),
            .carryout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_0_s1 ),
            .clk(N__16907),
            .ce(),
            .sr(N__14642));
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_0_s1_THRU_LUT4_0_LC_16_18_1 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_0_s1_THRU_LUT4_0_LC_16_18_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_0_s1_THRU_LUT4_0_LC_16_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_0_s1_THRU_LUT4_0_LC_16_18_1  (
            .in0(_gnd_net_),
            .in1(N__14398),
            .in2(N__12449),
            .in3(N__11804),
            .lcout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_0_s1_THRU_CO ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_0_s1 ),
            .carryout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_1_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_1_s1_THRU_LUT4_0_LC_16_18_2 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_1_s1_THRU_LUT4_0_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_1_s1_THRU_LUT4_0_LC_16_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_1_s1_THRU_LUT4_0_LC_16_18_2  (
            .in0(_gnd_net_),
            .in1(N__14449),
            .in2(N__12453),
            .in3(N__11795),
            .lcout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_1_s1_THRU_CO ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_1_s1 ),
            .carryout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_2_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_2_s1_THRU_LUT4_0_LC_16_18_3 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_2_s1_THRU_LUT4_0_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_2_s1_THRU_LUT4_0_LC_16_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_2_s1_THRU_LUT4_0_LC_16_18_3  (
            .in0(_gnd_net_),
            .in1(N__14418),
            .in2(N__12450),
            .in3(N__11792),
            .lcout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_2_s1_THRU_CO ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_2_s1 ),
            .carryout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_3_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_3_s1_THRU_LUT4_0_LC_16_18_4 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_3_s1_THRU_LUT4_0_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_3_s1_THRU_LUT4_0_LC_16_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_3_s1_THRU_LUT4_0_LC_16_18_4  (
            .in0(_gnd_net_),
            .in1(N__11788),
            .in2(N__12454),
            .in3(N__11765),
            .lcout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_3_s1_THRU_CO ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_3_s1 ),
            .carryout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_4_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_4_s1_THRU_LUT4_0_LC_16_18_5 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_4_s1_THRU_LUT4_0_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_4_s1_THRU_LUT4_0_LC_16_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_4_s1_THRU_LUT4_0_LC_16_18_5  (
            .in0(_gnd_net_),
            .in1(N__12075),
            .in2(N__12451),
            .in3(N__12050),
            .lcout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_4_s1_THRU_CO ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_4_s1 ),
            .carryout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_5_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_5_s1_THRU_LUT4_0_LC_16_18_6 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_5_s1_THRU_LUT4_0_LC_16_18_6 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_5_s1_THRU_LUT4_0_LC_16_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_5_s1_THRU_LUT4_0_LC_16_18_6  (
            .in0(_gnd_net_),
            .in1(N__12046),
            .in2(N__12455),
            .in3(N__12023),
            .lcout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_5_s1_THRU_CO ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_5_s1 ),
            .carryout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_6_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_6_s1_THRU_LUT4_0_LC_16_18_7 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_6_s1_THRU_LUT4_0_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_6_s1_THRU_LUT4_0_LC_16_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_6_s1_THRU_LUT4_0_LC_16_18_7  (
            .in0(_gnd_net_),
            .in1(N__12019),
            .in2(N__12452),
            .in3(N__11996),
            .lcout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_6_s1_THRU_CO ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_6_s1 ),
            .carryout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_7_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_7_s1_THRU_LUT4_0_LC_16_19_0 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_7_s1_THRU_LUT4_0_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_7_s1_THRU_LUT4_0_LC_16_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_7_s1_THRU_LUT4_0_LC_16_19_0  (
            .in0(_gnd_net_),
            .in1(N__11993),
            .in2(N__12459),
            .in3(N__11963),
            .lcout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_7_s1_THRU_CO ),
            .ltout(),
            .carryin(bfn_16_19_0_),
            .carryout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_8_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_8_s1_THRU_LUT4_0_LC_16_19_1 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_8_s1_THRU_LUT4_0_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_8_s1_THRU_LUT4_0_LC_16_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_8_s1_THRU_LUT4_0_LC_16_19_1  (
            .in0(_gnd_net_),
            .in1(N__11960),
            .in2(N__12457),
            .in3(N__11930),
            .lcout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_8_s1_THRU_CO ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_8_s1 ),
            .carryout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_9_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_9_s1_THRU_LUT4_0_LC_16_19_2 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_9_s1_THRU_LUT4_0_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_9_s1_THRU_LUT4_0_LC_16_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_9_s1_THRU_LUT4_0_LC_16_19_2  (
            .in0(_gnd_net_),
            .in1(N__11927),
            .in2(N__12460),
            .in3(N__11906),
            .lcout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_9_s1_THRU_CO ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_9_s1 ),
            .carryout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_10_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_10_s1_THRU_LUT4_0_LC_16_19_3 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_10_s1_THRU_LUT4_0_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_10_s1_THRU_LUT4_0_LC_16_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_10_s1_THRU_LUT4_0_LC_16_19_3  (
            .in0(_gnd_net_),
            .in1(N__11903),
            .in2(N__12456),
            .in3(N__11882),
            .lcout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_10_s1_THRU_CO ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_10_s1 ),
            .carryout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_11_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_11_s1_THRU_LUT4_0_LC_16_19_4 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_11_s1_THRU_LUT4_0_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_11_s1_THRU_LUT4_0_LC_16_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_11_s1_THRU_LUT4_0_LC_16_19_4  (
            .in0(_gnd_net_),
            .in1(N__12503),
            .in2(N__12458),
            .in3(N__12473),
            .lcout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_11_s1_THRU_CO ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_11_s1 ),
            .carryout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_12_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_12_s1_THRU_LUT4_0_LC_16_19_5 .C_ON=1'b1;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_12_s1_THRU_LUT4_0_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_12_s1_THRU_LUT4_0_LC_16_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_12_s1_THRU_LUT4_0_LC_16_19_5  (
            .in0(_gnd_net_),
            .in1(N__12439),
            .in2(N__12149),
            .in3(N__12122),
            .lcout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_12_s1_THRU_CO ),
            .ltout(),
            .carryin(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_12_s1 ),
            .carryout(\uart_inst0.uart_inst0.un1_tx_clk_divider_1_cry_13_s1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_clk_divider_esr_14_LC_16_19_6 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_esr_14_LC_16_19_6 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_esr_14_LC_16_19_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \uart_inst0.uart_inst0.tx_clk_divider_esr_14_LC_16_19_6  (
            .in0(_gnd_net_),
            .in1(N__12116),
            .in2(_gnd_net_),
            .in3(N__12119),
            .lcout(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16903),
            .ce(N__12104),
            .sr(N__14637));
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_RNI9D19_0_LC_17_2_0 .C_ON=1'b1;
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_RNI9D19_0_LC_17_2_0 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_RNI9D19_0_LC_17_2_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \fifo_inst.rx_fifo_inst.rRamWrAddr_RNI9D19_0_LC_17_2_0  (
            .in0(_gnd_net_),
            .in1(N__14797),
            .in2(N__14843),
            .in3(N__14840),
            .lcout(rRamWrAddr_RNI9D19_0),
            .ltout(),
            .carryin(bfn_17_2_0_),
            .carryout(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_1_LC_17_2_1 .C_ON=1'b1;
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_1_LC_17_2_1 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_1_LC_17_2_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.rx_fifo_inst.rRamWrAddr_1_LC_17_2_1  (
            .in0(N__16634),
            .in1(N__14155),
            .in2(_gnd_net_),
            .in3(N__12092),
            .lcout(fifo_inst_rx_fifo_inst_rRamWrAddr_1),
            .ltout(),
            .carryin(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_0 ),
            .carryout(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_1 ),
            .clk(N__16982),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_2_LC_17_2_2 .C_ON=1'b1;
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_2_LC_17_2_2 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_2_LC_17_2_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.rx_fifo_inst.rRamWrAddr_2_LC_17_2_2  (
            .in0(N__16637),
            .in1(N__14274),
            .in2(_gnd_net_),
            .in3(N__12089),
            .lcout(fifo_inst_rx_fifo_inst_rRamWrAddr_2),
            .ltout(),
            .carryin(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_1 ),
            .carryout(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_2 ),
            .clk(N__16982),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_2_c_RNIOTMG_LC_17_2_3 .C_ON=1'b1;
    defparam \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_2_c_RNIOTMG_LC_17_2_3 .SEQ_MODE=4'b0000;
    defparam \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_2_c_RNIOTMG_LC_17_2_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_2_c_RNIOTMG_LC_17_2_3  (
            .in0(_gnd_net_),
            .in1(N__14182),
            .in2(_gnd_net_),
            .in3(N__12086),
            .lcout(un1_rRamWrAddr_cry_2_c_RNIOTMG),
            .ltout(),
            .carryin(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_2 ),
            .carryout(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_4_LC_17_2_4 .C_ON=1'b1;
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_4_LC_17_2_4 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_4_LC_17_2_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.rx_fifo_inst.rRamWrAddr_4_LC_17_2_4  (
            .in0(N__16638),
            .in1(N__14308),
            .in2(_gnd_net_),
            .in3(N__12083),
            .lcout(fifo_inst_rx_fifo_inst_rRamWrAddr_4),
            .ltout(),
            .carryin(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_3 ),
            .carryout(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_4 ),
            .clk(N__16982),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_5_LC_17_2_5 .C_ON=1'b1;
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_5_LC_17_2_5 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_5_LC_17_2_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.rx_fifo_inst.rRamWrAddr_5_LC_17_2_5  (
            .in0(N__16635),
            .in1(N__14332),
            .in2(_gnd_net_),
            .in3(N__12080),
            .lcout(fifo_inst_rx_fifo_inst_rRamWrAddr_5),
            .ltout(),
            .carryin(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_4 ),
            .carryout(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_5 ),
            .clk(N__16982),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_6_LC_17_2_6 .C_ON=1'b1;
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_6_LC_17_2_6 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_6_LC_17_2_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.rx_fifo_inst.rRamWrAddr_6_LC_17_2_6  (
            .in0(N__16639),
            .in1(N__14218),
            .in2(_gnd_net_),
            .in3(N__12812),
            .lcout(fifo_inst_rx_fifo_inst_rRamWrAddr_6),
            .ltout(),
            .carryin(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_5 ),
            .carryout(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_6 ),
            .clk(N__16982),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_7_LC_17_2_7 .C_ON=1'b1;
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_7_LC_17_2_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_7_LC_17_2_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.rx_fifo_inst.rRamWrAddr_7_LC_17_2_7  (
            .in0(N__16636),
            .in1(N__14248),
            .in2(_gnd_net_),
            .in3(N__12809),
            .lcout(fifo_inst_rx_fifo_inst_rRamWrAddr_7),
            .ltout(),
            .carryin(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_6 ),
            .carryout(\fifo_inst.rx_fifo_inst.un1_rRamWrAddr_cry_7 ),
            .clk(N__16982),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_8_LC_17_3_0 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_8_LC_17_3_0 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_8_LC_17_3_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \fifo_inst.rx_fifo_inst.rRamWrAddr_8_LC_17_3_0  (
            .in0(N__16659),
            .in1(N__14130),
            .in2(_gnd_net_),
            .in3(N__12806),
            .lcout(fifo_inst_rx_fifo_inst_rRamWrAddr_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16979),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_2_LC_17_3_3 .C_ON=1'b0;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_2_LC_17_3_3 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.tx_fifo_inst.rRamRdAddr_2_LC_17_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \fifo_inst.tx_fifo_inst.rRamRdAddr_2_LC_17_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12796),
            .lcout(fifo_inst_tx_fifo_inst_rRamRdAddr_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16979),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.N_84_mux_i_LC_17_4_5 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.N_84_mux_i_LC_17_4_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.N_84_mux_i_LC_17_4_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.N_84_mux_i_LC_17_4_5  (
            .in0(N__12763),
            .in1(N__12695),
            .in2(N__12656),
            .in3(N__12599),
            .lcout(N_84_mux_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rRxData_6_LC_17_5_0.C_ON=1'b0;
    defparam rRxData_6_LC_17_5_0.SEQ_MODE=4'b1000;
    defparam rRxData_6_LC_17_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 rRxData_6_LC_17_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14653),
            .lcout(rRxDataZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16974),
            .ce(N__12851),
            .sr(_gnd_net_));
    defparam rRxData_1_LC_17_5_1.C_ON=1'b0;
    defparam rRxData_1_LC_17_5_1.SEQ_MODE=4'b1000;
    defparam rRxData_1_LC_17_5_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 rRxData_1_LC_17_5_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14689),
            .lcout(rRxDataZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16974),
            .ce(N__12851),
            .sr(_gnd_net_));
    defparam rRxData_2_LC_17_5_2.C_ON=1'b0;
    defparam rRxData_2_LC_17_5_2.SEQ_MODE=4'b1000;
    defparam rRxData_2_LC_17_5_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 rRxData_2_LC_17_5_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14671),
            .lcout(rRxDataZ0Z_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16974),
            .ce(N__12851),
            .sr(_gnd_net_));
    defparam rRxData_3_LC_17_5_3.C_ON=1'b0;
    defparam rRxData_3_LC_17_5_3.SEQ_MODE=4'b1000;
    defparam rRxData_3_LC_17_5_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 rRxData_3_LC_17_5_3 (
            .in0(N__14750),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(rRxDataZ0Z_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16974),
            .ce(N__12851),
            .sr(_gnd_net_));
    defparam rRxData_0_LC_17_5_4.C_ON=1'b0;
    defparam rRxData_0_LC_17_5_4.SEQ_MODE=4'b1000;
    defparam rRxData_0_LC_17_5_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 rRxData_0_LC_17_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15319),
            .lcout(rRxDataZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16974),
            .ce(N__12851),
            .sr(_gnd_net_));
    defparam rRxData_5_LC_17_5_5.C_ON=1'b0;
    defparam rRxData_5_LC_17_5_5.SEQ_MODE=4'b1000;
    defparam rRxData_5_LC_17_5_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 rRxData_5_LC_17_5_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14710),
            .lcout(rRxDataZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16974),
            .ce(N__12851),
            .sr(_gnd_net_));
    defparam rRxData_7_LC_17_5_7.C_ON=1'b0;
    defparam rRxData_7_LC_17_5_7.SEQ_MODE=4'b1000;
    defparam rRxData_7_LC_17_5_7.LUT_INIT=16'b1100110011001100;
    LogicCell40 rRxData_7_LC_17_5_7 (
            .in0(_gnd_net_),
            .in1(N__14728),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(rRxDataZ0Z_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16974),
            .ce(N__12851),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNO_0_0_LC_17_6_0 .C_ON=1'b1;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNO_0_0_LC_17_6_0 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNO_0_0_LC_17_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNO_0_0_LC_17_6_0  (
            .in0(_gnd_net_),
            .in1(N__15168),
            .in2(N__13157),
            .in3(N__13154),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNO_0_0_0 ),
            .ltout(),
            .carryin(bfn_17_6_0_),
            .carryout(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_1_LC_17_6_1 .C_ON=1'b1;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_1_LC_17_6_1 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_1_LC_17_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_1_LC_17_6_1  (
            .in0(_gnd_net_),
            .in1(N__15198),
            .in2(_gnd_net_),
            .in3(N__12827),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_1 ),
            .ltout(),
            .carryin(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_0 ),
            .carryout(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_1 ),
            .clk(N__16970),
            .ce(),
            .sr(N__13604));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_2_LC_17_6_2 .C_ON=1'b1;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_2_LC_17_6_2 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_2_LC_17_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_2_LC_17_6_2  (
            .in0(_gnd_net_),
            .in1(N__15225),
            .in2(_gnd_net_),
            .in3(N__12824),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_2 ),
            .ltout(),
            .carryin(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_1 ),
            .carryout(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_2 ),
            .clk(N__16970),
            .ce(),
            .sr(N__13604));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNO_0_3_LC_17_6_3 .C_ON=1'b1;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNO_0_3_LC_17_6_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNO_0_3_LC_17_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNO_0_3_LC_17_6_3  (
            .in0(_gnd_net_),
            .in1(N__15253),
            .in2(_gnd_net_),
            .in3(N__12821),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNO_0_0_3 ),
            .ltout(),
            .carryin(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_2 ),
            .carryout(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_4_LC_17_6_4 .C_ON=1'b1;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_4_LC_17_6_4 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_4_LC_17_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_4_LC_17_6_4  (
            .in0(_gnd_net_),
            .in1(N__15042),
            .in2(_gnd_net_),
            .in3(N__12818),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_4 ),
            .ltout(),
            .carryin(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_3 ),
            .carryout(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_4 ),
            .clk(N__16970),
            .ce(),
            .sr(N__13604));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_5_LC_17_6_5 .C_ON=1'b1;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_5_LC_17_6_5 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_5_LC_17_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_5_LC_17_6_5  (
            .in0(_gnd_net_),
            .in1(N__15099),
            .in2(_gnd_net_),
            .in3(N__12815),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_5 ),
            .ltout(),
            .carryin(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_4 ),
            .carryout(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_5 ),
            .clk(N__16970),
            .ce(),
            .sr(N__13604));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_6_LC_17_6_6 .C_ON=1'b1;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_6_LC_17_6_6 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_6_LC_17_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_6_LC_17_6_6  (
            .in0(_gnd_net_),
            .in1(N__15126),
            .in2(_gnd_net_),
            .in3(N__12905),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_6 ),
            .ltout(),
            .carryin(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_5 ),
            .carryout(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_6 ),
            .clk(N__16970),
            .ce(),
            .sr(N__13604));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_7_LC_17_6_7 .C_ON=1'b1;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_7_LC_17_6_7 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_7_LC_17_6_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_7_LC_17_6_7  (
            .in0(_gnd_net_),
            .in1(N__15072),
            .in2(_gnd_net_),
            .in3(N__12902),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_7 ),
            .ltout(),
            .carryin(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_6 ),
            .carryout(\uart_inst0.rx_uart_fifo_inst.un1_rRamWrAddr_cry_7 ),
            .clk(N__16970),
            .ce(),
            .sr(N__13604));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_8_LC_17_7_0 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_8_LC_17_7_0 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_8_LC_17_7_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_8_LC_17_7_0  (
            .in0(_gnd_net_),
            .in1(N__15286),
            .in2(_gnd_net_),
            .in3(N__12899),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16962),
            .ce(),
            .sr(N__13603));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_3_LC_17_7_2 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_3_LC_17_7_2 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_3_LC_17_7_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_3_LC_17_7_2  (
            .in0(N__13146),
            .in1(N__15025),
            .in2(N__15152),
            .in3(N__12896),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16962),
            .ce(),
            .sr(N__13603));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_0_LC_17_7_3 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_0_LC_17_7_3 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_0_LC_17_7_3 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_0_LC_17_7_3  (
            .in0(N__15148),
            .in1(N__12890),
            .in2(N__15026),
            .in3(N__13147),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rRamWrAddrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16962),
            .ce(),
            .sr(N__13603));
    defparam rUartRxState_0_LC_17_8_0.C_ON=1'b0;
    defparam rUartRxState_0_LC_17_8_0.SEQ_MODE=4'b1000;
    defparam rUartRxState_0_LC_17_8_0.LUT_INIT=16'b0000000000100010;
    LogicCell40 rUartRxState_0_LC_17_8_0 (
            .in0(N__14024),
            .in1(N__13041),
            .in2(_gnd_net_),
            .in3(N__13372),
            .lcout(rUartRxStateZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16956),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNO_0_2_LC_17_8_1 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNO_0_2_LC_17_8_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNO_0_2_LC_17_8_1 .LUT_INIT=16'b0000100011100000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rDataCount_RNO_0_2_LC_17_8_1  (
            .in0(N__12966),
            .in1(N__13092),
            .in2(N__14961),
            .in3(N__13142),
            .lcout(\uart_inst0.rx_uart_fifo_inst.un1_rDataCount_c2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNI2JT81_0_2_LC_17_8_2 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNI2JT81_0_2_LC_17_8_2 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNI2JT81_0_2_LC_17_8_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rDataCount_RNI2JT81_0_2_LC_17_8_2  (
            .in0(N__13091),
            .in1(N__12934),
            .in2(N__12968),
            .in3(N__13001),
            .lcout(wUartRxEmpty),
            .ltout(wUartRxEmpty_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNITL9D2_2_LC_17_8_3 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNITL9D2_2_LC_17_8_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNITL9D2_2_LC_17_8_3 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rDataCount_RNITL9D2_2_LC_17_8_3  (
            .in0(_gnd_net_),
            .in1(N__13141),
            .in2(N__12884),
            .in3(N__14950),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rDataCount_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNI2JT81_2_LC_17_8_5 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNI2JT81_2_LC_17_8_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNI2JT81_2_LC_17_8_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rDataCount_RNI2JT81_2_LC_17_8_5  (
            .in0(N__13000),
            .in1(N__12962),
            .in2(N__12935),
            .in3(N__13090),
            .lcout(\uart_inst0.rx_uart_fifo_inst.wUartRxEmpty_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_0_LC_17_9_1 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_0_LC_17_9_1 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_0_LC_17_9_1 .LUT_INIT=16'b0100101110110100;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rDataCount_0_LC_17_9_1  (
            .in0(N__13371),
            .in1(N__14960),
            .in2(N__13156),
            .in3(N__13089),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16949),
            .ce(),
            .sr(N__16429));
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNI3V391_2_LC_17_9_2 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNI3V391_2_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNI3V391_2_LC_17_9_2 .LUT_INIT=16'b1100110011001000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rDataCount_RNI3V391_2_LC_17_9_2  (
            .in0(N__13088),
            .in1(N__14943),
            .in2(N__13003),
            .in3(N__12957),
            .lcout(),
            .ltout(\uart_inst0.rx_uart_fifo_inst.rDataCount_RNI3V391Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNIO7PT1_3_LC_17_9_3 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNIO7PT1_3_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_RNIO7PT1_3_LC_17_9_3 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rDataCount_RNIO7PT1_3_LC_17_9_3  (
            .in0(N__14944),
            .in1(_gnd_net_),
            .in2(N__13061),
            .in3(N__12927),
            .lcout(\uart_inst0.rx_uart_fifo_inst.wRamRdEn ),
            .ltout(\uart_inst0.rx_uart_fifo_inst.wRamRdEn_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_1_LC_17_9_4 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_1_LC_17_9_4 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_1_LC_17_9_4 .LUT_INIT=16'b1011100101000110;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rDataCount_1_LC_17_9_4  (
            .in0(N__13058),
            .in1(N__13012),
            .in2(N__13052),
            .in3(N__12958),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16949),
            .ce(),
            .sr(N__16429));
    defparam rUartRxEn_LC_17_9_5.C_ON=1'b0;
    defparam rUartRxEn_LC_17_9_5.SEQ_MODE=4'b1000;
    defparam rUartRxEn_LC_17_9_5.LUT_INIT=16'b0001000100010001;
    LogicCell40 rUartRxEn_LC_17_9_5 (
            .in0(N__13370),
            .in1(N__13042),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(rUartRxEnZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16949),
            .ce(),
            .sr(N__16429));
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_2_LC_17_9_6 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_2_LC_17_9_6 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_2_LC_17_9_6 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rDataCount_2_LC_17_9_6  (
            .in0(N__13019),
            .in1(N__13013),
            .in2(N__13004),
            .in3(_gnd_net_),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rDataCountZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16949),
            .ce(),
            .sr(N__16429));
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_3_LC_17_9_7 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_3_LC_17_9_7 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.rDataCount_3_LC_17_9_7 .LUT_INIT=16'b1111011100010000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rDataCount_3_LC_17_9_7  (
            .in0(N__14945),
            .in1(N__12974),
            .in2(N__12967),
            .in3(N__12928),
            .lcout(\uart_inst0.wRxWrFull_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16949),
            .ce(),
            .sr(N__16429));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNID4JC2_0_LC_17_10_0 .C_ON=1'b1;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNID4JC2_0_LC_17_10_0 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNID4JC2_0_LC_17_10_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNID4JC2_0_LC_17_10_0  (
            .in0(_gnd_net_),
            .in1(N__13352),
            .in2(N__15798),
            .in3(N__15790),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNID4JC2Z0Z_0 ),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIK0HS_LC_17_10_1 .C_ON=1'b1;
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIK0HS_LC_17_10_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIK0HS_LC_17_10_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIK0HS_LC_17_10_1  (
            .in0(_gnd_net_),
            .in1(N__13180),
            .in2(_gnd_net_),
            .in3(N__13205),
            .lcout(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_0_c_RNIK0HSZ0 ),
            .ltout(),
            .carryin(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_0 ),
            .carryout(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIM3IS_LC_17_10_2 .C_ON=1'b1;
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIM3IS_LC_17_10_2 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIM3IS_LC_17_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIM3IS_LC_17_10_2  (
            .in0(_gnd_net_),
            .in1(N__13168),
            .in2(_gnd_net_),
            .in3(N__13202),
            .lcout(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_1_c_RNIM3ISZ0 ),
            .ltout(),
            .carryin(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_1 ),
            .carryout(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNIO6JS_LC_17_10_3 .C_ON=1'b1;
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNIO6JS_LC_17_10_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNIO6JS_LC_17_10_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNIO6JS_LC_17_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13337),
            .in3(N__13199),
            .lcout(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_2_c_RNIO6JSZ0 ),
            .ltout(),
            .carryin(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_2 ),
            .carryout(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIQ9KS_LC_17_10_4 .C_ON=1'b1;
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIQ9KS_LC_17_10_4 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIQ9KS_LC_17_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIQ9KS_LC_17_10_4  (
            .in0(_gnd_net_),
            .in1(N__13414),
            .in2(_gnd_net_),
            .in3(N__13196),
            .lcout(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_3_c_RNIQ9KSZ0 ),
            .ltout(),
            .carryin(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_3 ),
            .carryout(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNISCLS_LC_17_10_5 .C_ON=1'b1;
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNISCLS_LC_17_10_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNISCLS_LC_17_10_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNISCLS_LC_17_10_5  (
            .in0(_gnd_net_),
            .in1(N__13441),
            .in2(_gnd_net_),
            .in3(N__13193),
            .lcout(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_4_c_RNISCLSZ0 ),
            .ltout(),
            .carryin(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_4 ),
            .carryout(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIUFMS_LC_17_10_6 .C_ON=1'b1;
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIUFMS_LC_17_10_6 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIUFMS_LC_17_10_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIUFMS_LC_17_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13457),
            .in3(N__13190),
            .lcout(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_5_c_RNIUFMSZ0 ),
            .ltout(),
            .carryin(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_5 ),
            .carryout(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI0JNS_LC_17_10_7 .C_ON=1'b1;
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI0JNS_LC_17_10_7 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI0JNS_LC_17_10_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI0JNS_LC_17_10_7  (
            .in0(_gnd_net_),
            .in1(N__13426),
            .in2(_gnd_net_),
            .in3(N__13187),
            .lcout(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_6_c_RNI0JNSZ0 ),
            .ltout(),
            .carryin(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_6 ),
            .carryout(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI2MOS_LC_17_11_0 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI2MOS_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI2MOS_LC_17_11_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI2MOS_LC_17_11_0  (
            .in0(_gnd_net_),
            .in1(N__13394),
            .in2(_gnd_net_),
            .in3(N__13184),
            .lcout(\uart_inst0.rx_uart_fifo_inst.un1_rRamRdAddr_cry_7_c_RNI2MOSZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNI17A54_1_LC_17_11_1 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNI17A54_1_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNI17A54_1_LC_17_11_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNI17A54_1_LC_17_11_1  (
            .in0(N__13385),
            .in1(N__13181),
            .in2(N__13403),
            .in3(N__13169),
            .lcout(\uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_0_LC_17_11_2 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_0_LC_17_11_2 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_0_LC_17_11_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_0_LC_17_11_2  (
            .in0(_gnd_net_),
            .in1(N__16693),
            .in2(_gnd_net_),
            .in3(N__13483),
            .lcout(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNIA98R1_4_LC_17_11_6 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNIA98R1_4_LC_17_11_6 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNIA98R1_4_LC_17_11_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNIA98R1_4_LC_17_11_6  (
            .in0(N__13456),
            .in1(N__13442),
            .in2(N__13430),
            .in3(N__13415),
            .lcout(\uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNIA1EC1_8_LC_17_11_7 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNIA1EC1_8_LC_17_11_7 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNIA1EC1_8_LC_17_11_7 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_RNIA1EC1_8_LC_17_11_7  (
            .in0(N__13393),
            .in1(N__13333),
            .in2(_gnd_net_),
            .in3(N__13351),
            .lcout(\uart_inst0.rx_uart_fifo_inst.un20_rRamRdAddr_0_sqmuxa_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_0_LC_17_12_2 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_0_LC_17_12_2 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_0_LC_17_12_2 .LUT_INIT=16'b1100010011001100;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_0_LC_17_12_2  (
            .in0(N__15824),
            .in1(N__15470),
            .in2(N__13379),
            .in3(N__14963),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16936),
            .ce(),
            .sr(N__13602));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_3_LC_17_12_7 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_3_LC_17_12_7 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_3_LC_17_12_7 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamRdAddr_3_LC_17_12_7  (
            .in0(N__15823),
            .in1(N__15755),
            .in2(_gnd_net_),
            .in3(N__15800),
            .lcout(\uart_inst0.rx_uart_fifo_inst.rRamRdAddrZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16936),
            .ce(),
            .sr(N__13602));
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_RNINTCJ_2_LC_17_13_1 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_RNINTCJ_2_LC_17_13_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_RNINTCJ_2_LC_17_13_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \uart_inst0.uart_inst0.rx_bits_remaining_RNINTCJ_2_LC_17_13_1  (
            .in0(N__15891),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15637),
            .lcout(\uart_inst0.uart_inst0.N_274_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_RNO_0_2_LC_17_13_3 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_RNO_0_2_LC_17_13_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_RNO_0_2_LC_17_13_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uart_inst0.uart_inst0.rx_bits_remaining_RNO_0_2_LC_17_13_3  (
            .in0(N__16035),
            .in1(N__15969),
            .in2(_gnd_net_),
            .in3(N__15922),
            .lcout(\uart_inst0.uart_inst0.un1_rx_bits_remaining_c1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_state_RNID5M13_2_LC_17_13_5 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_state_RNID5M13_2_LC_17_13_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_state_RNID5M13_2_LC_17_13_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uart_inst0.uart_inst0.rx_state_RNID5M13_2_LC_17_13_5  (
            .in0(N__16036),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15920),
            .lcout(\uart_inst0.uart_inst0.rx_bits_remaining_2_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_state_RNI4UTC3_1_LC_17_13_6 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_state_RNI4UTC3_1_LC_17_13_6 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_state_RNI4UTC3_1_LC_17_13_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \uart_inst0.uart_inst0.rx_state_RNI4UTC3_1_LC_17_13_6  (
            .in0(N__15921),
            .in1(N__13298),
            .in2(_gnd_net_),
            .in3(N__13265),
            .lcout(\uart_inst0.uart_inst0.rx_state_2_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_countdown_RNID5M13_0_LC_17_13_7 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_countdown_RNID5M13_0_LC_17_13_7 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_countdown_RNID5M13_0_LC_17_13_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \uart_inst0.uart_inst0.rx_countdown_RNID5M13_0_LC_17_13_7  (
            .in0(N__14081),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14035),
            .lcout(\uart_inst0.uart_inst0.rRxData_0_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_state_RNO_0_3_LC_17_14_1 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_state_RNO_0_3_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_state_RNO_0_3_LC_17_14_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uart_inst0.uart_inst0.rx_state_RNO_0_3_LC_17_14_1  (
            .in0(N__13946),
            .in1(N__13771),
            .in2(_gnd_net_),
            .in3(N__13829),
            .lcout(),
            .ltout(\uart_inst0.uart_inst0.N_273_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_state_3_LC_17_14_2 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_state_3_LC_17_14_2 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_state_3_LC_17_14_2 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \uart_inst0.uart_inst0.rx_state_3_LC_17_14_2  (
            .in0(N__15655),
            .in1(N__13720),
            .in2(N__13790),
            .in3(N__13738),
            .lcout(\uart_inst0.uart_inst0.rx_stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16929),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_RNINTCJ_3_LC_17_14_3 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_RNINTCJ_3_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_RNINTCJ_3_LC_17_14_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uart_inst0.uart_inst0.rx_bits_remaining_RNINTCJ_3_LC_17_14_3  (
            .in0(_gnd_net_),
            .in1(N__13696),
            .in2(_gnd_net_),
            .in3(N__15965),
            .lcout(\uart_inst0.uart_inst0.rx_state_srsts_0_a5_0_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_RNO_0_3_LC_17_14_6 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_RNO_0_3_LC_17_14_6 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_RNO_0_3_LC_17_14_6 .LUT_INIT=16'b1100010000000000;
    LogicCell40 \uart_inst0.uart_inst0.rx_bits_remaining_RNO_0_3_LC_17_14_6  (
            .in0(N__13719),
            .in1(N__16037),
            .in2(N__15973),
            .in3(N__15923),
            .lcout(),
            .ltout(\uart_inst0.uart_inst0.un1_rx_bits_remaining_c3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_3_LC_17_14_7 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_3_LC_17_14_7 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_3_LC_17_14_7 .LUT_INIT=16'b0010000100010010;
    LogicCell40 \uart_inst0.uart_inst0.rx_bits_remaining_3_LC_17_14_7  (
            .in0(N__13697),
            .in1(N__15864),
            .in2(N__13700),
            .in3(N__15654),
            .lcout(\uart_inst0.uart_inst0.rx_bits_remainingZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16929),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_countdown_2_LC_17_16_4 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_countdown_2_LC_17_16_4 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.tx_countdown_2_LC_17_16_4 .LUT_INIT=16'b0011001011011100;
    LogicCell40 \uart_inst0.uart_inst0.tx_countdown_2_LC_17_16_4  (
            .in0(N__13685),
            .in1(N__13629),
            .in2(N__13643),
            .in3(N__14459),
            .lcout(\uart_inst0.uart_inst0.tx_countdownZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16922),
            .ce(),
            .sr(N__13597));
    defparam \uart_inst0.uart_inst0.tx_clk_divider_3_LC_17_17_4 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_3_LC_17_17_4 .SEQ_MODE=4'b1001;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_3_LC_17_17_4 .LUT_INIT=16'b1101110100100010;
    LogicCell40 \uart_inst0.uart_inst0.tx_clk_divider_3_LC_17_17_4  (
            .in0(N__13548),
            .in1(N__13490),
            .in2(_gnd_net_),
            .in3(N__14419),
            .lcout(\uart_inst0.uart_inst0.tx_clk_dividerZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16916),
            .ce(),
            .sr(N__14638));
    defparam \uart_inst0.uart_inst0.tx_countdown_RNO_2_2_LC_17_18_3 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_countdown_RNO_2_2_LC_17_18_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_countdown_RNO_2_2_LC_17_18_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uart_inst0.uart_inst0.tx_countdown_RNO_2_2_LC_17_18_3  (
            .in0(N__14593),
            .in1(N__14551),
            .in2(_gnd_net_),
            .in3(N__14504),
            .lcout(),
            .ltout(\uart_inst0.uart_inst0.tx_m5_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_countdown_RNO_1_2_LC_17_18_4 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_countdown_RNO_1_2_LC_17_18_4 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_countdown_RNO_1_2_LC_17_18_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uart_inst0.uart_inst0.tx_countdown_RNO_1_2_LC_17_18_4  (
            .in0(N__14489),
            .in1(N__14380),
            .in2(N__14480),
            .in3(N__14477),
            .lcout(\uart_inst0.uart_inst0.tx_N_11_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.tx_clk_divider_RNIAEQ11_0_LC_17_18_5 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_RNIAEQ11_0_LC_17_18_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.uart_inst0.tx_clk_divider_RNIAEQ11_0_LC_17_18_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_inst0.uart_inst0.tx_clk_divider_RNIAEQ11_0_LC_17_18_5  (
            .in0(N__14448),
            .in1(N__14431),
            .in2(N__14420),
            .in3(N__14397),
            .lcout(\uart_inst0.uart_inst0.tx_m5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.ft2232h_inst.rRxData_5_LC_18_1_1 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rRxData_5_LC_18_1_1 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rRxData_5_LC_18_1_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_inst.ft2232h_inst.rRxData_5_LC_18_1_1  (
            .in0(N__14366),
            .in1(N__17040),
            .in2(_gnd_net_),
            .in3(N__14356),
            .lcout(\fifo_inst.wRxWrData_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16988),
            .ce(),
            .sr(N__16368));
    defparam \uart_inst0.tx_uart_fifo_inst.m54_e_5_LC_18_2_0 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m54_e_5_LC_18_2_0 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m54_e_5_LC_18_2_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m54_e_5_LC_18_2_0  (
            .in0(N__14331),
            .in1(N__14307),
            .in2(N__14287),
            .in3(N__16658),
            .lcout(),
            .ltout(\uart_inst0.tx_uart_fifo_inst.m54_eZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m54_e_LC_18_2_1 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m54_e_LC_18_2_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m54_e_LC_18_2_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m54_e_LC_18_2_1  (
            .in0(N__14244),
            .in1(N__14217),
            .in2(N__14201),
            .in3(N__14108),
            .lcout(\uart_inst0.tx_uart_fifo_inst.N_91 ),
            .ltout(\uart_inst0.tx_uart_fifo_inst.N_91_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_3_LC_18_2_2 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_3_LC_18_2_2 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_3_LC_18_2_2 .LUT_INIT=16'b0101001100000000;
    LogicCell40 \fifo_inst.rx_fifo_inst.rRamWrAddr_3_LC_18_2_2  (
            .in0(N__14842),
            .in1(N__16657),
            .in2(N__14198),
            .in3(N__14195),
            .lcout(fifo_inst_rx_fifo_inst_rRamWrAddr_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16984),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.m54_e_6_LC_18_2_4 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.m54_e_6_LC_18_2_4 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.m54_e_6_LC_18_2_4 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.m54_e_6_LC_18_2_4  (
            .in0(N__14181),
            .in1(N__14154),
            .in2(N__14131),
            .in3(N__14796),
            .lcout(\uart_inst0.tx_uart_fifo_inst.m54_eZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_0_LC_18_2_7 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_0_LC_18_2_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.rRamWrAddr_0_LC_18_2_7 .LUT_INIT=16'b0000001010001010;
    LogicCell40 \fifo_inst.rx_fifo_inst.rRamWrAddr_0_LC_18_2_7  (
            .in0(N__14855),
            .in1(N__14849),
            .in2(N__16700),
            .in3(N__14841),
            .lcout(fifo_inst_rx_fifo_inst_rRamWrAddr_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16984),
            .ce(),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_4_LC_18_3_1 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_4_LC_18_3_1 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_4_LC_18_3_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_4_LC_18_3_1  (
            .in0(N__15412),
            .in1(N__14770),
            .in2(_gnd_net_),
            .in3(N__14780),
            .lcout(wRxData_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_4C_net ),
            .ce(N__15308),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_3_LC_18_3_7 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_3_LC_18_3_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_3_LC_18_3_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_3_LC_18_3_7  (
            .in0(N__15411),
            .in1(N__14749),
            .in2(_gnd_net_),
            .in3(N__14756),
            .lcout(wRxData_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_4C_net ),
            .ce(N__15308),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7_LC_18_4_0 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7_LC_18_4_0 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7_LC_18_4_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7_LC_18_4_0  (
            .in0(N__15402),
            .in1(N__14735),
            .in2(_gnd_net_),
            .in3(N__14729),
            .lcout(wRxData_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7C_net ),
            .ce(N__15304),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_5_LC_18_4_2 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_5_LC_18_4_2 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_5_LC_18_4_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_5_LC_18_4_2  (
            .in0(N__15400),
            .in1(N__14711),
            .in2(_gnd_net_),
            .in3(N__14717),
            .lcout(wRxData_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7C_net ),
            .ce(N__15304),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_1_LC_18_4_3 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_1_LC_18_4_3 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_1_LC_18_4_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_1_LC_18_4_3  (
            .in0(N__14693),
            .in1(N__14699),
            .in2(_gnd_net_),
            .in3(N__15398),
            .lcout(wRxData_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7C_net ),
            .ce(N__15304),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_2_LC_18_4_4 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_2_LC_18_4_4 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_2_LC_18_4_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_2_LC_18_4_4  (
            .in0(N__15399),
            .in1(N__14672),
            .in2(_gnd_net_),
            .in3(N__14678),
            .lcout(wRxData_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7C_net ),
            .ce(N__15304),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_6_LC_18_4_6 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_6_LC_18_4_6 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_6_LC_18_4_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_6_LC_18_4_6  (
            .in0(N__15401),
            .in1(N__14654),
            .in2(_gnd_net_),
            .in3(N__14660),
            .lcout(wRxData_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7C_net ),
            .ce(N__15304),
            .sr(_gnd_net_));
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_0_LC_18_4_7 .C_ON=1'b0;
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_0_LC_18_4_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_0_LC_18_4_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \fifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_0_LC_18_4_7  (
            .in0(N__15320),
            .in1(N__15425),
            .in2(_gnd_net_),
            .in3(N__15397),
            .lcout(wRxData_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVfifo_inst.rx_fifo_inst.ram512x8_inst.RDATA_7C_net ),
            .ce(N__15304),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNIRP0T_8_LC_18_7_1 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNIRP0T_8_LC_18_7_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNIRP0T_8_LC_18_7_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNIRP0T_8_LC_18_7_1  (
            .in0(_gnd_net_),
            .in1(N__15276),
            .in2(_gnd_net_),
            .in3(N__15252),
            .lcout(),
            .ltout(\uart_inst0.rx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNIMIH82_0_LC_18_7_2 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNIMIH82_0_LC_18_7_2 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNIMIH82_0_LC_18_7_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNIMIH82_0_LC_18_7_2  (
            .in0(N__15229),
            .in1(N__15202),
            .in2(N__15182),
            .in3(N__15172),
            .lcout(\uart_inst0.rx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNIMJ1Q1_4_LC_18_7_5 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNIMJ1Q1_4_LC_18_7_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNIMJ1Q1_4_LC_18_7_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.rRamWrAddr_RNIMJ1Q1_4_LC_18_7_5  (
            .in0(N__15127),
            .in1(N__15100),
            .in2(N__15079),
            .in3(N__15043),
            .lcout(\uart_inst0.rx_uart_fifo_inst.un24_rRamWrAddr_0_sqmuxa_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_5_LC_18_8_0 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_5_LC_18_8_0 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_5_LC_18_8_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_5_LC_18_8_0  (
            .in0(N__15014),
            .in1(N__15007),
            .in2(_gnd_net_),
            .in3(N__14947),
            .lcout(wUartRxData_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_5C_net ),
            .ce(N__14879),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_6_LC_18_8_1 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_6_LC_18_8_1 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_6_LC_18_8_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_6_LC_18_8_1  (
            .in0(N__14946),
            .in1(_gnd_net_),
            .in2(N__14993),
            .in3(N__14983),
            .lcout(wUartRxData_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_5C_net ),
            .ce(N__14879),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_7_LC_18_8_2 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_7_LC_18_8_2 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_7_LC_18_8_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_7_LC_18_8_2  (
            .in0(N__14893),
            .in1(N__14969),
            .in2(_gnd_net_),
            .in3(N__14948),
            .lcout(wUartRxData_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_5C_net ),
            .ce(N__14879),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_0_LC_18_9_0 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_0_LC_18_9_0 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_0_LC_18_9_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_0_LC_18_9_0  (
            .in0(N__14870),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(wUartRxData_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net ),
            .ce(N__15789),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_1_LC_18_9_1 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_1_LC_18_9_1 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_1_LC_18_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_1_LC_18_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15572),
            .lcout(wUartRxData_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net ),
            .ce(N__15789),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_2_LC_18_9_2 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_2_LC_18_9_2 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_2_LC_18_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_2_LC_18_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15557),
            .lcout(wUartRxData_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net ),
            .ce(N__15789),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_3_LC_18_9_3 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_3_LC_18_9_3 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_3_LC_18_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_3_LC_18_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15542),
            .lcout(wUartRxData_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net ),
            .ce(N__15789),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_4_LC_18_9_4 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_4_LC_18_9_4 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_4_LC_18_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_4_LC_18_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15527),
            .lcout(wUartRxData_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuart_inst0.rx_uart_fifo_inst.ram512x8_inst.RDATA_0C_net ),
            .ce(N__15789),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_5_LC_18_10_0 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_5_LC_18_10_0 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_5_LC_18_10_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_5_LC_18_10_0  (
            .in0(_gnd_net_),
            .in1(N__16684),
            .in2(_gnd_net_),
            .in3(N__15511),
            .lcout(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_3_LC_18_10_1 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_3_LC_18_10_1 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_3_LC_18_10_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_3_LC_18_10_1  (
            .in0(_gnd_net_),
            .in1(N__16686),
            .in2(_gnd_net_),
            .in3(N__15490),
            .lcout(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_LC_18_10_2 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_LC_18_10_2 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_LC_18_10_2 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_LC_18_10_2  (
            .in0(N__15822),
            .in1(N__15466),
            .in2(N__16703),
            .in3(N__15794),
            .lcout(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_4_LC_18_10_3 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_4_LC_18_10_3 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_4_LC_18_10_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_4_LC_18_10_3  (
            .in0(_gnd_net_),
            .in1(N__16687),
            .in2(_gnd_net_),
            .in3(N__15445),
            .lcout(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_2_LC_18_10_4 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_2_LC_18_10_4 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_2_LC_18_10_4 .LUT_INIT=16'b0001010100000000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_2_LC_18_10_4  (
            .in0(N__16685),
            .in1(N__15821),
            .in2(N__15799),
            .in3(N__15751),
            .lcout(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_6_LC_18_10_5 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_6_LC_18_10_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_6_LC_18_10_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_6_LC_18_10_5  (
            .in0(_gnd_net_),
            .in1(N__16688),
            .in2(_gnd_net_),
            .in3(N__15730),
            .lcout(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_1_LC_18_10_6 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_1_LC_18_10_6 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_1_LC_18_10_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_1_LC_18_10_6  (
            .in0(_gnd_net_),
            .in1(N__16683),
            .in2(_gnd_net_),
            .in3(N__15709),
            .lcout(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_7_LC_18_10_7 .C_ON=1'b0;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_7_LC_18_10_7 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_7_LC_18_10_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_7_LC_18_10_7  (
            .in0(_gnd_net_),
            .in1(N__16689),
            .in2(_gnd_net_),
            .in3(N__15688),
            .lcout(\uart_inst0.rx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_2_LC_18_11_2 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_2_LC_18_11_2 .SEQ_MODE=4'b1001;
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_2_LC_18_11_2 .LUT_INIT=16'b1110000101111000;
    LogicCell40 \uart_inst0.uart_inst0.rx_bits_remaining_2_LC_18_11_2  (
            .in0(N__15896),
            .in1(N__15668),
            .in2(N__15641),
            .in3(N__15659),
            .lcout(\uart_inst0.uart_inst0.rx_bits_remainingZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16945),
            .ce(),
            .sr(N__15874));
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_0_LC_18_11_3 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_0_LC_18_11_3 .SEQ_MODE=4'b1001;
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_0_LC_18_11_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \uart_inst0.uart_inst0.rx_bits_remaining_0_LC_18_11_3  (
            .in0(N__15938),
            .in1(N__15964),
            .in2(_gnd_net_),
            .in3(N__16049),
            .lcout(\uart_inst0.uart_inst0.rx_bits_remainingZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16945),
            .ce(),
            .sr(N__15874));
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_1_LC_18_11_5 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_1_LC_18_11_5 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_1_LC_18_11_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_1_LC_18_11_5  (
            .in0(_gnd_net_),
            .in1(N__16694),
            .in2(_gnd_net_),
            .in3(N__15622),
            .lcout(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_4_LC_18_11_7 .C_ON=1'b0;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_4_LC_18_11_7 .SEQ_MODE=4'b0000;
    defparam \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_4_LC_18_11_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNO_4_LC_18_11_7  (
            .in0(_gnd_net_),
            .in1(N__16695),
            .in2(_gnd_net_),
            .in3(N__15596),
            .lcout(\uart_inst0.tx_uart_fifo_inst.ram512x8_inst.mem_mem_0_0_RNOZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uart_inst0.uart_inst0.rRxData_esr_1_LC_18_12_0 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rRxData_esr_1_LC_18_12_0 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rRxData_esr_1_LC_18_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.uart_inst0.rRxData_esr_1_LC_18_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16081),
            .lcout(\uart_inst0.wRxWrData_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16940),
            .ce(N__16067),
            .sr(N__16454));
    defparam \uart_inst0.uart_inst0.rRxData_esr_4_LC_18_12_1 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rRxData_esr_4_LC_18_12_1 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rRxData_esr_4_LC_18_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.uart_inst0.rRxData_esr_4_LC_18_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16162),
            .lcout(\uart_inst0.wRxWrData_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16940),
            .ce(N__16067),
            .sr(N__16454));
    defparam \uart_inst0.uart_inst0.rRxData_esr_3_LC_18_12_3 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rRxData_esr_3_LC_18_12_3 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rRxData_esr_3_LC_18_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.uart_inst0.rRxData_esr_3_LC_18_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16210),
            .lcout(\uart_inst0.wRxWrData_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16940),
            .ce(N__16067),
            .sr(N__16454));
    defparam \uart_inst0.uart_inst0.rRxData_esr_0_LC_18_12_4 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rRxData_esr_0_LC_18_12_4 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rRxData_esr_0_LC_18_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.uart_inst0.rRxData_esr_0_LC_18_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16192),
            .lcout(\uart_inst0.wRxWrData_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16940),
            .ce(N__16067),
            .sr(N__16454));
    defparam \uart_inst0.uart_inst0.rRxData_esr_5_LC_18_12_5 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rRxData_esr_5_LC_18_12_5 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rRxData_esr_5_LC_18_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.uart_inst0.rRxData_esr_5_LC_18_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16114),
            .lcout(\uart_inst0.wRxWrData_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16940),
            .ce(N__16067),
            .sr(N__16454));
    defparam \uart_inst0.uart_inst0.rRxData_esr_6_LC_18_12_6 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rRxData_esr_6_LC_18_12_6 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rRxData_esr_6_LC_18_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.uart_inst0.rRxData_esr_6_LC_18_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16148),
            .lcout(\uart_inst0.wRxWrData_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16940),
            .ce(N__16067),
            .sr(N__16454));
    defparam \uart_inst0.uart_inst0.rRxData_esr_2_LC_18_13_5 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rRxData_esr_2_LC_18_13_5 .SEQ_MODE=4'b1000;
    defparam \uart_inst0.uart_inst0.rRxData_esr_2_LC_18_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uart_inst0.uart_inst0.rRxData_esr_2_LC_18_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16096),
            .lcout(\uart_inst0.wRxWrData_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16937),
            .ce(N__16066),
            .sr(N__16455));
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_1_LC_18_14_5 .C_ON=1'b0;
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_1_LC_18_14_5 .SEQ_MODE=4'b1001;
    defparam \uart_inst0.uart_inst0.rx_bits_remaining_1_LC_18_14_5 .LUT_INIT=16'b1010011010101010;
    LogicCell40 \uart_inst0.uart_inst0.rx_bits_remaining_1_LC_18_14_5  (
            .in0(N__15895),
            .in1(N__16048),
            .in2(N__15974),
            .in3(N__15933),
            .lcout(\uart_inst0.uart_inst0.rx_bits_remainingZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16932),
            .ce(),
            .sr(N__15875));
    defparam \fifo_inst.ft2232h_inst.rRxData_2_LC_20_3_0 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rRxData_2_LC_20_3_0 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rRxData_2_LC_20_3_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_inst.ft2232h_inst.rRxData_2_LC_20_3_0  (
            .in0(N__15848),
            .in1(N__17060),
            .in2(_gnd_net_),
            .in3(N__15836),
            .lcout(\fifo_inst.wRxWrData_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16989),
            .ce(),
            .sr(N__16419));
    defparam \fifo_inst.ft2232h_inst.rRxData_1_LC_20_3_2 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rRxData_1_LC_20_3_2 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rRxData_1_LC_20_3_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_inst.ft2232h_inst.rRxData_1_LC_20_3_2  (
            .in0(N__17225),
            .in1(N__17059),
            .in2(_gnd_net_),
            .in3(N__17209),
            .lcout(\fifo_inst.wRxWrData_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16989),
            .ce(),
            .sr(N__16419));
    defparam \fifo_inst.ft2232h_inst.rRxData_3_LC_20_3_3 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rRxData_3_LC_20_3_3 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rRxData_3_LC_20_3_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_inst.ft2232h_inst.rRxData_3_LC_20_3_3  (
            .in0(N__17061),
            .in1(N__17195),
            .in2(_gnd_net_),
            .in3(N__17182),
            .lcout(\fifo_inst.wRxWrData_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16989),
            .ce(),
            .sr(N__16419));
    defparam \fifo_inst.ft2232h_inst.rRxData_4_LC_20_3_4 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rRxData_4_LC_20_3_4 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rRxData_4_LC_20_3_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_inst.ft2232h_inst.rRxData_4_LC_20_3_4  (
            .in0(N__17168),
            .in1(N__17062),
            .in2(_gnd_net_),
            .in3(N__17156),
            .lcout(\fifo_inst.wRxWrData_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16989),
            .ce(),
            .sr(N__16419));
    defparam \fifo_inst.ft2232h_inst.rRxData_0_LC_20_3_6 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rRxData_0_LC_20_3_6 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rRxData_0_LC_20_3_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_inst.ft2232h_inst.rRxData_0_LC_20_3_6  (
            .in0(N__17144),
            .in1(N__17058),
            .in2(_gnd_net_),
            .in3(N__17129),
            .lcout(\fifo_inst.wRxWrData_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16989),
            .ce(),
            .sr(N__16419));
    defparam \fifo_inst.ft2232h_inst.rRxData_7_LC_20_3_7 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rRxData_7_LC_20_3_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rRxData_7_LC_20_3_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \fifo_inst.ft2232h_inst.rRxData_7_LC_20_3_7  (
            .in0(N__17063),
            .in1(N__17117),
            .in2(_gnd_net_),
            .in3(N__17096),
            .lcout(\fifo_inst.wRxWrData_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16989),
            .ce(),
            .sr(N__16419));
    defparam \fifo_inst.ft2232h_inst.rRxData_6_LC_20_4_7 .C_ON=1'b0;
    defparam \fifo_inst.ft2232h_inst.rRxData_6_LC_20_4_7 .SEQ_MODE=4'b1000;
    defparam \fifo_inst.ft2232h_inst.rRxData_6_LC_20_4_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \fifo_inst.ft2232h_inst.rRxData_6_LC_20_4_7  (
            .in0(N__17084),
            .in1(N__17057),
            .in2(_gnd_net_),
            .in3(N__17005),
            .lcout(\fifo_inst.wRxWrData_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__16987),
            .ce(),
            .sr(N__16421));
endmodule // top
